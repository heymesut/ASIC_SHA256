
module message_schedule_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module message_schedule_DW01_add_2 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3;
  wire   [31:2] carry;

  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX4 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX4 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX4 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX4 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX4 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX4 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX4 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX4 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  NOR2X1 U1 ( .A(n2), .B(n3), .Y(n1) );
  CLKINVX4 U2 ( .A(A[0]), .Y(n2) );
  INVXL U3 ( .A(B[0]), .Y(n3) );
  XOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module message_schedule_DW01_add_1 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n19, n21, n23, n16, n17, n18, n20, n22, n24, n25, n26, n27;
  wire   [31:2] carry;

  ADDFHX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX4 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(n27), .CO(carry[21]), .S(SUM[20])
         );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX4 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX4 U1_18 ( .A(A[18]), .B(B[18]), .CI(n22), .CO(carry[19]), .S(SUM[18])
         );
  ADDFHX4 U1_26 ( .A(A[26]), .B(B[26]), .CI(n26), .CO(carry[27]), .S(SUM[26])
         );
  ADDFHX4 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX4 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX4 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  INVX1 U1 ( .A(A[17]), .Y(n25) );
  INVX1 U2 ( .A(B[17]), .Y(n24) );
  XOR3X2 U3 ( .A(A[8]), .B(B[8]), .C(carry[8]), .Y(SUM[8]) );
  OAI2BB2X4 U4 ( .B0(n16), .B1(n17), .A0N(n21), .A1N(carry[19]), .Y(n27) );
  INVX1 U5 ( .A(B[19]), .Y(n16) );
  INVX1 U6 ( .A(A[19]), .Y(n17) );
  OAI2BB2X4 U7 ( .B0(n18), .B1(n20), .A0N(n19), .A1N(carry[25]), .Y(n26) );
  INVX1 U8 ( .A(B[25]), .Y(n18) );
  INVX1 U9 ( .A(A[25]), .Y(n20) );
  AND2X2 U10 ( .A(A[0]), .B(B[0]), .Y(n1) );
  OAI2BB2X4 U11 ( .B0(n24), .B1(n25), .A0N(n23), .A1N(carry[17]), .Y(n22) );
  XOR2X4 U12 ( .A(carry[17]), .B(n23), .Y(SUM[17]) );
  XOR2X1 U13 ( .A(carry[19]), .B(n21), .Y(SUM[19]) );
  XOR2X1 U14 ( .A(carry[25]), .B(n19), .Y(SUM[25]) );
  XOR2X1 U15 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  XOR2X1 U16 ( .A(A[17]), .B(B[17]), .Y(n23) );
  XOR2X1 U17 ( .A(A[19]), .B(B[19]), .Y(n21) );
  XOR2X1 U18 ( .A(A[25]), .B(B[25]), .Y(n19) );
endmodule


module message_schedule_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n27, n41, n42, n43, n44, n45, n46, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n47, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74;
  wire   [31:2] carry;

  AND2X2 U1 ( .A(A[0]), .B(B[0]), .Y(n27) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX4 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX4 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX4 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX4 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n27), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  NAND2X2 U2 ( .A(n69), .B(carry[26]), .Y(n50) );
  CLKINVX3 U3 ( .A(B[26]), .Y(n68) );
  XOR2X4 U4 ( .A(A[5]), .B(B[5]), .Y(n46) );
  NAND2X4 U5 ( .A(n46), .B(carry[5]), .Y(n66) );
  XOR2X1 U6 ( .A(carry[5]), .B(n46), .Y(SUM[5]) );
  OAI2BB1X2 U7 ( .A0N(A[17]), .A1N(B[17]), .B0(n60), .Y(n73) );
  OAI2BB1X4 U8 ( .A0N(n73), .A1N(A[18]), .B0(n45), .Y(carry[19]) );
  OAI21X4 U9 ( .A0(A[18]), .A1(n44), .B0(B[18]), .Y(n45) );
  XNOR2X4 U10 ( .A(A[6]), .B(B[6]), .Y(n42) );
  OAI2BB1X4 U11 ( .A0N(A[17]), .A1N(B[17]), .B0(n60), .Y(n44) );
  AND2X2 U12 ( .A(A[27]), .B(carry[27]), .Y(n72) );
  OR2X2 U13 ( .A(carry[27]), .B(A[27]), .Y(n49) );
  OAI2BB1X4 U14 ( .A0N(A[26]), .A1N(B[26]), .B0(n50), .Y(carry[27]) );
  OR2X2 U15 ( .A(A[28]), .B(B[28]), .Y(n47) );
  NAND2X4 U16 ( .A(n47), .B(carry[28]), .Y(n43) );
  OAI2BB1X4 U17 ( .A0N(A[28]), .A1N(B[28]), .B0(n43), .Y(carry[29]) );
  OAI21X4 U18 ( .A0(A[23]), .A1(B[23]), .B0(carry[23]), .Y(n57) );
  OAI21X4 U19 ( .A0(A[24]), .A1(n54), .B0(B[24]), .Y(n55) );
  OAI2BB1X4 U20 ( .A0N(A[23]), .A1N(B[23]), .B0(n57), .Y(n54) );
  OAI2BB2X4 U21 ( .B0(n41), .B1(n42), .A0N(B[6]), .A1N(A[6]), .Y(carry[7]) );
  AND2X4 U22 ( .A(n65), .B(n66), .Y(n41) );
  CMPR32X1 U23 ( .A(A[22]), .B(B[22]), .C(carry[22]), .CO(n64) );
  NAND2X1 U24 ( .A(B[5]), .B(A[5]), .Y(n65) );
  XOR2X1 U25 ( .A(n42), .B(n41), .Y(SUM[6]) );
  NOR2X2 U26 ( .A(n71), .B(n72), .Y(n48) );
  NAND2X1 U27 ( .A(n67), .B(n68), .Y(n69) );
  INVXL U28 ( .A(A[26]), .Y(n67) );
  XNOR2X1 U29 ( .A(n70), .B(n48), .Y(SUM[28]) );
  XOR2XL U30 ( .A(A[28]), .B(B[28]), .Y(n70) );
  AND2X2 U31 ( .A(B[27]), .B(n49), .Y(n71) );
  OAI2BB1X4 U32 ( .A0N(n54), .A1N(A[24]), .B0(n55), .Y(carry[25]) );
  OAI2BB1XL U33 ( .A0N(A[17]), .A1N(B[17]), .B0(n60), .Y(n74) );
  OAI21X4 U34 ( .A0(A[17]), .A1(B[17]), .B0(carry[17]), .Y(n60) );
  XNOR2X1 U35 ( .A(A[26]), .B(B[26]), .Y(n51) );
  OR2XL U36 ( .A(carry[25]), .B(A[25]), .Y(n53) );
  OAI2BB1X1 U37 ( .A0N(A[16]), .A1N(B[16]), .B0(n63), .Y(n61) );
  OAI21XL U38 ( .A0(A[16]), .A1(B[16]), .B0(carry[16]), .Y(n63) );
  XOR2X1 U39 ( .A(n51), .B(n52), .Y(SUM[26]) );
  AOI22XL U40 ( .A0(B[25]), .A1(n53), .B0(A[25]), .B1(carry[25]), .Y(n52) );
  XOR2X1 U41 ( .A(n54), .B(n56), .Y(SUM[24]) );
  XOR2X1 U42 ( .A(B[24]), .B(A[24]), .Y(n56) );
  XOR2X1 U43 ( .A(A[23]), .B(n58), .Y(SUM[23]) );
  XOR2X1 U44 ( .A(n64), .B(B[23]), .Y(n58) );
  XOR2X1 U45 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U46 ( .A(n61), .B(n62), .Y(SUM[17]) );
  XOR2X1 U47 ( .A(B[17]), .B(A[17]), .Y(n62) );
  XOR2X1 U48 ( .A(n74), .B(n59), .Y(SUM[18]) );
  XOR2X1 U49 ( .A(B[18]), .B(A[18]), .Y(n59) );
endmodule


module message_schedule ( clk, reset, data, write_enable, inner_busy, Wt );
  input [31:0] data;
  output [31:0] Wt;
  input clk, reset, write_enable, inner_busy;
  wire   n1761, n1762, N622, N623, N624, N625, N626, N627, N628, n5, n8, n9,
         n11, n12, n13, n14, n15, n16, n20, n24, n26, n28, n30, n32, n36, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n400, n401, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n439, n440, n441, n442,
         n445, n446, n447, n457, n458, n459, n460, n470, n488, n489, n490,
         n491, n492, n493, N9, N8, N7, N67, N66, N65, N64, N63, N62, N61, N60,
         N6, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N5, N49, N48,
         N47, N46, N45, N44, N43, N42, N41, N40, N4, N39, N38, N37, N36, N35,
         N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21,
         N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, n676, n677,
         n678, n1188, n1195, n1196, n1199, n1553, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760;
  wire   [31:0] R14;
  wire   [31:0] sigma0;
  wire   [31:0] R1;
  wire   [31:0] sigma1;
  wire   [31:0] R15;
  wire   [31:0] R6;
  wire   [31:0] logic_result;
  wire   [6:0] counter;
  wire   [31:0] R2;
  wire   [31:0] R3;
  wire   [31:0] R4;
  wire   [31:0] R5;
  wire   [31:0] R7;
  wire   [31:0] R8;
  wire   [31:0] R9;
  wire   [31:0] R10;
  wire   [31:0] R11;
  wire   [31:0] R12;
  wire   [31:0] R13;

  DFFTRX4 R1_reg_18_ ( .D(Wt[18]), .RN(n1661), .CK(clk), .Q(R1[18]), .QN(n15)
         );
  DFFTRX4 R1_reg_17_ ( .D(Wt[17]), .RN(n1661), .CK(clk), .Q(R1[17]), .QN(n14)
         );
  DFFTRX4 R14_reg_18_ ( .D(R13[18]), .RN(n1661), .CK(clk), .Q(R14[18]), .QN(n8) );
  DFFHQX4 Wt_reg_15_ ( .D(n1744), .CK(clk), .Q(Wt[15]) );
  DFFHQX4 Wt_reg_14_ ( .D(n1743), .CK(clk), .Q(Wt[14]) );
  DFFHQX4 Wt_reg_13_ ( .D(n1742), .CK(clk), .Q(Wt[13]) );
  DFFHQX4 Wt_reg_12_ ( .D(n1741), .CK(clk), .Q(Wt[12]) );
  DFFHQX4 Wt_reg_11_ ( .D(n1740), .CK(clk), .Q(Wt[11]) );
  DFFHQX4 Wt_reg_10_ ( .D(n1739), .CK(clk), .Q(Wt[10]) );
  DFFHQX4 Wt_reg_0_ ( .D(n1729), .CK(clk), .Q(n1762) );
  DFFHQX4 Wt_reg_2_ ( .D(n1731), .CK(clk), .Q(Wt[2]) );
  DFFHQX4 Wt_reg_8_ ( .D(n1737), .CK(clk), .Q(Wt[8]) );
  DFFHQX4 Wt_reg_9_ ( .D(n1738), .CK(clk), .Q(Wt[9]) );
  DFFHQX4 Wt_reg_7_ ( .D(n1736), .CK(clk), .Q(Wt[7]) );
  DFFHQX4 Wt_reg_6_ ( .D(n1735), .CK(clk), .Q(Wt[6]) );
  DFFHQX4 Wt_reg_5_ ( .D(n1734), .CK(clk), .Q(Wt[5]) );
  DFFHQX4 Wt_reg_4_ ( .D(n1733), .CK(clk), .Q(Wt[4]) );
  DFFTRX4 R14_reg_3_ ( .D(R13[3]), .RN(n1629), .CK(clk), .Q(R14[3]), .QN(n20)
         );
  DFFTRX4 R1_reg_19_ ( .D(Wt[19]), .RN(n1629), .CK(clk), .Q(R1[19]), .QN(n12)
         );
  DFFTRX4 R14_reg_5_ ( .D(R13[5]), .RN(n1630), .CK(clk), .Q(R14[5]), .QN(n11)
         );
  DFFTRX4 R14_reg_4_ ( .D(R13[4]), .RN(n1660), .CK(clk), .Q(R14[4]), .QN(n9)
         );
  DFFTRX4 R14_reg_7_ ( .D(R13[7]), .RN(n1660), .CK(clk), .Q(R14[7]) );
  DFFTRX4 R14_reg_19_ ( .D(R13[19]), .RN(n1660), .CK(clk), .Q(R14[19]) );
  DFFHQX4 Wt_reg_3_ ( .D(n1732), .CK(clk), .Q(Wt[3]) );
  DFFHQX4 Wt_reg_1_ ( .D(n1730), .CK(clk), .Q(n1761) );
  message_schedule_DW01_inc_0 add_110 ( .A(counter), .SUM({N628, N627, N626, 
        N625, N624, N623, N622}) );
  message_schedule_DW01_add_2 add_2_root_add_0_root_add_34_3 ( .A(R15), .B(R6), 
        .SUM({N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, 
        N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, 
        N40, N39, N38, N37, N36}) );
  message_schedule_DW01_add_1 add_1_root_add_0_root_add_34_3 ( .A(sigma1), .B(
        sigma0), .SUM({N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4}) );
  message_schedule_DW01_add_0 add_0_root_add_0_root_add_34_3 ( .A({N67, N66, 
        N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, 
        N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, 
        N37, N36}), .B({N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4}), .SUM(logic_result) );
  DFFTRX1 R15_reg_30_ ( .D(R14[30]), .RN(n1626), .CK(clk), .Q(R15[30]) );
  DFFTRX1 R15_reg_31_ ( .D(R14[31]), .RN(n1625), .CK(clk), .Q(R15[31]) );
  DFFTRX1 R6_reg_30_ ( .D(R5[30]), .RN(n1630), .CK(clk), .Q(R6[30]) );
  DFFTRX1 R6_reg_29_ ( .D(R5[29]), .RN(n1626), .CK(clk), .Q(R6[29]) );
  DFFTRX1 R6_reg_31_ ( .D(R5[31]), .RN(n1624), .CK(clk), .Q(R6[31]) );
  DFFTRX1 R15_reg_29_ ( .D(R14[29]), .RN(n1661), .CK(clk), .Q(R15[29]) );
  DFFTRX1 R15_reg_28_ ( .D(R14[28]), .RN(n1627), .CK(clk), .Q(R15[28]) );
  DFFTRX1 R15_reg_27_ ( .D(R14[27]), .RN(n1624), .CK(clk), .Q(R15[27]) );
  DFFTRX1 R15_reg_26_ ( .D(R14[26]), .RN(n1624), .CK(clk), .Q(R15[26]) );
  DFFTRX1 R6_reg_28_ ( .D(R5[28]), .RN(n1624), .CK(clk), .Q(R6[28]) );
  DFFTRX1 R6_reg_27_ ( .D(R5[27]), .RN(n1624), .CK(clk), .Q(R6[27]) );
  DFFTRX1 R6_reg_26_ ( .D(R5[26]), .RN(n1624), .CK(clk), .Q(R6[26]) );
  DFFTRX1 counter_reg_6_ ( .D(N628), .RN(n1624), .CK(clk), .Q(counter[6]) );
  DFFTRX1 R15_reg_25_ ( .D(R14[25]), .RN(n1624), .CK(clk), .Q(R15[25]) );
  DFFTRX1 R15_reg_24_ ( .D(R14[24]), .RN(n1624), .CK(clk), .Q(R15[24]) );
  DFFTRX1 R15_reg_23_ ( .D(R14[23]), .RN(n1624), .CK(clk), .Q(R15[23]) );
  DFFTRX1 R15_reg_22_ ( .D(R14[22]), .RN(n1625), .CK(clk), .Q(R15[22]) );
  DFFTRX1 R6_reg_25_ ( .D(R5[25]), .RN(n1624), .CK(clk), .Q(R6[25]) );
  DFFTRX1 R6_reg_24_ ( .D(R5[24]), .RN(n1624), .CK(clk), .Q(R6[24]) );
  DFFTRX1 R6_reg_23_ ( .D(R5[23]), .RN(n1625), .CK(clk), .Q(R6[23]) );
  DFFTRX1 R6_reg_22_ ( .D(R5[22]), .RN(n1625), .CK(clk), .Q(R6[22]) );
  DFFHQXL Wt_reg_31_ ( .D(n1760), .CK(clk), .Q(Wt[31]) );
  DFFHQXL Wt_reg_30_ ( .D(n1759), .CK(clk), .Q(Wt[30]) );
  DFFTRX1 R15_reg_21_ ( .D(R14[21]), .RN(n1625), .CK(clk), .Q(R15[21]) );
  DFFTRX1 R15_reg_20_ ( .D(R14[20]), .RN(n1625), .CK(clk), .Q(R15[20]) );
  DFFTRX1 R15_reg_19_ ( .D(R14[19]), .RN(n1625), .CK(clk), .Q(R15[19]) );
  DFFTRX1 R15_reg_18_ ( .D(R14[18]), .RN(n1625), .CK(clk), .Q(R15[18]) );
  DFFTRX1 R6_reg_21_ ( .D(R5[21]), .RN(n1625), .CK(clk), .Q(R6[21]) );
  DFFTRX1 R6_reg_20_ ( .D(R5[20]), .RN(n1625), .CK(clk), .Q(R6[20]) );
  DFFTRX1 R6_reg_19_ ( .D(R5[19]), .RN(n1627), .CK(clk), .Q(R6[19]) );
  DFFTRX1 R6_reg_18_ ( .D(R5[18]), .RN(n1625), .CK(clk), .Q(R6[18]) );
  DFFHQXL Wt_reg_28_ ( .D(n1757), .CK(clk), .Q(Wt[28]) );
  DFFHQXL Wt_reg_29_ ( .D(n1758), .CK(clk), .Q(Wt[29]) );
  DFFHQXL Wt_reg_27_ ( .D(n1756), .CK(clk), .Q(Wt[27]) );
  DFFTRX1 R15_reg_17_ ( .D(R14[17]), .RN(n1625), .CK(clk), .Q(R15[17]) );
  DFFTRX1 R15_reg_16_ ( .D(R14[16]), .RN(n1625), .CK(clk), .Q(R15[16]) );
  DFFTRX1 R15_reg_15_ ( .D(R14[15]), .RN(n1628), .CK(clk), .Q(R15[15]) );
  DFFTRX1 R6_reg_17_ ( .D(R5[17]), .RN(n1630), .CK(clk), .Q(R6[17]) );
  DFFTRX1 R6_reg_16_ ( .D(R5[16]), .RN(n1661), .CK(clk), .Q(R6[16]) );
  DFFTRX1 R6_reg_15_ ( .D(R5[15]), .RN(n1624), .CK(clk), .Q(R6[15]) );
  DFFHQXL Wt_reg_26_ ( .D(n1755), .CK(clk), .Q(Wt[26]) );
  DFFTRX1 R15_reg_14_ ( .D(R14[14]), .RN(n1627), .CK(clk), .Q(R15[14]) );
  DFFTRX1 R15_reg_13_ ( .D(R14[13]), .RN(n1625), .CK(clk), .Q(R15[13]) );
  DFFTRX1 R15_reg_12_ ( .D(R14[12]), .RN(n1626), .CK(clk), .Q(R15[12]) );
  DFFTRX1 R15_reg_11_ ( .D(R14[11]), .RN(n1627), .CK(clk), .Q(R15[11]) );
  DFFTRX1 R6_reg_14_ ( .D(R5[14]), .RN(n1626), .CK(clk), .Q(R6[14]) );
  DFFTRX1 R6_reg_13_ ( .D(R5[13]), .RN(n1626), .CK(clk), .Q(R6[13]) );
  DFFTRX1 R6_reg_12_ ( .D(R5[12]), .RN(n1626), .CK(clk), .Q(R6[12]) );
  DFFTRX1 R6_reg_11_ ( .D(R5[11]), .RN(n1626), .CK(clk), .Q(R6[11]) );
  DFFTRX1 R1_reg_4_ ( .D(Wt[4]), .RN(n1626), .CK(clk), .Q(R1[4]) );
  DFFTRX1 R15_reg_10_ ( .D(R14[10]), .RN(n1627), .CK(clk), .Q(R15[10]) );
  DFFTRX1 R15_reg_9_ ( .D(R14[9]), .RN(n1627), .CK(clk), .Q(R15[9]) );
  DFFTRX1 R15_reg_8_ ( .D(n1675), .RN(n1627), .CK(clk), .Q(R15[8]) );
  DFFTRX1 R15_reg_7_ ( .D(R14[7]), .RN(n1627), .CK(clk), .Q(R15[7]) );
  DFFTRX1 R6_reg_10_ ( .D(R5[10]), .RN(n1627), .CK(clk), .Q(R6[10]) );
  DFFTRX1 R6_reg_9_ ( .D(R5[9]), .RN(n1627), .CK(clk), .Q(R6[9]) );
  DFFTRX1 R6_reg_8_ ( .D(R5[8]), .RN(n1627), .CK(clk), .Q(R6[8]) );
  DFFTRX1 R6_reg_7_ ( .D(R5[7]), .RN(n1627), .CK(clk), .Q(R6[7]) );
  DFFTRX1 R15_reg_5_ ( .D(R14[5]), .RN(n1626), .CK(clk), .Q(R15[5]) );
  DFFTRX1 R15_reg_3_ ( .D(R14[3]), .RN(n1661), .CK(clk), .Q(R15[3]) );
  DFFTRX1 R15_reg_1_ ( .D(R14[1]), .RN(n1660), .CK(clk), .Q(R15[1]) );
  DFFTRX1 R15_reg_2_ ( .D(R14[2]), .RN(n1629), .CK(clk), .Q(R15[2]) );
  DFFTRX1 R14_reg_22_ ( .D(R13[22]), .RN(n1630), .CK(clk), .Q(R14[22]), .QN(
        n408) );
  DFFTRX1 R14_reg_20_ ( .D(R13[20]), .RN(n1630), .CK(clk), .Q(R14[20]), .QN(
        n395) );
  DFFTRX1 R14_reg_13_ ( .D(R13[13]), .RN(n1628), .CK(clk), .Q(R14[13]), .QN(
        n32) );
  DFFTRX1 R14_reg_11_ ( .D(R13[11]), .RN(n1630), .CK(clk), .Q(R14[11]), .QN(
        n28) );
  DFFTRX1 R14_reg_12_ ( .D(R13[12]), .RN(n1628), .CK(clk), .Q(R14[12]), .QN(
        n412) );
  DFFTRX1 R6_reg_6_ ( .D(R5[6]), .RN(n1628), .CK(clk), .Q(R6[6]) );
  DFFTRX1 R6_reg_5_ ( .D(R5[5]), .RN(n1628), .CK(clk), .Q(R6[5]) );
  DFFTRX1 R6_reg_4_ ( .D(R5[4]), .RN(n1628), .CK(clk), .Q(R6[4]) );
  DFFTRX1 R6_reg_3_ ( .D(R5[3]), .RN(n1628), .CK(clk), .Q(R6[3]) );
  DFFTRX1 R6_reg_1_ ( .D(R5[1]), .RN(n1660), .CK(clk), .Q(R6[1]) );
  DFFTRX1 R1_reg_27_ ( .D(Wt[27]), .RN(n1629), .CK(clk), .Q(R1[27]), .QN(n411)
         );
  DFFTRX1 R14_reg_26_ ( .D(R13[26]), .RN(n1628), .CK(clk), .Q(R14[26]), .QN(
        n410) );
  DFFHQX1 Wt_reg_18_ ( .D(n1747), .CK(clk), .Q(Wt[18]) );
  DFFTRX1 R14_reg_14_ ( .D(R13[14]), .RN(n1629), .CK(clk), .Q(R14[14]), .QN(
        n404) );
  DFFTRX1 R14_reg_25_ ( .D(R13[25]), .RN(n1629), .CK(clk), .Q(R14[25]), .QN(
        n409) );
  DFFHQX1 Wt_reg_17_ ( .D(n1746), .CK(clk), .Q(Wt[17]) );
  DFFTRX1 R14_reg_15_ ( .D(R13[15]), .RN(n1629), .CK(clk), .Q(R14[15]), .QN(
        n30) );
  DFFTRX1 R10_reg_4_ ( .D(R9[4]), .RN(n1656), .CK(clk), .Q(R10[4]) );
  DFFTRX1 R11_reg_4_ ( .D(R10[4]), .RN(n1656), .CK(clk), .Q(R11[4]) );
  DFFTRX1 R12_reg_4_ ( .D(R11[4]), .RN(n1656), .CK(clk), .Q(R12[4]) );
  DFFTRX1 R13_reg_4_ ( .D(R12[4]), .RN(n1656), .CK(clk), .Q(R13[4]) );
  DFFTRX1 R2_reg_3_ ( .D(R1[3]), .RN(n1656), .CK(clk), .Q(R2[3]) );
  DFFTRX1 R3_reg_3_ ( .D(R2[3]), .RN(n1656), .CK(clk), .Q(R3[3]) );
  DFFTRX1 R4_reg_3_ ( .D(R3[3]), .RN(n1656), .CK(clk), .Q(R4[3]) );
  DFFTRX1 R5_reg_3_ ( .D(R4[3]), .RN(n1656), .CK(clk), .Q(R5[3]) );
  DFFTRX1 R7_reg_3_ ( .D(R6[3]), .RN(n1656), .CK(clk), .Q(R7[3]) );
  DFFTRX1 R8_reg_3_ ( .D(R7[3]), .RN(n1656), .CK(clk), .Q(R8[3]) );
  DFFTRX1 R9_reg_3_ ( .D(R8[3]), .RN(n1656), .CK(clk), .Q(R9[3]) );
  DFFTRX1 R10_reg_3_ ( .D(R9[3]), .RN(n1656), .CK(clk), .Q(R10[3]) );
  DFFTRX1 R11_reg_3_ ( .D(R10[3]), .RN(n1657), .CK(clk), .Q(R11[3]) );
  DFFTRX1 R12_reg_3_ ( .D(R11[3]), .RN(n1657), .CK(clk), .Q(R12[3]) );
  DFFTRX1 R13_reg_3_ ( .D(R12[3]), .RN(n1657), .CK(clk), .Q(R13[3]) );
  DFFTRX1 R2_reg_2_ ( .D(R1[2]), .RN(n1657), .CK(clk), .Q(R2[2]) );
  DFFTRX1 R3_reg_2_ ( .D(R2[2]), .RN(n1657), .CK(clk), .Q(R3[2]) );
  DFFTRX1 R4_reg_2_ ( .D(R3[2]), .RN(n1657), .CK(clk), .Q(R4[2]) );
  DFFTRX1 R5_reg_2_ ( .D(R4[2]), .RN(n1657), .CK(clk), .Q(R5[2]) );
  DFFTRX1 R7_reg_2_ ( .D(R6[2]), .RN(n1657), .CK(clk), .Q(R7[2]) );
  DFFTRX1 R8_reg_2_ ( .D(R7[2]), .RN(n1657), .CK(clk), .Q(R8[2]) );
  DFFTRX1 R9_reg_2_ ( .D(R8[2]), .RN(n1657), .CK(clk), .Q(R9[2]) );
  DFFTRX1 R10_reg_2_ ( .D(R9[2]), .RN(n1657), .CK(clk), .Q(R10[2]) );
  DFFTRX1 R11_reg_2_ ( .D(R10[2]), .RN(n1657), .CK(clk), .Q(R11[2]) );
  DFFTRX1 R12_reg_2_ ( .D(R11[2]), .RN(n1658), .CK(clk), .Q(R12[2]) );
  DFFTRX1 R13_reg_2_ ( .D(R12[2]), .RN(n1658), .CK(clk), .Q(R13[2]) );
  DFFTRX1 R2_reg_1_ ( .D(R1[1]), .RN(n1658), .CK(clk), .Q(R2[1]) );
  DFFTRX1 R3_reg_1_ ( .D(R2[1]), .RN(n1658), .CK(clk), .Q(R3[1]) );
  DFFTRX1 R4_reg_1_ ( .D(R3[1]), .RN(n1658), .CK(clk), .Q(R4[1]) );
  DFFTRX1 R5_reg_1_ ( .D(R4[1]), .RN(n1658), .CK(clk), .Q(R5[1]) );
  DFFTRX1 R7_reg_1_ ( .D(R6[1]), .RN(n1658), .CK(clk), .Q(R7[1]) );
  DFFTRX1 R8_reg_1_ ( .D(R7[1]), .RN(n1658), .CK(clk), .Q(R8[1]) );
  DFFTRX1 R9_reg_1_ ( .D(R8[1]), .RN(n1658), .CK(clk), .Q(R9[1]) );
  DFFTRX1 R10_reg_1_ ( .D(R9[1]), .RN(n1658), .CK(clk), .Q(R10[1]) );
  DFFTRX1 R11_reg_1_ ( .D(R10[1]), .RN(n1658), .CK(clk), .Q(R11[1]) );
  DFFTRX1 R12_reg_1_ ( .D(R11[1]), .RN(n1658), .CK(clk), .Q(R12[1]) );
  DFFTRX1 R13_reg_1_ ( .D(R12[1]), .RN(n1659), .CK(clk), .Q(R13[1]) );
  DFFTRX1 R2_reg_0_ ( .D(R1[0]), .RN(n1659), .CK(clk), .Q(R2[0]) );
  DFFTRX1 R3_reg_0_ ( .D(R2[0]), .RN(n1659), .CK(clk), .Q(R3[0]) );
  DFFTRX1 R4_reg_0_ ( .D(R3[0]), .RN(n1659), .CK(clk), .Q(R4[0]) );
  DFFTRX1 R5_reg_0_ ( .D(R4[0]), .RN(n1659), .CK(clk), .Q(R5[0]) );
  DFFTRX1 R7_reg_0_ ( .D(R6[0]), .RN(n1659), .CK(clk), .Q(R7[0]) );
  DFFTRX1 R8_reg_0_ ( .D(R7[0]), .RN(n1659), .CK(clk), .Q(R8[0]) );
  DFFTRX1 R9_reg_0_ ( .D(R8[0]), .RN(n1659), .CK(clk), .Q(R9[0]) );
  DFFTRX1 R10_reg_0_ ( .D(R9[0]), .RN(n1659), .CK(clk), .Q(R10[0]) );
  DFFTRX1 R11_reg_0_ ( .D(R10[0]), .RN(n1659), .CK(clk), .Q(R11[0]) );
  DFFTRX1 R12_reg_0_ ( .D(R11[0]), .RN(n1659), .CK(clk), .Q(R12[0]) );
  DFFTRX1 R13_reg_0_ ( .D(R12[0]), .RN(n1659), .CK(clk), .Q(R13[0]) );
  DFFTRX1 R13_reg_8_ ( .D(R12[8]), .RN(n1660), .CK(clk), .Q(R13[8]) );
  DFFTRX1 R13_reg_31_ ( .D(R12[31]), .RN(n1630), .CK(clk), .Q(R13[31]) );
  DFFTRX1 R2_reg_30_ ( .D(R1[30]), .RN(n1630), .CK(clk), .Q(R2[30]) );
  DFFTRX1 R3_reg_30_ ( .D(R2[30]), .RN(n1630), .CK(clk), .Q(R3[30]) );
  DFFTRX1 R4_reg_30_ ( .D(R3[30]), .RN(n1631), .CK(clk), .Q(R4[30]) );
  DFFTRX1 R5_reg_30_ ( .D(R4[30]), .RN(n1631), .CK(clk), .Q(R5[30]) );
  DFFTRX1 R7_reg_30_ ( .D(R6[30]), .RN(n1631), .CK(clk), .Q(R7[30]) );
  DFFTRX1 R8_reg_30_ ( .D(R7[30]), .RN(n1631), .CK(clk), .Q(R8[30]) );
  DFFTRX1 R9_reg_30_ ( .D(R8[30]), .RN(n1631), .CK(clk), .Q(R9[30]) );
  DFFTRX1 R10_reg_30_ ( .D(R9[30]), .RN(n1631), .CK(clk), .Q(R10[30]) );
  DFFTRX1 R11_reg_30_ ( .D(R10[30]), .RN(n1631), .CK(clk), .Q(R11[30]) );
  DFFTRX1 R12_reg_30_ ( .D(R11[30]), .RN(n1631), .CK(clk), .Q(R12[30]) );
  DFFTRX1 R13_reg_30_ ( .D(R12[30]), .RN(n1631), .CK(clk), .Q(R13[30]) );
  DFFTRX1 R2_reg_29_ ( .D(R1[29]), .RN(n1631), .CK(clk), .Q(R2[29]) );
  DFFTRX1 R3_reg_29_ ( .D(R2[29]), .RN(n1631), .CK(clk), .Q(R3[29]) );
  DFFTRX1 R2_reg_31_ ( .D(R1[31]), .RN(n1631), .CK(clk), .Q(R2[31]) );
  DFFTRX1 R3_reg_31_ ( .D(R2[31]), .RN(n1632), .CK(clk), .Q(R3[31]) );
  DFFTRX1 R4_reg_31_ ( .D(R3[31]), .RN(n1632), .CK(clk), .Q(R4[31]) );
  DFFTRX1 R5_reg_31_ ( .D(R4[31]), .RN(n1632), .CK(clk), .Q(R5[31]) );
  DFFTRX1 R7_reg_31_ ( .D(R6[31]), .RN(n1632), .CK(clk), .Q(R7[31]) );
  DFFTRX1 R8_reg_31_ ( .D(R7[31]), .RN(n1632), .CK(clk), .Q(R8[31]) );
  DFFTRX1 R9_reg_31_ ( .D(R8[31]), .RN(n1632), .CK(clk), .Q(R9[31]) );
  DFFTRX1 R10_reg_31_ ( .D(R9[31]), .RN(n1632), .CK(clk), .Q(R10[31]) );
  DFFTRX1 R11_reg_31_ ( .D(R10[31]), .RN(n1632), .CK(clk), .Q(R11[31]) );
  DFFTRX1 R12_reg_31_ ( .D(R11[31]), .RN(n1632), .CK(clk), .Q(R12[31]) );
  DFFTRX1 R4_reg_29_ ( .D(R3[29]), .RN(n1632), .CK(clk), .Q(R4[29]) );
  DFFTRX1 R5_reg_29_ ( .D(R4[29]), .RN(n1632), .CK(clk), .Q(R5[29]) );
  DFFTRX1 R7_reg_29_ ( .D(R6[29]), .RN(n1632), .CK(clk), .Q(R7[29]) );
  DFFTRX1 R8_reg_29_ ( .D(R7[29]), .RN(n1633), .CK(clk), .Q(R8[29]) );
  DFFTRX1 R9_reg_29_ ( .D(R8[29]), .RN(n1633), .CK(clk), .Q(R9[29]) );
  DFFTRX1 R10_reg_29_ ( .D(R9[29]), .RN(n1633), .CK(clk), .Q(R10[29]) );
  DFFTRX1 R11_reg_29_ ( .D(R10[29]), .RN(n1633), .CK(clk), .Q(R11[29]) );
  DFFTRX1 R12_reg_29_ ( .D(R11[29]), .RN(n1633), .CK(clk), .Q(R12[29]) );
  DFFTRX1 R13_reg_29_ ( .D(R12[29]), .RN(n1633), .CK(clk), .Q(R13[29]) );
  DFFTRX1 R2_reg_28_ ( .D(R1[28]), .RN(n1633), .CK(clk), .Q(R2[28]) );
  DFFTRX1 R3_reg_28_ ( .D(R2[28]), .RN(n1633), .CK(clk), .Q(R3[28]) );
  DFFTRX1 R4_reg_28_ ( .D(R3[28]), .RN(n1633), .CK(clk), .Q(R4[28]) );
  DFFTRX1 R5_reg_28_ ( .D(R4[28]), .RN(n1633), .CK(clk), .Q(R5[28]) );
  DFFTRX1 R7_reg_28_ ( .D(R6[28]), .RN(n1633), .CK(clk), .Q(R7[28]) );
  DFFTRX1 R8_reg_28_ ( .D(R7[28]), .RN(n1633), .CK(clk), .Q(R8[28]) );
  DFFTRX1 R9_reg_28_ ( .D(R8[28]), .RN(n1634), .CK(clk), .Q(R9[28]) );
  DFFTRX1 R10_reg_28_ ( .D(R9[28]), .RN(n1634), .CK(clk), .Q(R10[28]) );
  DFFTRX1 R11_reg_28_ ( .D(R10[28]), .RN(n1634), .CK(clk), .Q(R11[28]) );
  DFFTRX1 R12_reg_28_ ( .D(R11[28]), .RN(n1634), .CK(clk), .Q(R12[28]) );
  DFFTRX1 R13_reg_28_ ( .D(R12[28]), .RN(n1634), .CK(clk), .Q(R13[28]) );
  DFFTRX1 R2_reg_27_ ( .D(R1[27]), .RN(n1634), .CK(clk), .Q(R2[27]) );
  DFFTRX1 R3_reg_27_ ( .D(R2[27]), .RN(n1634), .CK(clk), .Q(R3[27]) );
  DFFTRX1 R4_reg_27_ ( .D(R3[27]), .RN(n1634), .CK(clk), .Q(R4[27]) );
  DFFTRX1 R5_reg_27_ ( .D(R4[27]), .RN(n1634), .CK(clk), .Q(R5[27]) );
  DFFTRX1 R7_reg_27_ ( .D(R6[27]), .RN(n1634), .CK(clk), .Q(R7[27]) );
  DFFTRX1 R8_reg_27_ ( .D(R7[27]), .RN(n1634), .CK(clk), .Q(R8[27]) );
  DFFTRX1 R9_reg_27_ ( .D(R8[27]), .RN(n1634), .CK(clk), .Q(R9[27]) );
  DFFTRX1 R10_reg_27_ ( .D(R9[27]), .RN(n1635), .CK(clk), .Q(R10[27]) );
  DFFTRX1 R11_reg_27_ ( .D(R10[27]), .RN(n1635), .CK(clk), .Q(R11[27]) );
  DFFTRX1 R12_reg_27_ ( .D(R11[27]), .RN(n1635), .CK(clk), .Q(R12[27]) );
  DFFTRX1 R13_reg_27_ ( .D(R12[27]), .RN(n1635), .CK(clk), .Q(R13[27]) );
  DFFTRX1 R2_reg_26_ ( .D(R1[26]), .RN(n1635), .CK(clk), .Q(R2[26]) );
  DFFTRX1 R3_reg_26_ ( .D(R2[26]), .RN(n1635), .CK(clk), .Q(R3[26]) );
  DFFTRX1 R4_reg_26_ ( .D(R3[26]), .RN(n1635), .CK(clk), .Q(R4[26]) );
  DFFTRX1 R5_reg_26_ ( .D(R4[26]), .RN(n1635), .CK(clk), .Q(R5[26]) );
  DFFTRX1 R7_reg_26_ ( .D(R6[26]), .RN(n1635), .CK(clk), .Q(R7[26]) );
  DFFTRX1 R8_reg_26_ ( .D(R7[26]), .RN(n1635), .CK(clk), .Q(R8[26]) );
  DFFTRX1 R9_reg_26_ ( .D(R8[26]), .RN(n1635), .CK(clk), .Q(R9[26]) );
  DFFTRX1 R10_reg_26_ ( .D(R9[26]), .RN(n1635), .CK(clk), .Q(R10[26]) );
  DFFTRX1 R11_reg_26_ ( .D(R10[26]), .RN(n1636), .CK(clk), .Q(R11[26]) );
  DFFTRX1 R12_reg_26_ ( .D(R11[26]), .RN(n1636), .CK(clk), .Q(R12[26]) );
  DFFTRX1 R13_reg_26_ ( .D(R12[26]), .RN(n1636), .CK(clk), .Q(R13[26]) );
  DFFTRX1 R2_reg_25_ ( .D(R1[25]), .RN(n1636), .CK(clk), .Q(R2[25]) );
  DFFTRX1 R3_reg_25_ ( .D(R2[25]), .RN(n1636), .CK(clk), .Q(R3[25]) );
  DFFTRX1 R4_reg_25_ ( .D(R3[25]), .RN(n1636), .CK(clk), .Q(R4[25]) );
  DFFTRX1 R5_reg_25_ ( .D(R4[25]), .RN(n1636), .CK(clk), .Q(R5[25]) );
  DFFTRX1 R7_reg_25_ ( .D(R6[25]), .RN(n1636), .CK(clk), .Q(R7[25]) );
  DFFTRX1 R8_reg_25_ ( .D(R7[25]), .RN(n1636), .CK(clk), .Q(R8[25]) );
  DFFTRX1 R9_reg_25_ ( .D(R8[25]), .RN(n1636), .CK(clk), .Q(R9[25]) );
  DFFTRX1 R10_reg_25_ ( .D(R9[25]), .RN(n1636), .CK(clk), .Q(R10[25]) );
  DFFTRX1 R11_reg_25_ ( .D(R10[25]), .RN(n1636), .CK(clk), .Q(R11[25]) );
  DFFTRX1 R12_reg_25_ ( .D(R11[25]), .RN(n1637), .CK(clk), .Q(R12[25]) );
  DFFTRX1 R13_reg_25_ ( .D(R12[25]), .RN(n1637), .CK(clk), .Q(R13[25]) );
  DFFTRX1 R2_reg_24_ ( .D(R1[24]), .RN(n1637), .CK(clk), .Q(R2[24]) );
  DFFTRX1 R3_reg_24_ ( .D(R2[24]), .RN(n1637), .CK(clk), .Q(R3[24]) );
  DFFTRX1 R4_reg_24_ ( .D(R3[24]), .RN(n1637), .CK(clk), .Q(R4[24]) );
  DFFTRX1 R5_reg_24_ ( .D(R4[24]), .RN(n1637), .CK(clk), .Q(R5[24]) );
  DFFTRX1 R7_reg_24_ ( .D(R6[24]), .RN(n1637), .CK(clk), .Q(R7[24]) );
  DFFTRX1 R8_reg_24_ ( .D(R7[24]), .RN(n1637), .CK(clk), .Q(R8[24]) );
  DFFTRX1 R9_reg_24_ ( .D(R8[24]), .RN(n1637), .CK(clk), .Q(R9[24]) );
  DFFTRX1 R10_reg_24_ ( .D(R9[24]), .RN(n1637), .CK(clk), .Q(R10[24]) );
  DFFTRX1 R11_reg_24_ ( .D(R10[24]), .RN(n1637), .CK(clk), .Q(R11[24]) );
  DFFTRX1 R12_reg_24_ ( .D(R11[24]), .RN(n1637), .CK(clk), .Q(R12[24]) );
  DFFTRX1 R13_reg_24_ ( .D(R12[24]), .RN(n1638), .CK(clk), .Q(R13[24]) );
  DFFTRX1 R2_reg_23_ ( .D(R1[23]), .RN(n1638), .CK(clk), .Q(R2[23]) );
  DFFTRX1 R3_reg_23_ ( .D(R2[23]), .RN(n1638), .CK(clk), .Q(R3[23]) );
  DFFTRX1 R4_reg_23_ ( .D(R3[23]), .RN(n1638), .CK(clk), .Q(R4[23]) );
  DFFTRX1 R5_reg_23_ ( .D(R4[23]), .RN(n1638), .CK(clk), .Q(R5[23]) );
  DFFTRX1 R7_reg_23_ ( .D(R6[23]), .RN(n1638), .CK(clk), .Q(R7[23]) );
  DFFTRX1 R8_reg_23_ ( .D(R7[23]), .RN(n1638), .CK(clk), .Q(R8[23]) );
  DFFTRX1 R9_reg_23_ ( .D(R8[23]), .RN(n1638), .CK(clk), .Q(R9[23]) );
  DFFTRX1 R10_reg_23_ ( .D(R9[23]), .RN(n1638), .CK(clk), .Q(R10[23]) );
  DFFTRX1 R11_reg_23_ ( .D(R10[23]), .RN(n1638), .CK(clk), .Q(R11[23]) );
  DFFTRX1 R12_reg_23_ ( .D(R11[23]), .RN(n1638), .CK(clk), .Q(R12[23]) );
  DFFTRX1 R13_reg_23_ ( .D(R12[23]), .RN(n1638), .CK(clk), .Q(R13[23]) );
  DFFTRX1 R2_reg_22_ ( .D(R1[22]), .RN(n1639), .CK(clk), .Q(R2[22]) );
  DFFTRX1 R3_reg_22_ ( .D(R2[22]), .RN(n1639), .CK(clk), .Q(R3[22]) );
  DFFTRX1 R4_reg_22_ ( .D(R3[22]), .RN(n1639), .CK(clk), .Q(R4[22]) );
  DFFTRX1 R5_reg_22_ ( .D(R4[22]), .RN(n1639), .CK(clk), .Q(R5[22]) );
  DFFTRX1 R7_reg_22_ ( .D(R6[22]), .RN(n1639), .CK(clk), .Q(R7[22]) );
  DFFTRX1 R8_reg_22_ ( .D(R7[22]), .RN(n1639), .CK(clk), .Q(R8[22]) );
  DFFTRX1 R9_reg_22_ ( .D(R8[22]), .RN(n1639), .CK(clk), .Q(R9[22]) );
  DFFTRX1 R10_reg_22_ ( .D(R9[22]), .RN(n1639), .CK(clk), .Q(R10[22]) );
  DFFTRX1 R11_reg_22_ ( .D(R10[22]), .RN(n1639), .CK(clk), .Q(R11[22]) );
  DFFTRX1 R12_reg_22_ ( .D(R11[22]), .RN(n1639), .CK(clk), .Q(R12[22]) );
  DFFTRX1 R13_reg_22_ ( .D(R12[22]), .RN(n1639), .CK(clk), .Q(R13[22]) );
  DFFTRX1 R2_reg_21_ ( .D(R1[21]), .RN(n1639), .CK(clk), .Q(R2[21]) );
  DFFTRX1 R3_reg_21_ ( .D(R2[21]), .RN(n1640), .CK(clk), .Q(R3[21]) );
  DFFTRX1 R4_reg_21_ ( .D(R3[21]), .RN(n1640), .CK(clk), .Q(R4[21]) );
  DFFTRX1 R5_reg_21_ ( .D(R4[21]), .RN(n1640), .CK(clk), .Q(R5[21]) );
  DFFTRX1 R7_reg_21_ ( .D(R6[21]), .RN(n1640), .CK(clk), .Q(R7[21]) );
  DFFTRX1 R8_reg_21_ ( .D(R7[21]), .RN(n1640), .CK(clk), .Q(R8[21]) );
  DFFTRX1 R9_reg_21_ ( .D(R8[21]), .RN(n1640), .CK(clk), .Q(R9[21]) );
  DFFTRX1 R10_reg_21_ ( .D(R9[21]), .RN(n1640), .CK(clk), .Q(R10[21]) );
  DFFTRX1 R11_reg_21_ ( .D(R10[21]), .RN(n1640), .CK(clk), .Q(R11[21]) );
  DFFTRX1 R12_reg_21_ ( .D(R11[21]), .RN(n1640), .CK(clk), .Q(R12[21]) );
  DFFTRX1 R13_reg_21_ ( .D(R12[21]), .RN(n1640), .CK(clk), .Q(R13[21]) );
  DFFTRX1 R2_reg_20_ ( .D(R1[20]), .RN(n1640), .CK(clk), .Q(R2[20]) );
  DFFTRX1 R3_reg_20_ ( .D(R2[20]), .RN(n1640), .CK(clk), .Q(R3[20]) );
  DFFTRX1 R4_reg_20_ ( .D(R3[20]), .RN(n1641), .CK(clk), .Q(R4[20]) );
  DFFTRX1 R5_reg_20_ ( .D(R4[20]), .RN(n1641), .CK(clk), .Q(R5[20]) );
  DFFTRX1 R7_reg_20_ ( .D(R6[20]), .RN(n1641), .CK(clk), .Q(R7[20]) );
  DFFTRX1 R8_reg_20_ ( .D(R7[20]), .RN(n1641), .CK(clk), .Q(R8[20]) );
  DFFTRX1 R9_reg_20_ ( .D(R8[20]), .RN(n1641), .CK(clk), .Q(R9[20]) );
  DFFTRX1 R10_reg_20_ ( .D(R9[20]), .RN(n1641), .CK(clk), .Q(R10[20]) );
  DFFTRX1 R11_reg_20_ ( .D(R10[20]), .RN(n1641), .CK(clk), .Q(R11[20]) );
  DFFTRX1 R12_reg_20_ ( .D(R11[20]), .RN(n1641), .CK(clk), .Q(R12[20]) );
  DFFTRX1 R13_reg_20_ ( .D(R12[20]), .RN(n1641), .CK(clk), .Q(R13[20]) );
  DFFTRX1 R2_reg_19_ ( .D(R1[19]), .RN(n1641), .CK(clk), .Q(R2[19]) );
  DFFTRX1 R3_reg_19_ ( .D(R2[19]), .RN(n1641), .CK(clk), .Q(R3[19]) );
  DFFTRX1 R4_reg_19_ ( .D(R3[19]), .RN(n1641), .CK(clk), .Q(R4[19]) );
  DFFTRX1 R5_reg_19_ ( .D(R4[19]), .RN(n1642), .CK(clk), .Q(R5[19]) );
  DFFTRX1 R7_reg_19_ ( .D(R6[19]), .RN(n1642), .CK(clk), .Q(R7[19]) );
  DFFTRX1 R8_reg_19_ ( .D(R7[19]), .RN(n1642), .CK(clk), .Q(R8[19]) );
  DFFTRX1 R9_reg_19_ ( .D(R8[19]), .RN(n1642), .CK(clk), .Q(R9[19]) );
  DFFTRX1 R10_reg_19_ ( .D(R9[19]), .RN(n1642), .CK(clk), .Q(R10[19]) );
  DFFTRX1 R11_reg_19_ ( .D(R10[19]), .RN(n1642), .CK(clk), .Q(R11[19]) );
  DFFTRX1 R12_reg_19_ ( .D(R11[19]), .RN(n1642), .CK(clk), .Q(R12[19]) );
  DFFTRX1 R13_reg_19_ ( .D(R12[19]), .RN(n1642), .CK(clk), .Q(R13[19]) );
  DFFTRX1 R2_reg_18_ ( .D(R1[18]), .RN(n1642), .CK(clk), .Q(R2[18]) );
  DFFTRX1 R3_reg_18_ ( .D(R2[18]), .RN(n1642), .CK(clk), .Q(R3[18]) );
  DFFTRX1 R4_reg_18_ ( .D(R3[18]), .RN(n1642), .CK(clk), .Q(R4[18]) );
  DFFTRX1 R5_reg_18_ ( .D(R4[18]), .RN(n1642), .CK(clk), .Q(R5[18]) );
  DFFTRX1 R7_reg_18_ ( .D(R6[18]), .RN(n1643), .CK(clk), .Q(R7[18]) );
  DFFTRX1 R8_reg_18_ ( .D(R7[18]), .RN(n1643), .CK(clk), .Q(R8[18]) );
  DFFTRX1 R9_reg_18_ ( .D(R8[18]), .RN(n1643), .CK(clk), .Q(R9[18]) );
  DFFTRX1 R10_reg_18_ ( .D(R9[18]), .RN(n1643), .CK(clk), .Q(R10[18]) );
  DFFTRX1 R11_reg_18_ ( .D(R10[18]), .RN(n1643), .CK(clk), .Q(R11[18]) );
  DFFTRX1 R12_reg_18_ ( .D(R11[18]), .RN(n1643), .CK(clk), .Q(R12[18]) );
  DFFTRX1 R13_reg_18_ ( .D(R12[18]), .RN(n1643), .CK(clk), .Q(R13[18]) );
  DFFTRX1 R2_reg_17_ ( .D(R1[17]), .RN(n1643), .CK(clk), .Q(R2[17]) );
  DFFTRX1 R3_reg_17_ ( .D(R2[17]), .RN(n1643), .CK(clk), .Q(R3[17]) );
  DFFTRX1 R4_reg_17_ ( .D(R3[17]), .RN(n1643), .CK(clk), .Q(R4[17]) );
  DFFTRX1 R5_reg_17_ ( .D(R4[17]), .RN(n1643), .CK(clk), .Q(R5[17]) );
  DFFTRX1 R7_reg_17_ ( .D(R6[17]), .RN(n1643), .CK(clk), .Q(R7[17]) );
  DFFTRX1 R8_reg_17_ ( .D(R7[17]), .RN(n1644), .CK(clk), .Q(R8[17]) );
  DFFTRX1 R9_reg_17_ ( .D(R8[17]), .RN(n1644), .CK(clk), .Q(R9[17]) );
  DFFTRX1 R10_reg_17_ ( .D(R9[17]), .RN(n1644), .CK(clk), .Q(R10[17]) );
  DFFTRX1 R11_reg_17_ ( .D(R10[17]), .RN(n1644), .CK(clk), .Q(R11[17]) );
  DFFTRX1 R12_reg_17_ ( .D(R11[17]), .RN(n1644), .CK(clk), .Q(R12[17]) );
  DFFTRX1 R13_reg_17_ ( .D(R12[17]), .RN(n1644), .CK(clk), .Q(R13[17]) );
  DFFTRX1 R2_reg_16_ ( .D(R1[16]), .RN(n1644), .CK(clk), .Q(R2[16]) );
  DFFTRX1 R3_reg_16_ ( .D(R2[16]), .RN(n1644), .CK(clk), .Q(R3[16]) );
  DFFTRX1 R4_reg_16_ ( .D(R3[16]), .RN(n1644), .CK(clk), .Q(R4[16]) );
  DFFTRX1 R5_reg_16_ ( .D(R4[16]), .RN(n1644), .CK(clk), .Q(R5[16]) );
  DFFTRX1 R7_reg_16_ ( .D(R6[16]), .RN(n1644), .CK(clk), .Q(R7[16]) );
  DFFTRX1 R8_reg_16_ ( .D(R7[16]), .RN(n1644), .CK(clk), .Q(R8[16]) );
  DFFTRX1 R9_reg_16_ ( .D(R8[16]), .RN(n1645), .CK(clk), .Q(R9[16]) );
  DFFTRX1 R10_reg_16_ ( .D(R9[16]), .RN(n1645), .CK(clk), .Q(R10[16]) );
  DFFTRX1 R11_reg_16_ ( .D(R10[16]), .RN(n1645), .CK(clk), .Q(R11[16]) );
  DFFTRX1 R12_reg_16_ ( .D(R11[16]), .RN(n1645), .CK(clk), .Q(R12[16]) );
  DFFTRX1 R13_reg_16_ ( .D(R12[16]), .RN(n1645), .CK(clk), .Q(R13[16]) );
  DFFTRX1 R2_reg_15_ ( .D(R1[15]), .RN(n1645), .CK(clk), .Q(R2[15]) );
  DFFTRX1 R3_reg_15_ ( .D(R2[15]), .RN(n1645), .CK(clk), .Q(R3[15]) );
  DFFTRX1 R4_reg_15_ ( .D(R3[15]), .RN(n1645), .CK(clk), .Q(R4[15]) );
  DFFTRX1 R5_reg_15_ ( .D(R4[15]), .RN(n1645), .CK(clk), .Q(R5[15]) );
  DFFTRX1 R7_reg_15_ ( .D(R6[15]), .RN(n1645), .CK(clk), .Q(R7[15]) );
  DFFTRX1 R8_reg_15_ ( .D(R7[15]), .RN(n1645), .CK(clk), .Q(R8[15]) );
  DFFTRX1 R9_reg_15_ ( .D(R8[15]), .RN(n1645), .CK(clk), .Q(R9[15]) );
  DFFTRX1 R10_reg_15_ ( .D(R9[15]), .RN(n1646), .CK(clk), .Q(R10[15]) );
  DFFTRX1 R11_reg_15_ ( .D(R10[15]), .RN(n1646), .CK(clk), .Q(R11[15]) );
  DFFTRX1 R12_reg_15_ ( .D(R11[15]), .RN(n1646), .CK(clk), .Q(R12[15]) );
  DFFTRX1 R13_reg_15_ ( .D(R12[15]), .RN(n1646), .CK(clk), .Q(R13[15]) );
  DFFTRX1 R2_reg_14_ ( .D(R1[14]), .RN(n1646), .CK(clk), .Q(R2[14]) );
  DFFTRX1 R3_reg_14_ ( .D(R2[14]), .RN(n1646), .CK(clk), .Q(R3[14]) );
  DFFTRX1 R4_reg_14_ ( .D(R3[14]), .RN(n1646), .CK(clk), .Q(R4[14]) );
  DFFTRX1 R5_reg_14_ ( .D(R4[14]), .RN(n1646), .CK(clk), .Q(R5[14]) );
  DFFTRX1 R7_reg_14_ ( .D(R6[14]), .RN(n1646), .CK(clk), .Q(R7[14]) );
  DFFTRX1 R8_reg_14_ ( .D(R7[14]), .RN(n1646), .CK(clk), .Q(R8[14]) );
  DFFTRX1 R9_reg_14_ ( .D(R8[14]), .RN(n1646), .CK(clk), .Q(R9[14]) );
  DFFTRX1 R10_reg_14_ ( .D(R9[14]), .RN(n1646), .CK(clk), .Q(R10[14]) );
  DFFTRX1 R11_reg_14_ ( .D(R10[14]), .RN(n1647), .CK(clk), .Q(R11[14]) );
  DFFTRX1 R12_reg_14_ ( .D(R11[14]), .RN(n1647), .CK(clk), .Q(R12[14]) );
  DFFTRX1 R13_reg_14_ ( .D(R12[14]), .RN(n1647), .CK(clk), .Q(R13[14]) );
  DFFTRX1 R2_reg_13_ ( .D(R1[13]), .RN(n1647), .CK(clk), .Q(R2[13]) );
  DFFTRX1 R3_reg_13_ ( .D(R2[13]), .RN(n1647), .CK(clk), .Q(R3[13]) );
  DFFTRX1 R4_reg_13_ ( .D(R3[13]), .RN(n1647), .CK(clk), .Q(R4[13]) );
  DFFTRX1 R5_reg_13_ ( .D(R4[13]), .RN(n1647), .CK(clk), .Q(R5[13]) );
  DFFTRX1 R7_reg_13_ ( .D(R6[13]), .RN(n1647), .CK(clk), .Q(R7[13]) );
  DFFTRX1 R8_reg_13_ ( .D(R7[13]), .RN(n1647), .CK(clk), .Q(R8[13]) );
  DFFTRX1 R9_reg_13_ ( .D(R8[13]), .RN(n1647), .CK(clk), .Q(R9[13]) );
  DFFTRX1 R10_reg_13_ ( .D(R9[13]), .RN(n1647), .CK(clk), .Q(R10[13]) );
  DFFTRX1 R11_reg_13_ ( .D(R10[13]), .RN(n1647), .CK(clk), .Q(R11[13]) );
  DFFTRX1 R12_reg_13_ ( .D(R11[13]), .RN(n1648), .CK(clk), .Q(R12[13]) );
  DFFTRX1 R13_reg_13_ ( .D(R12[13]), .RN(n1648), .CK(clk), .Q(R13[13]) );
  DFFTRX1 R2_reg_12_ ( .D(R1[12]), .RN(n1648), .CK(clk), .Q(R2[12]) );
  DFFTRX1 R3_reg_12_ ( .D(R2[12]), .RN(n1648), .CK(clk), .Q(R3[12]) );
  DFFTRX1 R4_reg_12_ ( .D(R3[12]), .RN(n1648), .CK(clk), .Q(R4[12]) );
  DFFTRX1 R5_reg_12_ ( .D(R4[12]), .RN(n1648), .CK(clk), .Q(R5[12]) );
  DFFTRX1 R7_reg_12_ ( .D(R6[12]), .RN(n1648), .CK(clk), .Q(R7[12]) );
  DFFTRX1 R8_reg_12_ ( .D(R7[12]), .RN(n1648), .CK(clk), .Q(R8[12]) );
  DFFTRX1 R9_reg_12_ ( .D(R8[12]), .RN(n1648), .CK(clk), .Q(R9[12]) );
  DFFTRX1 R10_reg_12_ ( .D(R9[12]), .RN(n1648), .CK(clk), .Q(R10[12]) );
  DFFTRX1 R11_reg_12_ ( .D(R10[12]), .RN(n1648), .CK(clk), .Q(R11[12]) );
  DFFTRX1 R12_reg_12_ ( .D(R11[12]), .RN(n1648), .CK(clk), .Q(R12[12]) );
  DFFTRX1 R13_reg_12_ ( .D(R12[12]), .RN(n1649), .CK(clk), .Q(R13[12]) );
  DFFTRX1 R2_reg_11_ ( .D(R1[11]), .RN(n1649), .CK(clk), .Q(R2[11]) );
  DFFTRX1 R3_reg_11_ ( .D(R2[11]), .RN(n1649), .CK(clk), .Q(R3[11]) );
  DFFTRX1 R4_reg_11_ ( .D(R3[11]), .RN(n1649), .CK(clk), .Q(R4[11]) );
  DFFTRX1 R5_reg_11_ ( .D(R4[11]), .RN(n1649), .CK(clk), .Q(R5[11]) );
  DFFTRX1 R7_reg_11_ ( .D(R6[11]), .RN(n1649), .CK(clk), .Q(R7[11]) );
  DFFTRX1 R8_reg_11_ ( .D(R7[11]), .RN(n1649), .CK(clk), .Q(R8[11]) );
  DFFTRX1 R9_reg_11_ ( .D(R8[11]), .RN(n1649), .CK(clk), .Q(R9[11]) );
  DFFTRX1 R10_reg_11_ ( .D(R9[11]), .RN(n1649), .CK(clk), .Q(R10[11]) );
  DFFTRX1 R11_reg_11_ ( .D(R10[11]), .RN(n1649), .CK(clk), .Q(R11[11]) );
  DFFTRX1 R12_reg_11_ ( .D(R11[11]), .RN(n1649), .CK(clk), .Q(R12[11]) );
  DFFTRX1 R13_reg_11_ ( .D(R12[11]), .RN(n1649), .CK(clk), .Q(R13[11]) );
  DFFTRX1 R2_reg_10_ ( .D(R1[10]), .RN(n1650), .CK(clk), .Q(R2[10]) );
  DFFTRX1 R3_reg_10_ ( .D(R2[10]), .RN(n1650), .CK(clk), .Q(R3[10]) );
  DFFTRX1 R4_reg_10_ ( .D(R3[10]), .RN(n1650), .CK(clk), .Q(R4[10]) );
  DFFTRX1 R5_reg_10_ ( .D(R4[10]), .RN(n1650), .CK(clk), .Q(R5[10]) );
  DFFTRX1 R7_reg_10_ ( .D(R6[10]), .RN(n1650), .CK(clk), .Q(R7[10]) );
  DFFTRX1 R8_reg_10_ ( .D(R7[10]), .RN(n1650), .CK(clk), .Q(R8[10]) );
  DFFTRX1 R9_reg_10_ ( .D(R8[10]), .RN(n1650), .CK(clk), .Q(R9[10]) );
  DFFTRX1 R10_reg_10_ ( .D(R9[10]), .RN(n1650), .CK(clk), .Q(R10[10]) );
  DFFTRX1 R11_reg_10_ ( .D(R10[10]), .RN(n1650), .CK(clk), .Q(R11[10]) );
  DFFTRX1 R12_reg_10_ ( .D(R11[10]), .RN(n1650), .CK(clk), .Q(R12[10]) );
  DFFTRX1 R13_reg_10_ ( .D(R12[10]), .RN(n1650), .CK(clk), .Q(R13[10]) );
  DFFTRX1 R2_reg_9_ ( .D(R1[9]), .RN(n1650), .CK(clk), .Q(R2[9]) );
  DFFTRX1 R3_reg_9_ ( .D(R2[9]), .RN(n1651), .CK(clk), .Q(R3[9]) );
  DFFTRX1 R4_reg_9_ ( .D(R3[9]), .RN(n1651), .CK(clk), .Q(R4[9]) );
  DFFTRX1 R5_reg_9_ ( .D(R4[9]), .RN(n1651), .CK(clk), .Q(R5[9]) );
  DFFTRX1 R7_reg_9_ ( .D(R6[9]), .RN(n1651), .CK(clk), .Q(R7[9]) );
  DFFTRX1 R8_reg_9_ ( .D(R7[9]), .RN(n1651), .CK(clk), .Q(R8[9]) );
  DFFTRX1 R9_reg_9_ ( .D(R8[9]), .RN(n1651), .CK(clk), .Q(R9[9]) );
  DFFTRX1 R10_reg_9_ ( .D(R9[9]), .RN(n1651), .CK(clk), .Q(R10[9]) );
  DFFTRX1 R11_reg_9_ ( .D(R10[9]), .RN(n1651), .CK(clk), .Q(R11[9]) );
  DFFTRX1 R12_reg_9_ ( .D(R11[9]), .RN(n1651), .CK(clk), .Q(R12[9]) );
  DFFTRX1 R13_reg_9_ ( .D(R12[9]), .RN(n1651), .CK(clk), .Q(R13[9]) );
  DFFTRX1 R2_reg_8_ ( .D(R1[8]), .RN(n1651), .CK(clk), .Q(R2[8]) );
  DFFTRX1 R3_reg_8_ ( .D(R2[8]), .RN(n1651), .CK(clk), .Q(R3[8]) );
  DFFTRX1 R4_reg_8_ ( .D(R3[8]), .RN(n1652), .CK(clk), .Q(R4[8]) );
  DFFTRX1 R5_reg_8_ ( .D(R4[8]), .RN(n1652), .CK(clk), .Q(R5[8]) );
  DFFTRX1 R7_reg_8_ ( .D(R6[8]), .RN(n1652), .CK(clk), .Q(R7[8]) );
  DFFTRX1 R8_reg_8_ ( .D(R7[8]), .RN(n1652), .CK(clk), .Q(R8[8]) );
  DFFTRX1 R9_reg_8_ ( .D(R8[8]), .RN(n1652), .CK(clk), .Q(R9[8]) );
  DFFTRX1 R10_reg_8_ ( .D(R9[8]), .RN(n1652), .CK(clk), .Q(R10[8]) );
  DFFTRX1 R11_reg_8_ ( .D(R10[8]), .RN(n1652), .CK(clk), .Q(R11[8]) );
  DFFTRX1 R12_reg_8_ ( .D(R11[8]), .RN(n1652), .CK(clk), .Q(R12[8]) );
  DFFTRX1 R2_reg_7_ ( .D(R1[7]), .RN(n1652), .CK(clk), .Q(R2[7]) );
  DFFTRX1 R3_reg_7_ ( .D(R2[7]), .RN(n1652), .CK(clk), .Q(R3[7]) );
  DFFTRX1 R4_reg_7_ ( .D(R3[7]), .RN(n1652), .CK(clk), .Q(R4[7]) );
  DFFTRX1 R5_reg_7_ ( .D(R4[7]), .RN(n1652), .CK(clk), .Q(R5[7]) );
  DFFTRX1 R7_reg_7_ ( .D(R6[7]), .RN(n1653), .CK(clk), .Q(R7[7]) );
  DFFTRX1 R8_reg_7_ ( .D(R7[7]), .RN(n1653), .CK(clk), .Q(R8[7]) );
  DFFTRX1 R9_reg_7_ ( .D(R8[7]), .RN(n1653), .CK(clk), .Q(R9[7]) );
  DFFTRX1 R10_reg_7_ ( .D(R9[7]), .RN(n1653), .CK(clk), .Q(R10[7]) );
  DFFTRX1 R11_reg_7_ ( .D(R10[7]), .RN(n1653), .CK(clk), .Q(R11[7]) );
  DFFTRX1 R12_reg_7_ ( .D(R11[7]), .RN(n1653), .CK(clk), .Q(R12[7]) );
  DFFTRX1 R13_reg_7_ ( .D(R12[7]), .RN(n1653), .CK(clk), .Q(R13[7]) );
  DFFTRX1 R2_reg_6_ ( .D(R1[6]), .RN(n1653), .CK(clk), .Q(R2[6]) );
  DFFTRX1 R3_reg_6_ ( .D(R2[6]), .RN(n1653), .CK(clk), .Q(R3[6]) );
  DFFTRX1 R4_reg_6_ ( .D(R3[6]), .RN(n1653), .CK(clk), .Q(R4[6]) );
  DFFTRX1 R5_reg_6_ ( .D(R4[6]), .RN(n1653), .CK(clk), .Q(R5[6]) );
  DFFTRX1 R7_reg_6_ ( .D(R6[6]), .RN(n1653), .CK(clk), .Q(R7[6]) );
  DFFTRX1 R8_reg_6_ ( .D(R7[6]), .RN(n1654), .CK(clk), .Q(R8[6]) );
  DFFTRX1 R9_reg_6_ ( .D(R8[6]), .RN(n1654), .CK(clk), .Q(R9[6]) );
  DFFTRX1 R10_reg_6_ ( .D(R9[6]), .RN(n1654), .CK(clk), .Q(R10[6]) );
  DFFTRX1 R11_reg_6_ ( .D(R10[6]), .RN(n1654), .CK(clk), .Q(R11[6]) );
  DFFTRX1 R12_reg_6_ ( .D(R11[6]), .RN(n1654), .CK(clk), .Q(R12[6]) );
  DFFTRX1 R13_reg_6_ ( .D(R12[6]), .RN(n1654), .CK(clk), .Q(R13[6]) );
  DFFTRX1 R2_reg_5_ ( .D(R1[5]), .RN(n1654), .CK(clk), .Q(R2[5]) );
  DFFTRX1 R3_reg_5_ ( .D(R2[5]), .RN(n1654), .CK(clk), .Q(R3[5]) );
  DFFTRX1 R4_reg_5_ ( .D(R3[5]), .RN(n1654), .CK(clk), .Q(R4[5]) );
  DFFTRX1 R5_reg_5_ ( .D(R4[5]), .RN(n1654), .CK(clk), .Q(R5[5]) );
  DFFTRX1 R7_reg_5_ ( .D(R6[5]), .RN(n1654), .CK(clk), .Q(R7[5]) );
  DFFTRX1 R8_reg_5_ ( .D(R7[5]), .RN(n1654), .CK(clk), .Q(R8[5]) );
  DFFTRX1 R9_reg_5_ ( .D(R8[5]), .RN(n1655), .CK(clk), .Q(R9[5]) );
  DFFTRX1 R10_reg_5_ ( .D(R9[5]), .RN(n1655), .CK(clk), .Q(R10[5]) );
  DFFTRX1 R11_reg_5_ ( .D(R10[5]), .RN(n1655), .CK(clk), .Q(R11[5]) );
  DFFTRX1 R12_reg_5_ ( .D(R11[5]), .RN(n1655), .CK(clk), .Q(R12[5]) );
  DFFTRX1 R13_reg_5_ ( .D(R12[5]), .RN(n1655), .CK(clk), .Q(R13[5]) );
  DFFTRX1 R2_reg_4_ ( .D(R1[4]), .RN(n1655), .CK(clk), .Q(R2[4]) );
  DFFTRX1 R3_reg_4_ ( .D(R2[4]), .RN(n1655), .CK(clk), .Q(R3[4]) );
  DFFTRX1 R4_reg_4_ ( .D(R3[4]), .RN(n1655), .CK(clk), .Q(R4[4]) );
  DFFTRX1 R5_reg_4_ ( .D(R4[4]), .RN(n1655), .CK(clk), .Q(R5[4]) );
  DFFTRX1 R7_reg_4_ ( .D(R6[4]), .RN(n1655), .CK(clk), .Q(R7[4]) );
  DFFTRX1 R8_reg_4_ ( .D(R7[4]), .RN(n1655), .CK(clk), .Q(R8[4]) );
  DFFTRX1 R9_reg_4_ ( .D(R8[4]), .RN(n1655), .CK(clk), .Q(R9[4]) );
  DFFTRX1 R15_reg_4_ ( .D(R14[4]), .RN(n1661), .CK(clk), .Q(R15[4]) );
  DFFTRX4 R14_reg_9_ ( .D(R13[9]), .RN(n1661), .CK(clk), .Q(R14[9]) );
  DFFTRX4 R1_reg_10_ ( .D(Wt[10]), .RN(n1661), .CK(clk), .Q(R1[10]), .QN(n390)
         );
  DFFHQX1 Wt_reg_19_ ( .D(n1748), .CK(clk), .Q(Wt[19]) );
  DFFTRX4 R1_reg_11_ ( .D(Wt[11]), .RN(n1661), .CK(clk), .Q(R1[11]), .QN(n391)
         );
  DFFTRX4 R14_reg_24_ ( .D(R13[24]), .RN(n1629), .CK(clk), .Q(R14[24]), .QN(
        n400) );
  DFFTRX4 R14_reg_23_ ( .D(R13[23]), .RN(n1629), .CK(clk), .Q(R14[23]), .QN(
        n36) );
  DFFTRX4 R1_reg_21_ ( .D(Wt[21]), .RN(n1660), .CK(clk), .Q(R1[21]), .QN(n5)
         );
  DFFTRX1 R1_reg_12_ ( .D(Wt[12]), .RN(n1660), .CK(clk), .Q(R1[12]), .QN(n393)
         );
  DFFTRX1 R1_reg_13_ ( .D(Wt[13]), .RN(n1630), .CK(clk), .Q(R1[13]), .QN(n394)
         );
  DFFTRX4 R14_reg_8_ ( .D(R13[8]), .RN(n1660), .CK(clk), .Q(R14[8]), .QN(n16)
         );
  DFFTRX4 R6_reg_0_ ( .D(R5[0]), .RN(n1661), .CK(clk), .Q(R6[0]) );
  DFFTRXL counter_reg_5_ ( .D(N627), .RN(n1728), .CK(clk), .Q(counter[5]), 
        .QN(n491) );
  DFFTRXL counter_reg_4_ ( .D(N626), .RN(n1728), .CK(clk), .Q(counter[4]), 
        .QN(n489) );
  DFFTRXL counter_reg_3_ ( .D(N625), .RN(n1728), .CK(clk), .Q(counter[3]), 
        .QN(n490) );
  DFFTRXL counter_reg_2_ ( .D(N624), .RN(n1728), .CK(clk), .Q(counter[2]), 
        .QN(n488) );
  DFFTRXL counter_reg_1_ ( .D(N623), .RN(n1728), .CK(clk), .Q(counter[1]), 
        .QN(n492) );
  DFFTRXL counter_reg_0_ ( .D(N622), .RN(n1728), .CK(clk), .Q(counter[0]), 
        .QN(n493) );
  DFFTRXL R14_reg_30_ ( .D(R13[30]), .RN(n1728), .CK(clk), .Q(R14[30]), .QN(
        n428) );
  DFFTRXL R14_reg_29_ ( .D(R13[29]), .RN(n1728), .CK(clk), .Q(R14[29]), .QN(
        n426) );
  DFFTRXL R14_reg_28_ ( .D(R13[28]), .RN(n1728), .CK(clk), .Q(R14[28]), .QN(
        n424) );
  DFFTRXL R14_reg_27_ ( .D(R13[27]), .RN(n1728), .CK(clk), .Q(R14[27]), .QN(
        n423) );
  DFFTRXL R14_reg_17_ ( .D(R13[17]), .RN(n1728), .CK(clk), .Q(R14[17]), .QN(
        n422) );
  DFFTRXL R1_reg_31_ ( .D(Wt[31]), .RN(n1728), .CK(clk), .Q(R1[31]), .QN(n430)
         );
  DFFTRXL R1_reg_30_ ( .D(Wt[30]), .RN(n1728), .CK(clk), .Q(R1[30]), .QN(n429)
         );
  DFFTRXL R1_reg_29_ ( .D(Wt[29]), .RN(n1728), .CK(clk), .Q(R1[29]), .QN(n427)
         );
  DFFTRXL R1_reg_9_ ( .D(Wt[9]), .RN(n1728), .CK(clk), .Q(R1[9]), .QN(n470) );
  DFFTRXL R1_reg_8_ ( .D(Wt[8]), .RN(n1728), .CK(clk), .Q(R1[8]), .QN(n460) );
  DFFTRXL R1_reg_7_ ( .D(Wt[7]), .RN(n1728), .CK(clk), .Q(R1[7]), .QN(n459) );
  DFFTRXL R1_reg_6_ ( .D(Wt[6]), .RN(n1728), .CK(clk), .Q(R1[6]), .QN(n458) );
  DFFTRXL R1_reg_5_ ( .D(Wt[5]), .RN(n1728), .CK(clk), .Q(R1[5]), .QN(n457) );
  DFFTRXL R14_reg_31_ ( .D(R13[31]), .RN(n1728), .CK(clk), .Q(R14[31]), .QN(
        n440) );
  DFFTRXL R14_reg_2_ ( .D(R13[2]), .RN(n1728), .CK(clk), .Q(R14[2]), .QN(n442)
         );
  DFFTRXL R14_reg_1_ ( .D(R13[1]), .RN(n1728), .CK(clk), .Q(R14[1]), .QN(n441)
         );
  DFFTRXL R14_reg_0_ ( .D(R13[0]), .RN(n1728), .CK(clk), .Q(R14[0]), .QN(n445)
         );
  DFFTRXL R1_reg_2_ ( .D(Wt[2]), .RN(n1728), .CK(clk), .Q(R1[2]), .QN(n439) );
  DFFTRXL R14_reg_16_ ( .D(R13[16]), .RN(n1728), .CK(clk), .Q(R14[16]), .QN(
        n24) );
  DFFTRXL R1_reg_28_ ( .D(Wt[28]), .RN(n1728), .CK(clk), .Q(R1[28]), .QN(n425)
         );
  DFFHQXL Wt_reg_16_ ( .D(n1745), .CK(clk), .Q(Wt[16]) );
  DFFHQXL Wt_reg_21_ ( .D(n1750), .CK(clk), .Q(Wt[21]) );
  DFFHQXL Wt_reg_20_ ( .D(n1749), .CK(clk), .Q(Wt[20]) );
  DFFHQXL Wt_reg_22_ ( .D(n1751), .CK(clk), .Q(Wt[22]) );
  DFFXL Wt_reg_24_ ( .D(n1753), .CK(clk), .Q(Wt[24]) );
  DFFXL Wt_reg_23_ ( .D(n1752), .CK(clk), .Q(Wt[23]) );
  DFFTRXL R1_reg_16_ ( .D(Wt[16]), .RN(n1628), .CK(clk), .Q(R1[16]), .QN(n407)
         );
  DFFTRXL R1_reg_15_ ( .D(Wt[15]), .RN(n1728), .CK(clk), .Q(R1[15]), .QN(n406)
         );
  DFFTRXL R1_reg_14_ ( .D(Wt[14]), .RN(n1728), .CK(clk), .Q(R1[14]), .QN(n405)
         );
  DFFTRXL R1_reg_23_ ( .D(Wt[23]), .RN(n1728), .CK(clk), .Q(R1[23]), .QN(n392)
         );
  DFFTRXL R14_reg_6_ ( .D(R13[6]), .RN(n1728), .CK(clk), .Q(R14[6]), .QN(n398)
         );
  DFFXL Wt_reg_25_ ( .D(n1754), .CK(clk), .Q(Wt[25]) );
  DFFTRXL R6_reg_2_ ( .D(R5[2]), .RN(n1628), .CK(clk), .Q(R6[2]) );
  DFFTRXL R1_reg_26_ ( .D(Wt[26]), .RN(n1728), .CK(clk), .Q(R1[26]), .QN(n403)
         );
  DFFTRXL R1_reg_25_ ( .D(Wt[25]), .RN(n1728), .CK(clk), .Q(R1[25]) );
  DFFTRXL R1_reg_24_ ( .D(Wt[24]), .RN(n1728), .CK(clk), .Q(R1[24]), .QN(n401)
         );
  DFFTRXL R14_reg_10_ ( .D(R13[10]), .RN(n1728), .CK(clk), .Q(R14[10]), .QN(
        n26) );
  DFFTRXL R15_reg_6_ ( .D(R14[6]), .RN(n1661), .CK(clk), .Q(R15[6]) );
  DFFTRXL R1_reg_22_ ( .D(Wt[22]), .RN(n1629), .CK(clk), .Q(R1[22]), .QN(n397)
         );
  AND2X1 R15_reg_0__U2 ( .A(R14[0]), .B(n1660), .Y(n1188) );
  DFFHQX4 R15_reg_0_ ( .D(n1188), .CK(clk), .Q(R15[0]) );
  DFFTRX4 R1_reg_20_ ( .D(Wt[20]), .RN(n1660), .CK(clk), .Q(R1[20]), .QN(n13)
         );
  DFFTRX2 R1_reg_3_ ( .D(Wt[3]), .RN(n1728), .CK(clk), .Q(R1[3]) );
  DFFTRX4 R14_reg_21_ ( .D(R13[21]), .RN(n1728), .CK(clk), .Q(R14[21]), .QN(
        n396) );
  DFFTRX2 R1_reg_0_ ( .D(Wt[0]), .RN(n1627), .CK(clk), .Q(R1[0]), .QN(n446) );
  DFFTRX1 R1_reg_1_ ( .D(Wt[1]), .RN(n1626), .CK(clk), .Q(R1[1]), .QN(n447) );
  BUFX16 U3 ( .A(n1762), .Y(Wt[0]) );
  CLKINVX3 U4 ( .A(n676), .Y(n1728) );
  NAND3BX4 U5 ( .AN(reset), .B(inner_busy), .C(n677), .Y(n676) );
  XOR3X4 U6 ( .A(R1[11]), .B(n15), .C(n13), .Y(sigma1[1]) );
  OAI21X4 U7 ( .A0(n1195), .A1(n1196), .B0(n1727), .Y(n1760) );
  CLKINVX8 U8 ( .A(logic_result[31]), .Y(n1195) );
  INVXL U9 ( .A(n1553), .Y(n1196) );
  XOR3X4 U10 ( .A(n390), .B(n14), .C(R1[19]), .Y(sigma1[0]) );
  XOR3X4 U11 ( .A(n8), .B(n20), .C(R14[7]), .Y(sigma0[0]) );
  BUFX20 U12 ( .A(n1761), .Y(Wt[1]) );
  CLKINVX8 U13 ( .A(n16), .Y(n1675) );
  XOR3X4 U14 ( .A(R14[8]), .B(R14[4]), .C(R14[19]), .Y(sigma0[1]) );
  NAND2XL U15 ( .A(data[31]), .B(n1616), .Y(n1727) );
  XOR3X2 U16 ( .A(n445), .B(R14[17]), .C(n396), .Y(sigma0[14]) );
  XOR3X2 U17 ( .A(R14[18]), .B(n426), .C(n404), .Y(sigma0[11]) );
  XOR2XL U18 ( .A(n460), .B(n390), .Y(sigma1[23]) );
  NAND2XL U19 ( .A(data[29]), .B(n1616), .Y(n1686) );
  XOR3X2 U20 ( .A(n446), .B(R1[30]), .C(n392), .Y(sigma1[13]) );
  XNOR3X2 U21 ( .A(n458), .B(n460), .C(n430), .Y(sigma1[21]) );
  XOR2XL U22 ( .A(n391), .B(n394), .Y(sigma1[26]) );
  XOR2XL U23 ( .A(n406), .B(n14), .Y(sigma1[30]) );
  NAND2XL U24 ( .A(data[27]), .B(n1616), .Y(n1684) );
  XOR2X1 U25 ( .A(n394), .B(n406), .Y(sigma1[28]) );
  NAND2XL U26 ( .A(data[20]), .B(n1616), .Y(n1723) );
  NAND2XL U27 ( .A(data[19]), .B(n1616), .Y(n1721) );
  XOR3X2 U28 ( .A(R1[2]), .B(R1[4]), .C(R1[27]), .Y(sigma1[17]) );
  NAND2X1 U29 ( .A(write_enable), .B(n1676), .Y(n1199) );
  INVX1 U30 ( .A(n1665), .Y(n1655) );
  INVX1 U31 ( .A(n1665), .Y(n1654) );
  INVX1 U32 ( .A(n1666), .Y(n1653) );
  INVX1 U33 ( .A(n1666), .Y(n1652) );
  INVX1 U34 ( .A(n1667), .Y(n1651) );
  INVX1 U35 ( .A(n1667), .Y(n1650) );
  INVX1 U36 ( .A(n1668), .Y(n1649) );
  INVX1 U37 ( .A(n1668), .Y(n1648) );
  INVX1 U38 ( .A(n1668), .Y(n1647) );
  INVX1 U39 ( .A(n1668), .Y(n1646) );
  INVX1 U40 ( .A(n1621), .Y(n1645) );
  INVX1 U41 ( .A(n1621), .Y(n1644) );
  INVX1 U42 ( .A(n1669), .Y(n1643) );
  INVX1 U43 ( .A(n1669), .Y(n1642) );
  INVX1 U44 ( .A(n1670), .Y(n1641) );
  INVX1 U45 ( .A(n1670), .Y(n1640) );
  INVX1 U46 ( .A(n1671), .Y(n1639) );
  INVX1 U47 ( .A(n1671), .Y(n1638) );
  INVX1 U48 ( .A(n1672), .Y(n1637) );
  INVX1 U49 ( .A(n1672), .Y(n1636) );
  INVX1 U50 ( .A(n1672), .Y(n1635) );
  INVX1 U51 ( .A(n1672), .Y(n1634) );
  INVX1 U52 ( .A(n1621), .Y(n1633) );
  INVX1 U53 ( .A(n1621), .Y(n1632) );
  INVX1 U54 ( .A(n1673), .Y(n1631) );
  INVX1 U55 ( .A(n1673), .Y(n1630) );
  INVX1 U56 ( .A(n1673), .Y(n1629) );
  INVX1 U57 ( .A(n1621), .Y(n1628) );
  INVX1 U58 ( .A(n1664), .Y(n1626) );
  INVX1 U59 ( .A(n1621), .Y(n1625) );
  INVX1 U60 ( .A(n1621), .Y(n1624) );
  INVX1 U61 ( .A(n1663), .Y(n1627) );
  INVX1 U62 ( .A(n1662), .Y(n1660) );
  INVX1 U63 ( .A(n1663), .Y(n1659) );
  INVX1 U64 ( .A(n1663), .Y(n1658) );
  INVX1 U65 ( .A(n1664), .Y(n1657) );
  INVX1 U66 ( .A(n1664), .Y(n1656) );
  INVX1 U67 ( .A(n1662), .Y(n1661) );
  INVX1 U68 ( .A(n1618), .Y(n1665) );
  INVX1 U69 ( .A(n1618), .Y(n1666) );
  INVX1 U70 ( .A(n1618), .Y(n1667) );
  INVX1 U71 ( .A(n1619), .Y(n1668) );
  INVX1 U72 ( .A(n1620), .Y(n1669) );
  INVX1 U73 ( .A(n1620), .Y(n1670) );
  INVX1 U74 ( .A(n1620), .Y(n1671) );
  INVX1 U75 ( .A(n1620), .Y(n1672) );
  INVX1 U76 ( .A(n1620), .Y(n1673) );
  INVX1 U77 ( .A(n1623), .Y(n1618) );
  INVX1 U78 ( .A(n1623), .Y(n1619) );
  INVX1 U79 ( .A(n1622), .Y(n1620) );
  INVX1 U80 ( .A(n1617), .Y(n1663) );
  INVX1 U81 ( .A(n1617), .Y(n1664) );
  INVX1 U82 ( .A(n1617), .Y(n1662) );
  INVX1 U83 ( .A(n1623), .Y(n1617) );
  INVX1 U84 ( .A(n1728), .Y(n1623) );
  INVX1 U85 ( .A(n1728), .Y(n1622) );
  INVX1 U86 ( .A(n1728), .Y(n1621) );
  INVX1 U87 ( .A(n676), .Y(n1676) );
  BUFX3 U88 ( .A(n1726), .Y(n1616) );
  INVXL U89 ( .A(n1199), .Y(n1726) );
  BUFX3 U90 ( .A(n1553), .Y(n1615) );
  XOR3X2 U91 ( .A(n426), .B(n441), .C(R14[12]), .Y(sigma0[26]) );
  XOR3X2 U92 ( .A(R14[14]), .B(n440), .C(n20), .Y(sigma0[28]) );
  XOR3X2 U93 ( .A(n36), .B(n412), .C(n1675), .Y(sigma0[5]) );
  XOR3X2 U94 ( .A(n401), .B(n406), .C(R1[22]), .Y(sigma1[5]) );
  XOR3X2 U95 ( .A(n400), .B(n32), .C(R14[9]), .Y(sigma0[6]) );
  XOR3X2 U96 ( .A(n392), .B(n407), .C(R1[25]), .Y(sigma1[6]) );
  XOR2X1 U97 ( .A(n11), .B(n24), .Y(sigma0[30]) );
  XOR2X1 U98 ( .A(n470), .B(n391), .Y(sigma1[24]) );
  XOR3X2 U99 ( .A(n423), .B(n440), .C(R14[10]), .Y(sigma0[24]) );
  XOR2X1 U100 ( .A(n398), .B(n422), .Y(sigma0[31]) );
  XOR2X1 U101 ( .A(n407), .B(n15), .Y(sigma1[31]) );
  XOR3X2 U102 ( .A(n36), .B(n442), .C(R14[19]), .Y(sigma0[16]) );
  XOR3X2 U103 ( .A(n403), .B(n447), .C(R1[3]), .Y(sigma1[16]) );
  XOR3X2 U104 ( .A(n8), .B(n441), .C(R14[22]), .Y(sigma0[15]) );
  XOR3X2 U105 ( .A(n446), .B(n439), .C(R1[25]), .Y(sigma1[15]) );
  XOR3X2 U106 ( .A(n410), .B(n428), .C(R14[9]), .Y(sigma0[23]) );
  XOR3X2 U107 ( .A(n400), .B(n424), .C(R14[7]), .Y(sigma0[21]) );
  XOR3X2 U108 ( .A(n408), .B(n28), .C(R14[7]), .Y(sigma0[4]) );
  XOR3X2 U109 ( .A(n392), .B(n405), .C(R1[21]), .Y(sigma1[4]) );
  XOR2X1 U110 ( .A(n459), .B(n470), .Y(sigma1[22]) );
  XOR3X2 U111 ( .A(n409), .B(n426), .C(n1675), .Y(sigma0[22]) );
  XOR3X2 U112 ( .A(n36), .B(n423), .C(R14[6]), .Y(sigma0[20]) );
  XOR3X2 U113 ( .A(n457), .B(n459), .C(R1[30]), .Y(sigma1[20]) );
  XOR3X2 U114 ( .A(n428), .B(n30), .C(R14[19]), .Y(sigma0[12]) );
  XOR3X2 U115 ( .A(n427), .B(n430), .C(R1[22]), .Y(sigma1[12]) );
  XOR3X2 U116 ( .A(n440), .B(n24), .C(R14[20]), .Y(sigma0[13]) );
  XOR3X2 U117 ( .A(n447), .B(n430), .C(R1[24]), .Y(sigma1[14]) );
  XOR3X2 U118 ( .A(n425), .B(n429), .C(R1[21]), .Y(sigma1[11]) );
  XOR2X1 U119 ( .A(n9), .B(n30), .Y(sigma0[29]) );
  XOR2X1 U120 ( .A(n405), .B(n407), .Y(sigma1[29]) );
  XOR3X2 U121 ( .A(n395), .B(n11), .C(R14[9]), .Y(sigma0[2]) );
  XOR3X2 U122 ( .A(n12), .B(n5), .C(R1[12]), .Y(sigma1[2]) );
  XOR3X2 U123 ( .A(n396), .B(n26), .C(R14[6]), .Y(sigma0[3]) );
  XOR3X2 U124 ( .A(n397), .B(n394), .C(R1[20]), .Y(sigma1[3]) );
  XOR3X2 U125 ( .A(n409), .B(n404), .C(R14[10]), .Y(sigma0[7]) );
  XOR3X2 U126 ( .A(n403), .B(n14), .C(R1[24]), .Y(sigma1[7]) );
  XOR3X2 U127 ( .A(n410), .B(n30), .C(R14[11]), .Y(sigma0[8]) );
  XOR3X2 U128 ( .A(n411), .B(n15), .C(R1[25]), .Y(sigma1[8]) );
  XOR3X2 U129 ( .A(n423), .B(n24), .C(R14[12]), .Y(sigma0[9]) );
  XOR3X2 U130 ( .A(n403), .B(n425), .C(R1[19]), .Y(sigma1[9]) );
  XOR3X2 U131 ( .A(n424), .B(n422), .C(R14[13]), .Y(sigma0[10]) );
  XOR3X2 U132 ( .A(n411), .B(n427), .C(R1[20]), .Y(sigma1[10]) );
  XOR2X1 U133 ( .A(n393), .B(n405), .Y(sigma1[27]) );
  XOR3X2 U134 ( .A(n428), .B(n442), .C(R14[13]), .Y(sigma0[27]) );
  XOR3X2 U135 ( .A(n396), .B(n409), .C(n1674), .Y(sigma0[18]) );
  XOR3X2 U136 ( .A(n425), .B(n457), .C(R1[3]), .Y(sigma1[18]) );
  OAI2BB1X1 U137 ( .A0N(logic_result[30]), .A1N(n1615), .B0(n1687), .Y(n1759)
         );
  NAND2X1 U138 ( .A(data[30]), .B(n1616), .Y(n1687) );
  OAI2BB1X1 U139 ( .A0N(logic_result[29]), .A1N(n1615), .B0(n1686), .Y(n1758)
         );
  OAI2BB1X1 U140 ( .A0N(logic_result[28]), .A1N(n1615), .B0(n1682), .Y(n1757)
         );
  NAND2X1 U141 ( .A(data[28]), .B(n1616), .Y(n1682) );
  OAI2BB1X1 U142 ( .A0N(logic_result[27]), .A1N(n1615), .B0(n1684), .Y(n1756)
         );
  OAI2BB1X1 U143 ( .A0N(logic_result[25]), .A1N(n1615), .B0(n1685), .Y(n1754)
         );
  NAND2X1 U144 ( .A(data[25]), .B(n1616), .Y(n1685) );
  OAI2BB1X1 U145 ( .A0N(logic_result[26]), .A1N(n1615), .B0(n1683), .Y(n1755)
         );
  NAND2X1 U146 ( .A(data[26]), .B(n1616), .Y(n1683) );
  OAI2BB1X1 U147 ( .A0N(logic_result[24]), .A1N(n1615), .B0(n1681), .Y(n1753)
         );
  NAND2X1 U148 ( .A(data[24]), .B(n1616), .Y(n1681) );
  OAI2BB1X1 U149 ( .A0N(logic_result[23]), .A1N(n1615), .B0(n1725), .Y(n1752)
         );
  NAND2X1 U150 ( .A(data[23]), .B(n1616), .Y(n1725) );
  OAI2BB1X1 U151 ( .A0N(logic_result[19]), .A1N(n1615), .B0(n1721), .Y(n1748)
         );
  OAI2BB1X1 U152 ( .A0N(logic_result[22]), .A1N(n1615), .B0(n1722), .Y(n1751)
         );
  NAND2X1 U153 ( .A(data[22]), .B(n1616), .Y(n1722) );
  OAI2BB1X1 U154 ( .A0N(logic_result[20]), .A1N(n1615), .B0(n1723), .Y(n1749)
         );
  OAI2BB1X1 U155 ( .A0N(logic_result[21]), .A1N(n1615), .B0(n1724), .Y(n1750)
         );
  NAND2X1 U156 ( .A(data[21]), .B(n1616), .Y(n1724) );
  NAND4BXL U157 ( .AN(n678), .B(n491), .C(n493), .D(n492), .Y(n677) );
  NAND4X1 U158 ( .A(n490), .B(n489), .C(n488), .D(counter[6]), .Y(n678) );
  OAI22XL U159 ( .A0(n1199), .A1(n1678), .B0(n1717), .B1(n1677), .Y(n1730) );
  INVX1 U160 ( .A(logic_result[1]), .Y(n1677) );
  INVX1 U161 ( .A(data[1]), .Y(n1678) );
  OAI22XL U162 ( .A0(n1199), .A1(n1680), .B0(n1717), .B1(n1679), .Y(n1732) );
  INVX1 U163 ( .A(logic_result[3]), .Y(n1679) );
  INVX1 U164 ( .A(data[3]), .Y(n1680) );
  OAI22XL U165 ( .A0(n1199), .A1(n1689), .B0(n1717), .B1(n1688), .Y(n1733) );
  INVX1 U166 ( .A(logic_result[4]), .Y(n1688) );
  INVX1 U167 ( .A(data[4]), .Y(n1689) );
  OAI22XL U168 ( .A0(n1199), .A1(n1691), .B0(n1717), .B1(n1690), .Y(n1734) );
  INVX1 U169 ( .A(logic_result[5]), .Y(n1690) );
  INVX1 U170 ( .A(data[5]), .Y(n1691) );
  OAI22XL U171 ( .A0(n1199), .A1(n1693), .B0(n1717), .B1(n1692), .Y(n1735) );
  INVX1 U172 ( .A(logic_result[6]), .Y(n1692) );
  INVX1 U173 ( .A(data[6]), .Y(n1693) );
  OAI22XL U174 ( .A0(n1199), .A1(n1695), .B0(n1717), .B1(n1694), .Y(n1736) );
  INVX1 U175 ( .A(logic_result[7]), .Y(n1694) );
  INVX1 U176 ( .A(data[7]), .Y(n1695) );
  OAI22XL U177 ( .A0(n1199), .A1(n1697), .B0(n1717), .B1(n1696), .Y(n1738) );
  INVX1 U178 ( .A(logic_result[9]), .Y(n1696) );
  INVX1 U179 ( .A(data[9]), .Y(n1697) );
  OAI22XL U180 ( .A0(n1199), .A1(n1699), .B0(n1717), .B1(n1698), .Y(n1737) );
  INVX1 U181 ( .A(logic_result[8]), .Y(n1698) );
  INVX1 U182 ( .A(data[8]), .Y(n1699) );
  OAI22XL U183 ( .A0(n1199), .A1(n1701), .B0(n1717), .B1(n1700), .Y(n1731) );
  INVX1 U184 ( .A(logic_result[2]), .Y(n1700) );
  INVX1 U185 ( .A(data[2]), .Y(n1701) );
  OAI22XL U186 ( .A0(n1199), .A1(n1703), .B0(n1717), .B1(n1702), .Y(n1729) );
  INVX1 U187 ( .A(logic_result[0]), .Y(n1702) );
  INVX1 U188 ( .A(data[0]), .Y(n1703) );
  OAI22XL U189 ( .A0(n1199), .A1(n1705), .B0(n1717), .B1(n1704), .Y(n1739) );
  INVX1 U190 ( .A(logic_result[10]), .Y(n1704) );
  INVX1 U191 ( .A(data[10]), .Y(n1705) );
  OAI22XL U192 ( .A0(n1199), .A1(n1707), .B0(n1717), .B1(n1706), .Y(n1740) );
  INVX1 U193 ( .A(logic_result[11]), .Y(n1706) );
  INVX1 U194 ( .A(data[11]), .Y(n1707) );
  OAI22XL U195 ( .A0(n1199), .A1(n1709), .B0(n1717), .B1(n1708), .Y(n1741) );
  INVX1 U196 ( .A(logic_result[12]), .Y(n1708) );
  INVX1 U197 ( .A(data[12]), .Y(n1709) );
  OAI22XL U198 ( .A0(n1199), .A1(n1711), .B0(n1717), .B1(n1710), .Y(n1742) );
  INVX1 U199 ( .A(logic_result[13]), .Y(n1710) );
  INVX1 U200 ( .A(data[13]), .Y(n1711) );
  OAI22XL U201 ( .A0(n1199), .A1(n1713), .B0(n1717), .B1(n1712), .Y(n1743) );
  INVX1 U202 ( .A(logic_result[14]), .Y(n1712) );
  INVX1 U203 ( .A(data[14]), .Y(n1713) );
  OAI22XL U204 ( .A0(n1199), .A1(n1715), .B0(n1717), .B1(n1714), .Y(n1744) );
  INVX1 U205 ( .A(logic_result[15]), .Y(n1714) );
  INVX1 U206 ( .A(data[15]), .Y(n1715) );
  OAI22XL U207 ( .A0(n1199), .A1(n1718), .B0(n1717), .B1(n1716), .Y(n1745) );
  INVX1 U208 ( .A(data[16]), .Y(n1718) );
  INVX1 U209 ( .A(logic_result[16]), .Y(n1716) );
  XOR3X2 U210 ( .A(n400), .B(n20), .C(R14[20]), .Y(sigma0[17]) );
  NOR2BX1 U211 ( .AN(n1676), .B(write_enable), .Y(n1553) );
  INVX1 U212 ( .A(n1553), .Y(n1717) );
  OAI2BB2X1 U213 ( .B0(n1199), .B1(n1719), .A0N(logic_result[17]), .A1N(n1615), 
        .Y(n1746) );
  INVX1 U214 ( .A(data[17]), .Y(n1719) );
  OAI2BB1X1 U215 ( .A0N(logic_result[18]), .A1N(n1615), .B0(n1720), .Y(n1747)
         );
  NAND2X1 U216 ( .A(data[18]), .B(n1616), .Y(n1720) );
  XOR3X2 U217 ( .A(n410), .B(n11), .C(R14[22]), .Y(sigma0[19]) );
  XOR3X2 U218 ( .A(R1[4]), .B(n458), .C(n427), .Y(sigma1[19]) );
  INVXL U219 ( .A(n9), .Y(n1674) );
  XOR3X2 U220 ( .A(n424), .B(n445), .C(R14[11]), .Y(sigma0[25]) );
  XOR2X1 U221 ( .A(n390), .B(n393), .Y(sigma1[25]) );
endmodule


module hash_core_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n34, n37, n38, n39, n24, n33,
         n35, n36, n40, n41, n42, n43, n44, n45;
  wire   [31:2] carry;

  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX4 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX4 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_4 ( .A(A[4]), .B(B[4]), .CI(n45), .CO(carry[5]), .S(SUM[4]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  NAND2X1 U1 ( .A(n36), .B(n40), .Y(n41) );
  INVX4 U2 ( .A(n25), .Y(n45) );
  OAI2BB2X4 U3 ( .B0(n24), .B1(n33), .A0N(n35), .A1N(carry[21]), .Y(carry[22])
         );
  INVX1 U4 ( .A(A[21]), .Y(n24) );
  INVX1 U5 ( .A(B[21]), .Y(n33) );
  AOI22X4 U6 ( .A0(B[3]), .A1(A[3]), .B0(n26), .B1(carry[3]), .Y(n25) );
  OAI211X4 U7 ( .A0(A[1]), .A1(B[1]), .B0(A[0]), .C0(B[0]), .Y(n27) );
  OAI2BB1X2 U8 ( .A0N(A[1]), .A1N(B[1]), .B0(n27), .Y(carry[2]) );
  OR2X2 U9 ( .A(A[21]), .B(B[21]), .Y(n35) );
  NAND2X4 U10 ( .A(n41), .B(carry[11]), .Y(n29) );
  INVXL U11 ( .A(A[11]), .Y(n36) );
  INVX1 U12 ( .A(B[11]), .Y(n40) );
  OAI2BB1X4 U13 ( .A0N(A[11]), .A1N(B[11]), .B0(n29), .Y(carry[12]) );
  OR2X2 U14 ( .A(A[23]), .B(B[23]), .Y(n42) );
  NAND2X4 U15 ( .A(n42), .B(carry[23]), .Y(n28) );
  OAI2BB1X4 U16 ( .A0N(A[23]), .A1N(B[23]), .B0(n28), .Y(carry[24]) );
  XOR2XL U17 ( .A(B[1]), .B(A[1]), .Y(n43) );
  XNOR2X1 U18 ( .A(n44), .B(n43), .Y(SUM[1]) );
  XOR2X1 U19 ( .A(A[3]), .B(B[3]), .Y(n26) );
  AOI22XL U20 ( .A0(B[22]), .A1(n32), .B0(A[22]), .B1(carry[22]), .Y(n31) );
  OR2XL U21 ( .A(carry[22]), .B(A[22]), .Y(n32) );
  XOR2X1 U22 ( .A(n37), .B(n38), .Y(SUM[11]) );
  XOR2X1 U23 ( .A(A[21]), .B(n34), .Y(SUM[21]) );
  XOR2X1 U24 ( .A(n30), .B(n31), .Y(SUM[23]) );
  XOR2X1 U25 ( .A(carry[3]), .B(n26), .Y(SUM[3]) );
  XOR2X1 U26 ( .A(carry[21]), .B(B[21]), .Y(n34) );
  OAI2BB1X1 U27 ( .A0N(A[10]), .A1N(B[10]), .B0(n39), .Y(n37) );
  OAI21XL U28 ( .A0(A[10]), .A1(B[10]), .B0(carry[10]), .Y(n39) );
  XOR2XL U29 ( .A(B[11]), .B(A[11]), .Y(n38) );
  NAND2XL U30 ( .A(A[0]), .B(B[0]), .Y(n44) );
  XNOR2X1 U31 ( .A(A[23]), .B(B[23]), .Y(n30) );
  XOR2XL U32 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module hash_core_DW01_add_1 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n11, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32;
  wire   [31:2] carry;

  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_13 ( .A(A[13]), .B(B[13]), .CI(n11), .CO(carry[14]), .S(SUM[13])
         );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX4 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX4 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  OAI2BB1X4 U1 ( .A0N(n29), .A1N(n30), .B0(carry[16]), .Y(n19) );
  CLKINVX20 U2 ( .A(A[16]), .Y(n29) );
  CLKINVX20 U3 ( .A(B[16]), .Y(n30) );
  OAI211X1 U4 ( .A0(A[1]), .A1(B[1]), .B0(A[0]), .C0(B[0]), .Y(n18) );
  OAI2BB1X4 U5 ( .A0N(A[12]), .A1N(B[12]), .B0(n17), .Y(n11) );
  XOR2XL U6 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X1 U7 ( .A(A[0]), .B(B[0]), .Y(n20) );
  OAI2BB1X4 U8 ( .A0N(A[16]), .A1N(B[16]), .B0(n19), .Y(carry[17]) );
  OAI21X4 U9 ( .A0(A[12]), .A1(B[12]), .B0(carry[12]), .Y(n17) );
  OR2X2 U10 ( .A(A[14]), .B(B[14]), .Y(n31) );
  NAND2X4 U11 ( .A(n31), .B(carry[14]), .Y(n25) );
  OAI2BB1X4 U12 ( .A0N(A[14]), .A1N(B[14]), .B0(n25), .Y(carry[15]) );
  OAI2BB1X2 U13 ( .A0N(A[1]), .A1N(B[1]), .B0(n18), .Y(carry[2]) );
  OAI2BB1XL U14 ( .A0N(A[14]), .A1N(B[14]), .B0(n25), .Y(n32) );
  AOI22XL U15 ( .A0(B[15]), .A1(n24), .B0(A[15]), .B1(n32), .Y(n23) );
  OR2XL U16 ( .A(n32), .B(A[15]), .Y(n24) );
  XOR2X1 U17 ( .A(n22), .B(n23), .Y(SUM[16]) );
  XNOR2X1 U18 ( .A(A[16]), .B(B[16]), .Y(n22) );
  XOR2X1 U19 ( .A(n26), .B(n27), .Y(SUM[14]) );
  XOR2X1 U20 ( .A(B[14]), .B(A[14]), .Y(n27) );
  OAI2BB1X1 U21 ( .A0N(A[13]), .A1N(B[13]), .B0(n28), .Y(n26) );
  OAI21XL U22 ( .A0(A[13]), .A1(B[13]), .B0(carry[13]), .Y(n28) );
  XOR2X1 U23 ( .A(n20), .B(n21), .Y(SUM[1]) );
  XOR2X1 U24 ( .A(B[1]), .B(A[1]), .Y(n21) );
endmodule


module hash_core_DW01_add_2 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n35, n36, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50,
         n32, n33, n34, n37, n46, n51, n52, n53, n54, n55;
  wire   [31:3] carry;

  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX4 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX4 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(n32), .CO(carry[29]), .S(SUM[28])
         );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(n55), .CO(carry[11]), .S(SUM[10])
         );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(n54), .CO(carry[22]), .S(SUM[21])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX4 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  OAI2BB2X4 U1 ( .B0(n33), .B1(n34), .A0N(n38), .A1N(carry[27]), .Y(n32) );
  CLKINVX20 U2 ( .A(B[27]), .Y(n33) );
  CLKINVX20 U3 ( .A(A[27]), .Y(n34) );
  AOI22X2 U4 ( .A0(B[9]), .A1(A[9]), .B0(n43), .B1(carry[9]), .Y(n42) );
  INVX1 U5 ( .A(n42), .Y(n55) );
  OAI2BB1X1 U6 ( .A0N(A[25]), .A1N(B[25]), .B0(n39), .Y(carry[26]) );
  NAND2X2 U7 ( .A(n37), .B(carry[25]), .Y(n39) );
  AOI22X4 U8 ( .A0(B[20]), .A1(A[20]), .B0(n41), .B1(carry[20]), .Y(n40) );
  OAI2BB1X4 U9 ( .A0N(A[23]), .A1N(B[23]), .B0(n49), .Y(carry[24]) );
  OAI211X2 U10 ( .A0(A[1]), .A1(B[1]), .B0(A[0]), .C0(B[0]), .Y(n45) );
  OAI21X2 U11 ( .A0(A[2]), .A1(n35), .B0(B[2]), .Y(n36) );
  OAI2BB1X1 U12 ( .A0N(n35), .A1N(A[2]), .B0(n36), .Y(carry[3]) );
  OAI21X4 U13 ( .A0(A[23]), .A1(B[23]), .B0(carry[23]), .Y(n49) );
  OR2XL U14 ( .A(A[25]), .B(B[25]), .Y(n37) );
  OAI2BB1X4 U15 ( .A0N(A[1]), .A1N(B[1]), .B0(n45), .Y(n35) );
  OAI2BB1XL U16 ( .A0N(A[23]), .A1N(B[23]), .B0(n49), .Y(n46) );
  XOR2XL U17 ( .A(B[2]), .B(A[2]), .Y(n44) );
  XNOR2X1 U18 ( .A(n51), .B(n47), .Y(SUM[25]) );
  XOR2X1 U19 ( .A(A[25]), .B(B[25]), .Y(n51) );
  AOI22XL U20 ( .A0(B[24]), .A1(n48), .B0(A[24]), .B1(n46), .Y(n47) );
  OR2XL U21 ( .A(n46), .B(A[24]), .Y(n48) );
  XNOR2XL U22 ( .A(B[1]), .B(A[1]), .Y(n53) );
  XOR2X1 U23 ( .A(A[23]), .B(n50), .Y(SUM[23]) );
  XOR2X1 U24 ( .A(carry[9]), .B(n43), .Y(SUM[9]) );
  XOR2X1 U25 ( .A(carry[27]), .B(n38), .Y(SUM[27]) );
  INVX2 U26 ( .A(n40), .Y(n54) );
  XOR2X1 U27 ( .A(A[9]), .B(B[9]), .Y(n43) );
  XOR2X1 U28 ( .A(carry[20]), .B(n41), .Y(SUM[20]) );
  XOR2X1 U29 ( .A(carry[23]), .B(B[23]), .Y(n50) );
  XOR2X1 U30 ( .A(A[20]), .B(B[20]), .Y(n41) );
  XOR2X1 U31 ( .A(A[27]), .B(B[27]), .Y(n38) );
  XOR2X1 U32 ( .A(n52), .B(n53), .Y(SUM[1]) );
  NAND2XL U33 ( .A(A[0]), .B(B[0]), .Y(n52) );
  XOR2X1 U34 ( .A(n35), .B(n44), .Y(SUM[2]) );
  XOR2XL U35 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module hash_core_DW01_add_4 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n5, n32, n33, n34, n36, n37, n38, n40, n42, n43, n44, n45, n27, n28,
         n29, n30, n31, n35, n39, n41, n46, n47, n48, n49;
  wire   [30:2] carry;

  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(n49), .CO(carry[8]), .S(SUM[7]) );
  ADDFHX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(n48), .CO(carry[24]), .S(SUM[23])
         );
  ADDFHX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(n30), .CO(carry[21]), .S(SUM[20])
         );
  ADDFHX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(n27), .CO(carry[17]), .S(SUM[16])
         );
  ADDFHXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX4 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(n39), .Y(SUM[31]) );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n5), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX4 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX4 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX4 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2X2 U1 ( .A(A[0]), .B(B[0]), .Y(n5) );
  INVX1 U2 ( .A(B[30]), .Y(n41) );
  ADDFHX2 U3 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(n47) );
  INVX1 U4 ( .A(A[30]), .Y(n46) );
  OAI2BB2X4 U5 ( .B0(n28), .B1(n29), .A0N(n42), .A1N(n47), .Y(n27) );
  CLKINVX20 U6 ( .A(B[15]), .Y(n28) );
  CLKINVX20 U7 ( .A(A[15]), .Y(n29) );
  OAI2BB2X4 U8 ( .B0(n31), .B1(n35), .A0N(n40), .A1N(carry[19]), .Y(n30) );
  CLKINVX20 U9 ( .A(B[19]), .Y(n31) );
  CLKINVX20 U10 ( .A(A[19]), .Y(n35) );
  OAI2BB2X4 U11 ( .B0(n41), .B1(n46), .A0N(n36), .A1N(carry[30]), .Y(n39) );
  OAI2BB1X4 U12 ( .A0N(A[4]), .A1N(B[4]), .B0(n34), .Y(carry[5]) );
  AOI22X4 U13 ( .A0(B[6]), .A1(A[6]), .B0(n33), .B1(carry[6]), .Y(n32) );
  AOI22X4 U14 ( .A0(B[22]), .A1(A[22]), .B0(n38), .B1(carry[22]), .Y(n37) );
  OAI21X4 U15 ( .A0(A[4]), .A1(B[4]), .B0(carry[4]), .Y(n34) );
  XOR2XL U16 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  INVX2 U17 ( .A(n37), .Y(n48) );
  XOR2X1 U18 ( .A(B[4]), .B(A[4]), .Y(n44) );
  XOR2X1 U19 ( .A(A[6]), .B(B[6]), .Y(n33) );
  XOR2X1 U20 ( .A(carry[30]), .B(n36), .Y(SUM[30]) );
  INVX1 U21 ( .A(n32), .Y(n49) );
  XOR2X1 U22 ( .A(n43), .B(n44), .Y(SUM[4]) );
  XOR2X1 U23 ( .A(carry[15]), .B(n42), .Y(SUM[15]) );
  XOR2X1 U24 ( .A(carry[22]), .B(n38), .Y(SUM[22]) );
  XOR2X1 U25 ( .A(carry[19]), .B(n40), .Y(SUM[19]) );
  XOR2X1 U26 ( .A(carry[6]), .B(n33), .Y(SUM[6]) );
  XOR2X1 U27 ( .A(A[15]), .B(B[15]), .Y(n42) );
  XOR2X1 U28 ( .A(A[19]), .B(B[19]), .Y(n40) );
  XOR2X1 U29 ( .A(A[22]), .B(B[22]), .Y(n38) );
  XOR2X1 U30 ( .A(A[30]), .B(B[30]), .Y(n36) );
  OAI2BB1X1 U31 ( .A0N(A[3]), .A1N(B[3]), .B0(n45), .Y(n43) );
  OAI21XL U32 ( .A0(A[3]), .A1(B[3]), .B0(carry[3]), .Y(n45) );
endmodule


module hash_core_DW01_add_5 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n21, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47;
  wire   [31:2] carry;

  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CMPR32X1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX4 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(n21), .CO(carry[16]), .S(SUM[15])
         );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  OAI21X4 U1 ( .A0(A[14]), .A1(B[14]), .B0(carry[14]), .Y(n28) );
  OAI2BB1X4 U2 ( .A0N(A[14]), .A1N(B[14]), .B0(n28), .Y(n21) );
  OAI2BB1X4 U3 ( .A0N(A[18]), .A1N(B[18]), .B0(n31), .Y(carry[19]) );
  OAI21X2 U4 ( .A0(A[5]), .A1(B[5]), .B0(carry[5]), .Y(n29) );
  OAI211X2 U5 ( .A0(A[1]), .A1(B[1]), .B0(A[0]), .C0(B[0]), .Y(n30) );
  OAI2BB1X2 U6 ( .A0N(A[9]), .A1N(B[9]), .B0(n32), .Y(carry[10]) );
  OAI21X2 U7 ( .A0(A[9]), .A1(B[9]), .B0(carry[9]), .Y(n32) );
  OAI2BB1X4 U8 ( .A0N(A[16]), .A1N(B[16]), .B0(n44), .Y(carry[17]) );
  OAI21X4 U9 ( .A0(A[16]), .A1(B[16]), .B0(carry[16]), .Y(n44) );
  OAI21X4 U10 ( .A0(A[18]), .A1(B[18]), .B0(carry[18]), .Y(n31) );
  AND2X1 U11 ( .A(A[0]), .B(B[0]), .Y(n39) );
  XOR2XL U12 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  OAI2BB1X2 U13 ( .A0N(A[1]), .A1N(B[1]), .B0(n30), .Y(carry[2]) );
  XOR2XL U14 ( .A(B[1]), .B(A[1]), .Y(n40) );
  XOR2XL U15 ( .A(B[9]), .B(A[9]), .Y(n34) );
  AOI22XL U16 ( .A0(B[17]), .A1(n43), .B0(A[17]), .B1(carry[17]), .Y(n42) );
  OR2XL U17 ( .A(carry[17]), .B(A[17]), .Y(n43) );
  XOR2X1 U18 ( .A(B[5]), .B(A[5]), .Y(n37) );
  OAI2BB1X1 U19 ( .A0N(A[5]), .A1N(B[5]), .B0(n29), .Y(carry[6]) );
  XOR2X1 U20 ( .A(n33), .B(n34), .Y(SUM[9]) );
  XOR2X1 U21 ( .A(n36), .B(n37), .Y(SUM[5]) );
  XOR2X1 U22 ( .A(n41), .B(n42), .Y(SUM[18]) );
  XOR2X1 U23 ( .A(n39), .B(n40), .Y(SUM[1]) );
  XOR2X1 U24 ( .A(n45), .B(n46), .Y(SUM[16]) );
  XOR2X1 U25 ( .A(B[16]), .B(A[16]), .Y(n46) );
  OAI2BB1X1 U26 ( .A0N(A[15]), .A1N(B[15]), .B0(n47), .Y(n45) );
  OAI21XL U27 ( .A0(A[15]), .A1(B[15]), .B0(carry[15]), .Y(n47) );
  OAI2BB1X1 U28 ( .A0N(A[8]), .A1N(B[8]), .B0(n35), .Y(n33) );
  OAI21XL U29 ( .A0(A[8]), .A1(B[8]), .B0(carry[8]), .Y(n35) );
  OAI2BB1X1 U30 ( .A0N(A[4]), .A1N(B[4]), .B0(n38), .Y(n36) );
  OAI21XL U31 ( .A0(A[4]), .A1(B[4]), .B0(carry[4]), .Y(n38) );
  XNOR2X1 U32 ( .A(A[18]), .B(B[18]), .Y(n41) );
endmodule


module hash_core_DW01_add_6 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n47, n46, n48, n49, n50, n51, n52, n53, n54, n55;
  wire   [31:2] carry;

  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  INVX1 U1 ( .A(B[18]), .Y(n49) );
  OAI21X1 U2 ( .A0(A[4]), .A1(B[4]), .B0(carry[4]), .Y(n36) );
  INVXL U3 ( .A(A[18]), .Y(n48) );
  DLY1X1 U4 ( .A(n43), .Y(n46) );
  OAI2BB1X4 U5 ( .A0N(n48), .A1N(n49), .B0(carry[18]), .Y(n31) );
  OAI2BB1X4 U6 ( .A0N(A[16]), .A1N(B[16]), .B0(n43), .Y(carry[17]) );
  OAI2BB1X4 U7 ( .A0N(A[18]), .A1N(B[18]), .B0(n31), .Y(carry[19]) );
  OAI21X4 U8 ( .A0(A[16]), .A1(B[16]), .B0(carry[16]), .Y(n43) );
  NAND2X2 U9 ( .A(n50), .B(n51), .Y(n52) );
  NAND2X4 U10 ( .A(n52), .B(carry[10]), .Y(n32) );
  INVXL U11 ( .A(A[10]), .Y(n50) );
  INVX1 U12 ( .A(B[10]), .Y(n51) );
  OAI2BB1X4 U13 ( .A0N(A[10]), .A1N(B[10]), .B0(n32), .Y(carry[11]) );
  AND2X1 U14 ( .A(A[0]), .B(B[0]), .Y(n38) );
  XOR2XL U15 ( .A(B[1]), .B(A[1]), .Y(n39) );
  OAI2BB1X4 U16 ( .A0N(A[1]), .A1N(B[1]), .B0(n30), .Y(carry[2]) );
  OAI21X2 U17 ( .A0(A[6]), .A1(B[6]), .B0(carry[6]), .Y(n29) );
  OAI2BB1X1 U18 ( .A0N(A[4]), .A1N(B[4]), .B0(n36), .Y(carry[5]) );
  XNOR2X1 U19 ( .A(n45), .B(n53), .Y(SUM[10]) );
  XNOR2XL U20 ( .A(B[10]), .B(A[10]), .Y(n53) );
  XNOR2XL U21 ( .A(A[6]), .B(B[6]), .Y(n33) );
  OAI2BB1XL U22 ( .A0N(A[4]), .A1N(B[4]), .B0(n36), .Y(n54) );
  OAI2BB1XL U23 ( .A0N(A[16]), .A1N(B[16]), .B0(n46), .Y(n55) );
  OAI211X2 U24 ( .A0(A[1]), .A1(B[1]), .B0(A[0]), .C0(B[0]), .Y(n30) );
  OAI2BB1X1 U25 ( .A0N(A[6]), .A1N(B[6]), .B0(n29), .Y(carry[7]) );
  XOR2X1 U26 ( .A(A[16]), .B(n44), .Y(SUM[16]) );
  XOR2X1 U27 ( .A(carry[16]), .B(B[16]), .Y(n44) );
  XOR2X1 U28 ( .A(n40), .B(n41), .Y(SUM[18]) );
  XOR2X1 U29 ( .A(n38), .B(n39), .Y(SUM[1]) );
  XOR2X1 U30 ( .A(A[4]), .B(n37), .Y(SUM[4]) );
  XOR2X1 U31 ( .A(carry[4]), .B(B[4]), .Y(n37) );
  AOI22XL U32 ( .A0(B[17]), .A1(n42), .B0(A[17]), .B1(n55), .Y(n41) );
  OR2XL U33 ( .A(n55), .B(A[17]), .Y(n42) );
  OAI2BB1X1 U34 ( .A0N(A[9]), .A1N(B[9]), .B0(n47), .Y(n45) );
  OAI21XL U35 ( .A0(A[9]), .A1(B[9]), .B0(carry[9]), .Y(n47) );
  XOR2X1 U36 ( .A(n33), .B(n34), .Y(SUM[6]) );
  AOI22XL U37 ( .A0(B[5]), .A1(n35), .B0(A[5]), .B1(n54), .Y(n34) );
  OR2XL U38 ( .A(n54), .B(A[5]), .Y(n35) );
  XNOR2X1 U39 ( .A(A[18]), .B(B[18]), .Y(n40) );
  XOR2XL U40 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module hash_core_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module hash_core_DW01_add_16 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n318,
         n319, n320, n321, n325, n326, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n349, n350, n351, n352, n353, n356, n357, n358,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n372, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n316, n317, n322, n323, n324, n327, n348, n354,
         n355, n359, n371, n373, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451;

  OAI211X2 U38 ( .A0(n334), .A1(n433), .B0(n335), .C0(n336), .Y(n331) );
  OAI221X2 U39 ( .A0(B[26]), .A1(A[26]), .B0(A[27]), .B1(B[27]), .C0(n337), 
        .Y(n336) );
  OR2X4 U42 ( .A(A[28]), .B(B[28]), .Y(n332) );
  OAI2BB1X4 U50 ( .A0N(n342), .A1N(n431), .B0(B[25]), .Y(n344) );
  OAI211X2 U51 ( .A0(A[25]), .A1(B[25]), .B0(n345), .C0(n346), .Y(n343) );
  OAI211X2 U58 ( .A0(n430), .A1(n350), .B0(n351), .C0(n352), .Y(n345) );
  OAI2BB1X4 U60 ( .A0N(n350), .A1N(n430), .B0(B[23]), .Y(n351) );
  OR2X4 U62 ( .A(A[24]), .B(B[24]), .Y(n346) );
  NAND2X4 U63 ( .A(B[24]), .B(A[24]), .Y(n342) );
  OAI2BB1X4 U70 ( .A0N(n358), .A1N(n429), .B0(B[21]), .Y(n360) );
  NAND2X4 U73 ( .A(B[22]), .B(A[22]), .Y(n350) );
  AOI211X2 U78 ( .A0(n366), .A1(A[19]), .B0(n368), .C0(n367), .Y(n364) );
  AOI2BB1X4 U80 ( .A0N(n366), .A1N(A[19]), .B0(n448), .Y(n367) );
  NAND2X4 U83 ( .A(B[20]), .B(A[20]), .Y(n358) );
  AOI21X4 U91 ( .A0(n376), .A1(n425), .B0(n377), .Y(n369) );
  NOR2X4 U93 ( .A(n447), .B(n426), .Y(n366) );
  AND2X2 U96 ( .A(B[17]), .B(A[17]), .Y(n377) );
  NOR2X4 U97 ( .A(B[17]), .B(A[17]), .Y(n378) );
  OAI21X4 U98 ( .A0(n380), .A1(n381), .B0(n382), .Y(n376) );
  OAI21X4 U101 ( .A0(B[15]), .A1(A[15]), .B0(n385), .Y(n384) );
  AOI31X2 U102 ( .A0(n386), .A1(n388), .A2(n387), .B0(n389), .Y(n385) );
  OAI222X2 U103 ( .A0(B[12]), .A1(A[12]), .B0(n390), .B1(n439), .C0(B[13]), 
        .C1(A[13]), .Y(n388) );
  NAND2X4 U105 ( .A(B[16]), .B(A[16]), .Y(n382) );
  NOR2X4 U106 ( .A(B[16]), .B(A[16]), .Y(n381) );
  NAND2X4 U115 ( .A(B[14]), .B(A[14]), .Y(n387) );
  AOI2BB2X4 U126 ( .B0(n450), .B1(n440), .A0N(A[10]), .A1N(B[10]), .Y(n404) );
  NAND2X4 U139 ( .A(B[8]), .B(A[8]), .Y(n298) );
  OAI32X4 U141 ( .A0(n415), .A1(n302), .A2(n311), .B0(n416), .B1(n302), .Y(
        n296) );
  AOI211X2 U142 ( .A0(n417), .A1(n418), .B0(n445), .C0(n301), .Y(n416) );
  AND2X2 U143 ( .A(B[7]), .B(A[7]), .Y(n301) );
  NAND2BX4 U145 ( .AN(n309), .B(n313), .Y(n418) );
  NAND2X4 U146 ( .A(B[4]), .B(A[4]), .Y(n313) );
  NOR2X4 U147 ( .A(n449), .B(n444), .Y(n309) );
  AOI21X4 U148 ( .A0(n315), .A1(A[3]), .B0(n442), .Y(n311) );
  AOI2BB1X4 U150 ( .A0N(A[2]), .A1N(n328), .B0(n420), .Y(n315) );
  AOI21X4 U151 ( .A0(n328), .A1(A[2]), .B0(B[2]), .Y(n420) );
  OAI2BB1X4 U152 ( .A0N(n370), .A1N(A[1]), .B0(n421), .Y(n328) );
  OAI21X4 U153 ( .A0(n370), .A1(A[1]), .B0(B[1]), .Y(n421) );
  OAI21X4 U155 ( .A0(B[4]), .A1(A[4]), .B0(n417), .Y(n415) );
  AOI21X4 U156 ( .A0(n449), .A1(n444), .B0(n303), .Y(n417) );
  NOR2X4 U157 ( .A(A[6]), .B(B[6]), .Y(n303) );
  NOR2X4 U161 ( .A(n451), .B(n443), .Y(n370) );
  INVX4 U2 ( .A(n405), .Y(n286) );
  OAI21X2 U3 ( .A0(n434), .A1(n326), .B0(n267), .Y(n325) );
  NAND2X2 U4 ( .A(n267), .B(n321), .Y(n329) );
  OAI21X2 U5 ( .A0(B[8]), .A1(A[8]), .B0(n404), .Y(n401) );
  XNOR2XL U6 ( .A(B[19]), .B(A[19]), .Y(n372) );
  XNOR2X2 U7 ( .A(B[23]), .B(A[23]), .Y(n327) );
  INVX8 U8 ( .A(A[23]), .Y(n430) );
  AOI2BB1XL U9 ( .A0N(n270), .A1N(n271), .B0(n436), .Y(n264) );
  INVX8 U10 ( .A(n384), .Y(n436) );
  OAI21XL U11 ( .A0(n264), .A1(n381), .B0(n382), .Y(n265) );
  NAND2X4 U12 ( .A(n430), .B(n266), .Y(n317) );
  CLKINVX20 U13 ( .A(B[23]), .Y(n266) );
  OAI211X1 U14 ( .A0(n350), .A1(n430), .B0(n268), .C0(n351), .Y(n291) );
  INVX8 U15 ( .A(A[18]), .Y(n426) );
  OR2X4 U16 ( .A(A[29]), .B(B[29]), .Y(n267) );
  INVX4 U17 ( .A(n334), .Y(n432) );
  DLY1X1 U18 ( .A(n352), .Y(n268) );
  DLY1X1 U19 ( .A(A[10]), .Y(n269) );
  AOI2BB1X4 U20 ( .A0N(n270), .A1N(n271), .B0(n436), .Y(n380) );
  CLKINVX20 U21 ( .A(A[15]), .Y(n270) );
  CLKINVX20 U22 ( .A(B[15]), .Y(n271) );
  DLY1X1 U23 ( .A(A[9]), .Y(n272) );
  INVX8 U24 ( .A(A[21]), .Y(n429) );
  NAND2X4 U25 ( .A(B[12]), .B(A[12]), .Y(n399) );
  OAI211X2 U26 ( .A0(B[21]), .A1(A[21]), .B0(n424), .C0(n428), .Y(n273) );
  INVX4 U27 ( .A(n363), .Y(n428) );
  NOR2X4 U28 ( .A(A[20]), .B(B[20]), .Y(n363) );
  INVX4 U29 ( .A(n296), .Y(n441) );
  INVX1 U30 ( .A(B[29]), .Y(n281) );
  INVX1 U31 ( .A(B[26]), .Y(n276) );
  OAI21X2 U32 ( .A0(n315), .A1(A[3]), .B0(B[3]), .Y(n419) );
  XOR2X1 U33 ( .A(n391), .B(n392), .Y(SUM[15]) );
  XNOR2XL U34 ( .A(n333), .B(n331), .Y(SUM[28]) );
  OAI211X4 U35 ( .A0(n358), .A1(n429), .B0(n360), .C0(n273), .Y(n282) );
  DLY1X1 U36 ( .A(n343), .Y(n290) );
  NAND2X2 U37 ( .A(n330), .B(n332), .Y(n333) );
  INVX4 U40 ( .A(n399), .Y(n439) );
  INVX1 U41 ( .A(n322), .Y(n274) );
  DLY1X1 U43 ( .A(n369), .Y(n275) );
  AOI21X4 U44 ( .A0(n340), .A1(n292), .B0(n277), .Y(n339) );
  NAND2BX4 U45 ( .AN(n276), .B(A[26]), .Y(n334) );
  DLY1X1 U46 ( .A(n432), .Y(n277) );
  INVXL U47 ( .A(n284), .Y(n278) );
  DLY1X1 U48 ( .A(n264), .Y(n279) );
  DLY1X1 U49 ( .A(n265), .Y(n280) );
  NAND2BX4 U52 ( .AN(n434), .B(n321), .Y(n289) );
  NAND2BX4 U53 ( .AN(n281), .B(A[29]), .Y(n321) );
  XOR2X2 U54 ( .A(n320), .B(n329), .Y(SUM[29]) );
  XOR2X4 U55 ( .A(n338), .B(n339), .Y(SUM[27]) );
  NAND2X2 U56 ( .A(n325), .B(n321), .Y(n323) );
  AND2X1 U57 ( .A(B[11]), .B(n278), .Y(n406) );
  NAND2X2 U59 ( .A(A[10]), .B(B[10]), .Y(n407) );
  OAI221X2 U61 ( .A0(n285), .A1(n286), .B0(n284), .B1(n283), .C0(n407), .Y(
        n287) );
  INVX1 U64 ( .A(B[11]), .Y(n283) );
  INVX4 U65 ( .A(A[11]), .Y(n284) );
  INVX4 U66 ( .A(n404), .Y(n285) );
  INVX4 U67 ( .A(n287), .Y(n403) );
  XNOR2X4 U68 ( .A(n318), .B(n288), .Y(SUM[31]) );
  XOR2X4 U69 ( .A(A[31]), .B(B[31]), .Y(n288) );
  OAI211X2 U71 ( .A0(n358), .A1(n429), .B0(n273), .C0(n360), .Y(n353) );
  CLKINVX8 U72 ( .A(A[30]), .Y(n435) );
  INVX4 U74 ( .A(n364), .Y(n424) );
  NAND2X4 U75 ( .A(n435), .B(n446), .Y(n294) );
  INVX8 U76 ( .A(A[25]), .Y(n431) );
  OAI211X2 U77 ( .A0(n342), .A1(n431), .B0(n290), .C0(n344), .Y(n292) );
  XNOR2X2 U79 ( .A(n341), .B(n292), .Y(SUM[26]) );
  OR2X4 U81 ( .A(n326), .B(n289), .Y(n293) );
  INVXL U82 ( .A(A[27]), .Y(n433) );
  NOR2X1 U84 ( .A(n434), .B(n326), .Y(n320) );
  INVX8 U85 ( .A(n330), .Y(n434) );
  AOI2BB1X4 U86 ( .A0N(n446), .A1N(n435), .B0(n319), .Y(n318) );
  OAI21X2 U87 ( .A0(n432), .A1(A[27]), .B0(B[27]), .Y(n335) );
  NAND3X4 U88 ( .A(n353), .B(n317), .C(n316), .Y(n352) );
  AND3X4 U89 ( .A(n293), .B(n294), .C(n267), .Y(n319) );
  OR2X2 U90 ( .A(B[22]), .B(A[22]), .Y(n316) );
  OAI211X2 U92 ( .A0(n342), .A1(n431), .B0(n343), .C0(n344), .Y(n337) );
  INVXL U94 ( .A(n424), .Y(n322) );
  INVX8 U95 ( .A(A[9]), .Y(n440) );
  OAI32X2 U99 ( .A0(n401), .A1(n441), .A2(n402), .B0(n403), .B1(n402), .Y(n390) );
  INVX4 U100 ( .A(A[0]), .Y(n443) );
  INVX8 U104 ( .A(A[5]), .Y(n444) );
  XNOR2X4 U107 ( .A(n323), .B(n373), .Y(SUM[30]) );
  INVX4 U108 ( .A(n378), .Y(n425) );
  CLKINVX4 U109 ( .A(n305), .Y(n445) );
  INVXL U110 ( .A(n389), .Y(n438) );
  NAND2X4 U111 ( .A(B[28]), .B(A[28]), .Y(n330) );
  XOR2X1 U112 ( .A(n347), .B(n324), .Y(SUM[25]) );
  XNOR2XL U113 ( .A(B[25]), .B(n431), .Y(n324) );
  XNOR2X1 U114 ( .A(n327), .B(n422), .Y(SUM[23]) );
  XNOR2X1 U116 ( .A(n372), .B(n348), .Y(SUM[19]) );
  OR2XL U117 ( .A(n374), .B(n366), .Y(n348) );
  AOI21X1 U118 ( .A0(n393), .A1(n438), .B0(n437), .Y(n392) );
  XOR2XL U119 ( .A(n354), .B(n295), .Y(SUM[9]) );
  XOR2X1 U120 ( .A(n272), .B(B[9]), .Y(n354) );
  XNOR2X1 U121 ( .A(n315), .B(n355), .Y(SUM[3]) );
  XNOR2XL U122 ( .A(B[3]), .B(A[3]), .Y(n355) );
  XOR2XL U123 ( .A(n359), .B(n328), .Y(SUM[2]) );
  XOR2X1 U124 ( .A(A[2]), .B(B[2]), .Y(n359) );
  XNOR2X1 U125 ( .A(n370), .B(n371), .Y(SUM[1]) );
  XNOR2XL U127 ( .A(B[1]), .B(A[1]), .Y(n371) );
  OAI21X2 U128 ( .A0(n450), .A1(n440), .B0(n298), .Y(n405) );
  XOR2X2 U129 ( .A(A[30]), .B(n446), .Y(n373) );
  NAND2XL U130 ( .A(n342), .B(n346), .Y(n349) );
  AOI21XL U131 ( .A0(n447), .A1(n426), .B0(n366), .Y(n375) );
  XNOR2XL U132 ( .A(n365), .B(n274), .Y(SUM[20]) );
  NAND2XL U133 ( .A(n358), .B(n428), .Y(n365) );
  XNOR2X1 U134 ( .A(n394), .B(n393), .Y(SUM[14]) );
  NAND2XL U135 ( .A(n387), .B(n438), .Y(n394) );
  XOR2X1 U136 ( .A(n280), .B(n379), .Y(SUM[17]) );
  NOR2XL U137 ( .A(n378), .B(n377), .Y(n379) );
  XOR2XL U138 ( .A(n383), .B(n279), .Y(SUM[16]) );
  NAND2BXL U140 ( .AN(n381), .B(n382), .Y(n383) );
  AOI21XL U144 ( .A0(n295), .A1(n272), .B0(n413), .Y(n410) );
  AOI2BB1X1 U149 ( .A0N(n272), .A1N(n295), .B0(n450), .Y(n413) );
  AOI21XL U154 ( .A0(n307), .A1(n308), .B0(n309), .Y(n304) );
  NAND2XL U158 ( .A(n444), .B(n449), .Y(n308) );
  XOR2X1 U159 ( .A(n299), .B(n300), .Y(SUM[7]) );
  NOR2XL U160 ( .A(n301), .B(n302), .Y(n300) );
  OAI21XL U162 ( .A0(n303), .A1(n304), .B0(n305), .Y(n299) );
  XOR2X1 U163 ( .A(n307), .B(n310), .Y(SUM[5]) );
  AOI21XL U164 ( .A0(n444), .A1(n449), .B0(n309), .Y(n310) );
  XOR2X1 U165 ( .A(n306), .B(n304), .Y(SUM[6]) );
  NAND2BXL U166 ( .AN(n303), .B(n305), .Y(n306) );
  AOI21XL U167 ( .A0(n451), .A1(n443), .B0(n370), .Y(SUM[0]) );
  INVX1 U168 ( .A(B[19]), .Y(n448) );
  NOR2X2 U169 ( .A(A[7]), .B(B[7]), .Y(n302) );
  NAND2X2 U170 ( .A(B[13]), .B(A[13]), .Y(n386) );
  NAND2X2 U171 ( .A(B[6]), .B(A[6]), .Y(n305) );
  NOR2X2 U172 ( .A(A[14]), .B(B[14]), .Y(n389) );
  OAI21XL U173 ( .A0(B[22]), .A1(A[22]), .B0(n350), .Y(n357) );
  OAI21XL U174 ( .A0(B[26]), .A1(A[26]), .B0(n334), .Y(n341) );
  XNOR2XL U175 ( .A(A[27]), .B(B[27]), .Y(n338) );
  OR2XL U176 ( .A(A[26]), .B(B[26]), .Y(n340) );
  NAND2XL U177 ( .A(n356), .B(n350), .Y(n422) );
  OR2XL U178 ( .A(A[12]), .B(B[12]), .Y(n398) );
  OAI21XL U179 ( .A0(n395), .A1(n396), .B0(n386), .Y(n393) );
  NOR2XL U180 ( .A(A[13]), .B(B[13]), .Y(n396) );
  INVX1 U181 ( .A(B[0]), .Y(n451) );
  XOR2X1 U182 ( .A(n397), .B(n395), .Y(SUM[13]) );
  OAI21XL U183 ( .A0(B[13]), .A1(A[13]), .B0(n386), .Y(n397) );
  XOR2X2 U184 ( .A(n361), .B(n362), .Y(SUM[21]) );
  XNOR2XL U185 ( .A(B[21]), .B(n429), .Y(n362) );
  XNOR2X1 U186 ( .A(A[15]), .B(B[15]), .Y(n391) );
  INVXL U187 ( .A(n387), .Y(n437) );
  OAI21XL U188 ( .A0(n441), .A1(n414), .B0(n298), .Y(n295) );
  NOR2XL U189 ( .A(A[8]), .B(B[8]), .Y(n414) );
  INVX1 U190 ( .A(B[5]), .Y(n449) );
  OAI21XL U191 ( .A0(B[12]), .A1(A[12]), .B0(n399), .Y(n400) );
  XOR2X1 U192 ( .A(n408), .B(n409), .Y(SUM[11]) );
  NOR2XL U193 ( .A(n406), .B(n402), .Y(n409) );
  OAI21XL U194 ( .A0(n410), .A1(n411), .B0(n407), .Y(n408) );
  NOR2XL U195 ( .A(n269), .B(B[10]), .Y(n411) );
  XOR2X1 U196 ( .A(n412), .B(n410), .Y(SUM[10]) );
  OAI21XL U197 ( .A0(B[10]), .A1(n269), .B0(n407), .Y(n412) );
  INVX1 U198 ( .A(B[9]), .Y(n450) );
  XNOR2X1 U199 ( .A(n296), .B(n297), .Y(SUM[8]) );
  OAI21XL U200 ( .A0(A[8]), .A1(B[8]), .B0(n298), .Y(n297) );
  OAI21XL U201 ( .A0(n311), .A1(n312), .B0(n313), .Y(n307) );
  NOR2XL U202 ( .A(A[4]), .B(B[4]), .Y(n312) );
  XOR2XL U203 ( .A(n314), .B(n311), .Y(SUM[4]) );
  OAI21XL U204 ( .A0(B[4]), .A1(A[4]), .B0(n313), .Y(n314) );
  INVX1 U205 ( .A(B[18]), .Y(n447) );
  INVX1 U206 ( .A(B[30]), .Y(n446) );
  AOI21XL U207 ( .A0(n447), .A1(n426), .B0(n275), .Y(n374) );
  XNOR2XL U208 ( .A(n375), .B(n275), .Y(SUM[18]) );
  OAI21XL U209 ( .A0(n363), .A1(n322), .B0(n358), .Y(n361) );
  OAI2BB1X1 U210 ( .A0N(n346), .A1N(n291), .B0(n342), .Y(n347) );
  XNOR2XL U211 ( .A(n349), .B(n291), .Y(SUM[24]) );
  DLY1X1 U212 ( .A(n390), .Y(n423) );
  INVX3 U213 ( .A(A[19]), .Y(n427) );
  XNOR2XL U214 ( .A(n357), .B(n282), .Y(SUM[22]) );
  XNOR2XL U215 ( .A(n400), .B(n423), .Y(SUM[12]) );
  OAI21XL U216 ( .A0(B[22]), .A1(A[22]), .B0(n282), .Y(n356) );
  AOI21XL U217 ( .A0(n423), .A1(n398), .B0(n439), .Y(n395) );
  NOR2X2 U218 ( .A(A[11]), .B(B[11]), .Y(n402) );
  AOI221X2 U219 ( .A0(n447), .A1(n426), .B0(n448), .B1(n427), .C0(n369), .Y(
        n368) );
  AND2X4 U220 ( .A(n331), .B(n332), .Y(n326) );
  CLKINVX4 U221 ( .A(n419), .Y(n442) );
endmodule


module hash_core_DW01_add_25 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n451, n452, n453, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n305, n306, n307, n308,
         n309, n310, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n333,
         n334, n336, n337, n339, n340, n341, n343, n344, n345, n346, n347,
         n348, n349, n350, n352, n353, n354, n355, n356, n358, n359, n361,
         n362, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n304, n311, n331, n332,
         n335, n338, n342, n351, n357, n360, n363, n388, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n418, n419, n420,
         n422, n423, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450;

  XOR2X4 U6 ( .A(n297), .B(n298), .Y(SUM[7]) );
  XOR2X4 U18 ( .A(n313), .B(n314), .Y(SUM[31]) );
  OAI21X4 U30 ( .A0(n327), .A1(n326), .B0(n328), .Y(n318) );
  NAND2BX4 U34 ( .AN(n326), .B(n328), .Y(n329) );
  AOI2BB1X4 U39 ( .A0N(A[26]), .A1N(n406), .B0(n334), .Y(n330) );
  AOI21X4 U46 ( .A0(n339), .A1(n439), .B0(n340), .Y(n336) );
  NOR2X4 U51 ( .A(B[24]), .B(A[24]), .Y(n341) );
  OAI2BB1X4 U52 ( .A0N(A[23]), .A1N(n343), .B0(n344), .Y(n339) );
  OAI21X4 U53 ( .A0(n343), .A1(A[23]), .B0(B[23]), .Y(n344) );
  AOI2BB1X4 U56 ( .A0N(n346), .A1N(A[22]), .B0(n347), .Y(n343) );
  AOI21X4 U57 ( .A0(n346), .A1(A[22]), .B0(B[22]), .Y(n347) );
  OAI2BB1X4 U60 ( .A0N(A[21]), .A1N(n349), .B0(n350), .Y(n346) );
  OAI21X4 U61 ( .A0(n349), .A1(A[21]), .B0(B[21]), .Y(n350) );
  OAI21X4 U64 ( .A0(n353), .A1(n352), .B0(n354), .Y(n349) );
  NAND2X4 U69 ( .A(B[20]), .B(A[20]), .Y(n354) );
  NOR2X4 U70 ( .A(B[20]), .B(A[20]), .Y(n352) );
  OAI2BB1X4 U74 ( .A0N(A[18]), .A1N(n361), .B0(n362), .Y(n356) );
  OAI21X4 U75 ( .A0(n361), .A1(A[18]), .B0(n282), .Y(n362) );
  OAI2BB1X4 U79 ( .A0N(A[17]), .A1N(n364), .B0(n365), .Y(n361) );
  OAI21X4 U80 ( .A0(n364), .A1(A[17]), .B0(B[17]), .Y(n365) );
  NAND2X4 U83 ( .A(n367), .B(n368), .Y(n364) );
  AOI31X2 U88 ( .A0(n374), .A1(n375), .A2(n376), .B0(n377), .Y(n373) );
  OAI211X2 U89 ( .A0(B[13]), .A1(A[13]), .B0(n378), .C0(n437), .Y(n374) );
  XOR2X4 U92 ( .A(n379), .B(n380), .Y(SUM[15]) );
  NOR2X4 U94 ( .A(n438), .B(n445), .Y(n370) );
  XOR2X4 U96 ( .A(n382), .B(n381), .Y(SUM[14]) );
  AND2X2 U97 ( .A(n383), .B(n376), .Y(n381) );
  NAND2X4 U100 ( .A(B[14]), .B(A[14]), .Y(n375) );
  NOR2X4 U101 ( .A(A[14]), .B(B[14]), .Y(n377) );
  NAND2X4 U104 ( .A(B[13]), .B(A[13]), .Y(n376) );
  XOR2X4 U114 ( .A(n397), .B(n398), .Y(SUM[11]) );
  NAND2X4 U124 ( .A(B[9]), .B(A[9]), .Y(n292) );
  NAND2X4 U126 ( .A(B[8]), .B(A[8]), .Y(n295) );
  NAND2BX4 U127 ( .AN(n293), .B(n296), .Y(n394) );
  OR2X4 U128 ( .A(B[8]), .B(A[8]), .Y(n296) );
  OAI31X2 U129 ( .A0(n401), .A1(n300), .A2(n302), .B0(n303), .Y(n293) );
  NOR2X4 U131 ( .A(n441), .B(n447), .Y(n302) );
  AND2X2 U132 ( .A(B[6]), .B(A[6]), .Y(n300) );
  NOR2X4 U134 ( .A(B[6]), .B(A[6]), .Y(n301) );
  OAI21X4 U138 ( .A0(n310), .A1(A[4]), .B0(B[4]), .Y(n402) );
  OAI21X4 U139 ( .A0(n276), .A1(n448), .B0(n403), .Y(n310) );
  OAI2BB1X4 U140 ( .A0N(n357), .A1N(n448), .B0(B[3]), .Y(n403) );
  NOR2X4 U142 ( .A(A[2]), .B(B[2]), .Y(n320) );
  NAND2BX4 U143 ( .AN(n324), .B(n323), .Y(n321) );
  NAND2X4 U144 ( .A(B[2]), .B(A[2]), .Y(n323) );
  OAI2BB1X4 U145 ( .A0N(n358), .A1N(A[1]), .B0(n404), .Y(n324) );
  NOR2X4 U149 ( .A(n442), .B(n449), .Y(n358) );
  DLY1X1 U2 ( .A(n396), .Y(n268) );
  DLY1X1 U3 ( .A(n411), .Y(n278) );
  AOI211X1 U4 ( .A0(n306), .A1(n307), .B0(n305), .C0(n301), .Y(n269) );
  DLY1X1 U5 ( .A(n291), .Y(n270) );
  NOR2X4 U7 ( .A(B[10]), .B(A[10]), .Y(n271) );
  NOR2XL U8 ( .A(B[10]), .B(A[10]), .Y(n272) );
  OAI31X4 U9 ( .A0(n269), .A1(n300), .A2(n302), .B0(n303), .Y(n273) );
  NOR2BX4 U10 ( .AN(n274), .B(B[9]), .Y(n291) );
  CLKINVX20 U11 ( .A(A[9]), .Y(n274) );
  OAI33X4 U12 ( .A0(n394), .A1(n272), .A2(n270), .B0(n268), .B1(n272), .B2(
        n291), .Y(n275) );
  NAND2X4 U13 ( .A(n321), .B(n444), .Y(n276) );
  NAND2XL U14 ( .A(B[12]), .B(A[12]), .Y(n277) );
  XOR2X2 U15 ( .A(n430), .B(n351), .Y(SUM[19]) );
  NAND2X4 U16 ( .A(n279), .B(n316), .Y(n315) );
  CLKINVX20 U17 ( .A(n281), .Y(n279) );
  XNOR2X2 U19 ( .A(n330), .B(n427), .Y(n451) );
  NAND2BX4 U20 ( .AN(n280), .B(B[5]), .Y(n307) );
  CLKINVX20 U21 ( .A(A[5]), .Y(n280) );
  CLKINVX20 U22 ( .A(A[30]), .Y(n281) );
  INVX1 U23 ( .A(A[19]), .Y(n412) );
  INVX2 U24 ( .A(A[3]), .Y(n448) );
  INVX1 U25 ( .A(A[15]), .Y(n445) );
  INVX4 U26 ( .A(B[0]), .Y(n442) );
  BUFX8 U27 ( .A(n451), .Y(SUM[27]) );
  CLKINVX3 U28 ( .A(n432), .Y(SUM[25]) );
  XOR2X2 U29 ( .A(n327), .B(n329), .Y(SUM[28]) );
  INVX1 U31 ( .A(n271), .Y(n436) );
  XNOR2X2 U32 ( .A(n316), .B(n317), .Y(SUM[30]) );
  NOR2X4 U33 ( .A(A[5]), .B(B[5]), .Y(n305) );
  BUFX8 U35 ( .A(B[18]), .Y(n282) );
  NOR2X4 U36 ( .A(B[10]), .B(A[10]), .Y(n283) );
  AND2X4 U37 ( .A(B[24]), .B(A[24]), .Y(n340) );
  OAI21X1 U38 ( .A0(A[13]), .A1(B[13]), .B0(n376), .Y(n385) );
  OAI21X1 U40 ( .A0(A[13]), .A1(B[13]), .B0(n384), .Y(n383) );
  OAI2BB1X4 U41 ( .A0N(n444), .A1N(n323), .B0(n324), .Y(n322) );
  NAND2X4 U42 ( .A(n321), .B(n444), .Y(n357) );
  INVX4 U43 ( .A(B[16]), .Y(n288) );
  XOR2X1 U44 ( .A(n423), .B(n406), .Y(n422) );
  NAND2BX2 U45 ( .AN(n352), .B(n354), .Y(n355) );
  INVX8 U47 ( .A(n434), .Y(n306) );
  XNOR2X2 U48 ( .A(A[26]), .B(B[26]), .Y(n423) );
  AOI21X4 U49 ( .A0(n284), .A1(n285), .B0(n286), .Y(n287) );
  INVX4 U50 ( .A(n381), .Y(n284) );
  INVXL U54 ( .A(n377), .Y(n285) );
  INVXL U55 ( .A(n375), .Y(n286) );
  INVX4 U58 ( .A(n287), .Y(n379) );
  OAI2BB2X4 U59 ( .B0(n369), .B1(n370), .A0N(n288), .A1N(n409), .Y(n367) );
  INVX1 U62 ( .A(A[16]), .Y(n409) );
  AOI21X4 U63 ( .A0(n277), .A1(n304), .B0(n389), .Y(n311) );
  INVXL U65 ( .A(n386), .Y(n304) );
  INVX4 U66 ( .A(n311), .Y(n387) );
  OAI2BB1X4 U67 ( .A0N(B[12]), .A1N(A[12]), .B0(n408), .Y(n378) );
  OAI2BB1X4 U68 ( .A0N(n450), .A1N(n336), .B0(B[25]), .Y(n337) );
  AOI211X2 U71 ( .A0(n306), .A1(n307), .B0(n305), .C0(n301), .Y(n401) );
  DLY1X1 U72 ( .A(n273), .Y(n331) );
  DLY1X1 U73 ( .A(n361), .Y(n332) );
  XNOR2X4 U76 ( .A(n342), .B(n431), .Y(SUM[21]) );
  DLY1X1 U77 ( .A(n349), .Y(n342) );
  NOR2BX4 U78 ( .AN(n373), .B(n410), .Y(n369) );
  INVXL U81 ( .A(n278), .Y(n351) );
  NOR2X1 U82 ( .A(n392), .B(n271), .Y(n400) );
  CLKBUFX2 U84 ( .A(n343), .Y(n338) );
  DLY1X1 U85 ( .A(n275), .Y(n335) );
  XOR2X1 U86 ( .A(n289), .B(n290), .Y(SUM[9]) );
  XOR2X4 U87 ( .A(n338), .B(n345), .Y(SUM[23]) );
  XNOR2X4 U90 ( .A(A[30]), .B(B[30]), .Y(n317) );
  INVX4 U91 ( .A(n422), .Y(SUM[26]) );
  NOR2X4 U93 ( .A(B[28]), .B(A[28]), .Y(n326) );
  INVX4 U95 ( .A(n356), .Y(n411) );
  NAND2BX4 U98 ( .AN(n336), .B(A[25]), .Y(n414) );
  INVX8 U99 ( .A(n320), .Y(n444) );
  INVX4 U102 ( .A(B[27]), .Y(n426) );
  NAND2X2 U103 ( .A(B[28]), .B(A[28]), .Y(n328) );
  INVXL U105 ( .A(n378), .Y(n360) );
  CLKINVX3 U106 ( .A(n360), .Y(n363) );
  OAI21X4 U107 ( .A0(n358), .A1(A[1]), .B0(B[1]), .Y(n404) );
  NAND2BXL U108 ( .AN(n305), .B(n307), .Y(n308) );
  DLY1X1 U109 ( .A(n369), .Y(n388) );
  DLY1X1 U110 ( .A(n364), .Y(n405) );
  XOR2XL U111 ( .A(n355), .B(n353), .Y(SUM[20]) );
  NAND2X4 U112 ( .A(n414), .B(n337), .Y(n406) );
  INVX8 U113 ( .A(B[7]), .Y(n441) );
  AOI21X1 U115 ( .A0(n399), .A1(n436), .B0(n392), .Y(n398) );
  AND2X2 U116 ( .A(B[10]), .B(A[10]), .Y(n392) );
  NAND2XL U117 ( .A(B[9]), .B(A[9]), .Y(n407) );
  NOR2X4 U118 ( .A(B[10]), .B(A[10]), .Y(n395) );
  NOR2X4 U119 ( .A(n411), .B(n412), .Y(n413) );
  OAI31X2 U120 ( .A0(n390), .A1(n391), .A2(n392), .B0(n393), .Y(n408) );
  OAI31X4 U121 ( .A0(n391), .A1(n392), .A2(n335), .B0(n393), .Y(n389) );
  AND2X4 U122 ( .A(n438), .B(n445), .Y(n410) );
  INVX8 U123 ( .A(B[15]), .Y(n438) );
  NOR2X4 U125 ( .A(n428), .B(n413), .Y(n353) );
  NAND2X4 U130 ( .A(n414), .B(n337), .Y(n333) );
  AND2X4 U133 ( .A(n330), .B(A[27]), .Y(n415) );
  NOR2X4 U135 ( .A(n425), .B(n415), .Y(n327) );
  XOR2X2 U136 ( .A(B[29]), .B(A[29]), .Y(n325) );
  NAND2X2 U137 ( .A(n447), .B(n441), .Y(n303) );
  AOI21X2 U141 ( .A0(n445), .A1(n438), .B0(n370), .Y(n380) );
  BUFX8 U146 ( .A(n452), .Y(SUM[24]) );
  OAI2BB1X4 U147 ( .A0N(A[29]), .A1N(n318), .B0(n319), .Y(n316) );
  AOI2BB2X4 U148 ( .B0(n315), .B1(n440), .A0N(n316), .A1N(A[30]), .Y(n313) );
  INVX4 U150 ( .A(n341), .Y(n439) );
  INVX4 U151 ( .A(n386), .Y(n437) );
  NOR2X4 U152 ( .A(A[12]), .B(B[12]), .Y(n386) );
  XOR2X1 U153 ( .A(n299), .B(n419), .Y(SUM[6]) );
  XOR2X1 U154 ( .A(B[22]), .B(A[22]), .Y(n348) );
  INVX3 U155 ( .A(B[19]), .Y(n429) );
  OAI2BB1X4 U156 ( .A0N(A[4]), .A1N(n310), .B0(n402), .Y(n434) );
  XOR2XL U157 ( .A(n433), .B(n336), .Y(n432) );
  XNOR2X1 U158 ( .A(n339), .B(n418), .Y(n452) );
  OR2XL U159 ( .A(n341), .B(n340), .Y(n418) );
  NAND2BXL U160 ( .AN(n391), .B(n393), .Y(n397) );
  NOR2XL U161 ( .A(n300), .B(n301), .Y(n419) );
  XOR2X1 U162 ( .A(n332), .B(n420), .Y(SUM[18]) );
  XOR2X1 U163 ( .A(n282), .B(A[18]), .Y(n420) );
  AOI21X4 U164 ( .A0(n333), .A1(A[26]), .B0(B[26]), .Y(n334) );
  NAND2X4 U165 ( .A(A[16]), .B(B[16]), .Y(n368) );
  XOR2X4 U166 ( .A(B[31]), .B(A[31]), .Y(n314) );
  NAND2XL U167 ( .A(n295), .B(n296), .Y(n294) );
  OAI21XL U168 ( .A0(n290), .A1(n270), .B0(n407), .Y(n399) );
  OR2X4 U169 ( .A(A[11]), .B(B[11]), .Y(n393) );
  NAND2BXL U170 ( .AN(n291), .B(n407), .Y(n289) );
  NAND2BXL U171 ( .AN(n377), .B(n375), .Y(n382) );
  NOR2BX4 U172 ( .AN(B[11]), .B(n446), .Y(n391) );
  OAI21XL U173 ( .A0(n305), .A1(n306), .B0(n307), .Y(n299) );
  XOR2X2 U174 ( .A(n399), .B(n400), .Y(SUM[10]) );
  XOR2X1 U175 ( .A(n308), .B(n306), .Y(SUM[5]) );
  AOI21XL U176 ( .A0(n443), .A1(n299), .B0(n300), .Y(n298) );
  NAND2BXL U177 ( .AN(n302), .B(n303), .Y(n297) );
  INVXL U178 ( .A(n301), .Y(n443) );
  AOI21XL U179 ( .A0(n442), .A1(n449), .B0(n358), .Y(SUM[0]) );
  XOR2X1 U180 ( .A(B[23]), .B(A[23]), .Y(n345) );
  INVX1 U181 ( .A(A[25]), .Y(n450) );
  AOI2BB1X4 U182 ( .A0N(n330), .A1N(A[27]), .B0(n426), .Y(n425) );
  XNOR2X4 U183 ( .A(B[27]), .B(A[27]), .Y(n427) );
  XNOR2X1 U184 ( .A(n384), .B(n385), .Y(SUM[13]) );
  INVXL U185 ( .A(B[30]), .Y(n440) );
  AOI2BB1X4 U186 ( .A0N(n356), .A1N(A[19]), .B0(n429), .Y(n428) );
  XOR2XL U187 ( .A(A[19]), .B(B[19]), .Y(n430) );
  XNOR2X1 U188 ( .A(B[21]), .B(A[21]), .Y(n431) );
  XOR2X1 U189 ( .A(A[25]), .B(B[25]), .Y(n433) );
  XOR2X1 U190 ( .A(B[17]), .B(A[17]), .Y(n366) );
  XOR2X2 U191 ( .A(n371), .B(n372), .Y(SUM[16]) );
  OAI21XL U192 ( .A0(A[16]), .A1(B[16]), .B0(n368), .Y(n371) );
  XOR2X1 U193 ( .A(n358), .B(n359), .Y(SUM[1]) );
  XOR2X1 U194 ( .A(n276), .B(n312), .Y(SUM[3]) );
  XNOR2XL U195 ( .A(A[3]), .B(B[3]), .Y(n312) );
  XNOR2XL U196 ( .A(n309), .B(n310), .Y(SUM[4]) );
  XNOR2XL U197 ( .A(A[4]), .B(B[4]), .Y(n309) );
  INVX1 U198 ( .A(A[7]), .Y(n447) );
  INVX1 U199 ( .A(A[11]), .Y(n446) );
  OAI21X4 U200 ( .A0(n318), .A1(A[29]), .B0(B[29]), .Y(n319) );
  XOR2X4 U201 ( .A(n318), .B(n325), .Y(SUM[29]) );
  BUFX4 U202 ( .A(n453), .Y(SUM[12]) );
  OAI21XL U203 ( .A0(n386), .A1(n363), .B0(n387), .Y(n453) );
  AND2X1 U204 ( .A(n363), .B(n437), .Y(n384) );
  NOR2XL U205 ( .A(n370), .B(n388), .Y(n372) );
  XOR2X1 U206 ( .A(n331), .B(n294), .Y(SUM[8]) );
  XOR2X1 U207 ( .A(B[1]), .B(A[1]), .Y(n359) );
  AND2X4 U208 ( .A(n292), .B(n295), .Y(n396) );
  AND2X1 U209 ( .A(n394), .B(n295), .Y(n290) );
  OAI33X2 U210 ( .A0(n394), .A1(n283), .A2(n291), .B0(n395), .B1(n396), .B2(
        n291), .Y(n390) );
  XOR2X1 U211 ( .A(n346), .B(n348), .Y(SUM[22]) );
  XOR2X1 U212 ( .A(n405), .B(n366), .Y(SUM[17]) );
  OAI21XL U213 ( .A0(n320), .A1(n321), .B0(n322), .Y(SUM[2]) );
  CLKINVX4 U214 ( .A(A[0]), .Y(n449) );
endmodule


module hash_core_DW01_add_26 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n276, n277, n278, n279, n280, n281, n282, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n299, n300,
         n301, n302, n303, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n317, n318, n320, n321, n323, n324, n326, n327,
         n329, n330, n331, n332, n333, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n369, n370, n371, n372, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n263, n264, n265, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n283, n297, n298, n304,
         n316, n319, n322, n325, n328, n334, n368, n373, n393, n394, n395,
         n396;

  OAI21X4 U8 ( .A0(n284), .A1(n285), .B0(n286), .Y(n282) );
  AND2X2 U10 ( .A(n288), .B(n289), .Y(n285) );
  XOR2X4 U21 ( .A(n302), .B(n303), .Y(SUM[31]) );
  XOR2X4 U25 ( .A(n305), .B(n306), .Y(SUM[30]) );
  OAI21X4 U33 ( .A0(A[28]), .A1(n314), .B0(B[28]), .Y(n315) );
  OAI2BB1X4 U36 ( .A0N(n317), .A1N(A[27]), .B0(n318), .Y(n314) );
  OAI21X4 U37 ( .A0(A[27]), .A1(n317), .B0(B[27]), .Y(n318) );
  OAI2BB1X4 U40 ( .A0N(n320), .A1N(A[26]), .B0(n321), .Y(n317) );
  OAI21X4 U41 ( .A0(A[26]), .A1(n320), .B0(B[26]), .Y(n321) );
  OAI2BB1X4 U44 ( .A0N(n323), .A1N(A[25]), .B0(n324), .Y(n320) );
  OAI21X4 U45 ( .A0(A[25]), .A1(n323), .B0(B[25]), .Y(n324) );
  OAI2BB1X4 U48 ( .A0N(n326), .A1N(A[24]), .B0(n327), .Y(n323) );
  OAI21X4 U49 ( .A0(A[24]), .A1(n326), .B0(B[24]), .Y(n327) );
  OAI2BB1X4 U52 ( .A0N(n329), .A1N(A[23]), .B0(n330), .Y(n326) );
  OAI21X4 U53 ( .A0(A[23]), .A1(n329), .B0(B[23]), .Y(n330) );
  OAI2BB1X4 U56 ( .A0N(n332), .A1N(A[22]), .B0(n333), .Y(n329) );
  OAI21X4 U57 ( .A0(A[22]), .A1(n332), .B0(B[22]), .Y(n333) );
  OAI2BB1X4 U60 ( .A0N(n335), .A1N(A[21]), .B0(n336), .Y(n332) );
  OAI21X4 U61 ( .A0(A[21]), .A1(n335), .B0(B[21]), .Y(n336) );
  OAI2BB1X4 U64 ( .A0N(n338), .A1N(A[20]), .B0(n339), .Y(n335) );
  OAI21X4 U65 ( .A0(A[20]), .A1(n338), .B0(B[20]), .Y(n339) );
  OAI2BB1X4 U68 ( .A0N(n341), .A1N(A[19]), .B0(n342), .Y(n338) );
  OAI21X4 U69 ( .A0(A[19]), .A1(n341), .B0(B[19]), .Y(n342) );
  OAI2BB1X4 U74 ( .A0N(n346), .A1N(A[18]), .B0(n347), .Y(n341) );
  OAI21X4 U75 ( .A0(A[18]), .A1(n346), .B0(B[18]), .Y(n347) );
  OAI2BB1X4 U78 ( .A0N(n349), .A1N(A[17]), .B0(n350), .Y(n346) );
  OAI21X4 U79 ( .A0(A[17]), .A1(n349), .B0(B[17]), .Y(n350) );
  OAI2BB1X4 U82 ( .A0N(n352), .A1N(A[16]), .B0(n353), .Y(n349) );
  OAI21X4 U83 ( .A0(n352), .A1(A[16]), .B0(B[16]), .Y(n353) );
  AOI2BB1X4 U87 ( .A0N(A[15]), .A1N(n355), .B0(n356), .Y(n352) );
  AOI21X4 U88 ( .A0(n355), .A1(A[15]), .B0(B[15]), .Y(n356) );
  OAI21X4 U89 ( .A0(n357), .A1(n358), .B0(n359), .Y(n355) );
  AOI31X2 U90 ( .A0(n395), .A1(n394), .A2(n360), .B0(n393), .Y(n358) );
  XOR2X4 U91 ( .A(n362), .B(n363), .Y(SUM[15]) );
  XOR2X4 U94 ( .A(n364), .B(n365), .Y(SUM[14]) );
  OAI21X4 U98 ( .A0(n366), .A1(n367), .B0(n361), .Y(n364) );
  NAND4BX4 U109 ( .AN(n280), .B(n368), .C(n319), .D(n376), .Y(n375) );
  AOI211X2 U112 ( .A0(n278), .A1(n281), .B0(n379), .C0(n380), .Y(n378) );
  AND2X2 U117 ( .A(B[11]), .B(A[11]), .Y(n377) );
  NAND2X4 U123 ( .A(B[8]), .B(A[8]), .Y(n281) );
  NOR3X4 U125 ( .A(n387), .B(n388), .C(n389), .Y(n280) );
  NAND2BX4 U127 ( .AN(n296), .B(n294), .Y(n292) );
  NAND2X4 U128 ( .A(n301), .B(n391), .Y(n294) );
  OAI21X4 U129 ( .A0(n299), .A1(n328), .B0(n300), .Y(n391) );
  OR2X4 U130 ( .A(A[3]), .B(B[3]), .Y(n300) );
  AND2X2 U132 ( .A(n310), .B(n312), .Y(n299) );
  OR2X4 U133 ( .A(B[2]), .B(A[2]), .Y(n312) );
  OAI2BB1X4 U134 ( .A0N(n343), .A1N(A[1]), .B0(n392), .Y(n310) );
  OAI21X4 U135 ( .A0(n343), .A1(A[1]), .B0(B[1]), .Y(n392) );
  NAND2X4 U139 ( .A(B[6]), .B(A[6]), .Y(n286) );
  NOR2X4 U141 ( .A(A[6]), .B(B[6]), .Y(n284) );
  OAI22X4 U142 ( .A0(B[7]), .A1(A[7]), .B0(B[5]), .B1(A[5]), .Y(n390) );
  NOR2X4 U145 ( .A(A[9]), .B(B[9]), .Y(n380) );
  NOR2X4 U147 ( .A(A[10]), .B(B[10]), .Y(n379) );
  NAND2X4 U148 ( .A(B[10]), .B(A[10]), .Y(n384) );
  NOR2X4 U150 ( .A(n396), .B(n304), .Y(n343) );
  INVX4 U2 ( .A(n380), .Y(n368) );
  XNOR2X2 U3 ( .A(n313), .B(n307), .Y(SUM[29]) );
  NOR2X2 U4 ( .A(A[13]), .B(B[13]), .Y(n366) );
  NOR2X2 U5 ( .A(A[12]), .B(B[12]), .Y(n369) );
  AOI211XL U6 ( .A0(n293), .A1(n289), .B0(n390), .C0(n284), .Y(n387) );
  INVX1 U7 ( .A(B[30]), .Y(n274) );
  XOR2X2 U9 ( .A(n381), .B(n382), .Y(SUM[11]) );
  XNOR2X1 U11 ( .A(n385), .B(n383), .Y(SUM[10]) );
  OAI21XL U12 ( .A0(A[5]), .A1(B[5]), .B0(n290), .Y(n288) );
  CLKINVX8 U13 ( .A(B[0]), .Y(n396) );
  AOI21X4 U14 ( .A0(n307), .A1(A[29]), .B0(B[29]), .Y(n308) );
  OAI2BB1X2 U15 ( .A0N(n314), .A1N(A[28]), .B0(n315), .Y(n307) );
  AOI2BB1X4 U16 ( .A0N(A[29]), .A1N(n307), .B0(n308), .Y(n305) );
  XNOR2X4 U17 ( .A(n345), .B(n341), .Y(SUM[19]) );
  NAND2XL U18 ( .A(B[13]), .B(A[13]), .Y(n361) );
  NAND2XL U19 ( .A(B[12]), .B(A[12]), .Y(n371) );
  XNOR2X2 U20 ( .A(n367), .B(n263), .Y(SUM[13]) );
  XNOR2X1 U22 ( .A(n265), .B(n314), .Y(SUM[28]) );
  NAND2X4 U23 ( .A(B[9]), .B(A[9]), .Y(n278) );
  XOR2X2 U24 ( .A(n283), .B(n323), .Y(SUM[25]) );
  INVXL U26 ( .A(n374), .Y(n268) );
  NAND2XL U27 ( .A(n292), .B(n293), .Y(n290) );
  XNOR2X1 U28 ( .A(n331), .B(n329), .Y(SUM[23]) );
  XNOR2X1 U29 ( .A(n264), .B(n320), .Y(SUM[26]) );
  CLKINVX2 U30 ( .A(A[7]), .Y(n334) );
  NAND2X2 U31 ( .A(B[5]), .B(A[5]), .Y(n289) );
  NAND2XL U32 ( .A(n360), .B(n395), .Y(n367) );
  NAND2BX4 U34 ( .AN(n372), .B(n371), .Y(n360) );
  OAI32X2 U35 ( .A0(n292), .A1(n284), .A2(n390), .B0(n286), .B1(n334), .Y(n389) );
  AOI21X2 U38 ( .A0(n334), .A1(n286), .B0(n373), .Y(n388) );
  XOR2X4 U39 ( .A(n287), .B(n285), .Y(SUM[6]) );
  AND2X1 U42 ( .A(n361), .B(n394), .Y(n263) );
  AOI21XL U43 ( .A0(n383), .A1(n319), .B0(n316), .Y(n382) );
  NOR2XL U46 ( .A(n322), .B(n357), .Y(n365) );
  XNOR2X1 U47 ( .A(A[26]), .B(B[26]), .Y(n264) );
  OAI21X4 U50 ( .A0(n280), .A1(n386), .B0(n281), .Y(n277) );
  NOR2XL U51 ( .A(A[8]), .B(B[8]), .Y(n386) );
  NOR2X2 U54 ( .A(B[4]), .B(A[4]), .Y(n296) );
  XNOR2X1 U55 ( .A(A[28]), .B(B[28]), .Y(n265) );
  NAND2X2 U58 ( .A(B[2]), .B(A[2]), .Y(n311) );
  INVX12 U59 ( .A(n272), .Y(SUM[24]) );
  NAND2X1 U62 ( .A(B[3]), .B(A[3]), .Y(n301) );
  XNOR2XL U63 ( .A(n267), .B(n332), .Y(SUM[22]) );
  XNOR2X1 U66 ( .A(A[22]), .B(B[22]), .Y(n267) );
  AOI2BB1X1 U67 ( .A0N(A[8]), .A1N(B[8]), .B0(n374), .Y(n376) );
  NOR2X4 U70 ( .A(A[11]), .B(B[11]), .Y(n374) );
  INVXL U71 ( .A(n357), .Y(n325) );
  AOI21X4 U72 ( .A0(n325), .A1(n364), .B0(n322), .Y(n363) );
  NAND2XL U73 ( .A(B[14]), .B(A[14]), .Y(n359) );
  OAI2BB1X4 U76 ( .A0N(n269), .A1N(n268), .B0(n375), .Y(n372) );
  OR3X4 U77 ( .A(n377), .B(n378), .C(n316), .Y(n269) );
  OAI2BB1X1 U80 ( .A0N(n368), .A1N(n277), .B0(n278), .Y(n383) );
  NAND2BXL U81 ( .AN(n284), .B(n286), .Y(n287) );
  XOR2X2 U84 ( .A(n270), .B(n271), .Y(SUM[3]) );
  AND2X1 U85 ( .A(n300), .B(n301), .Y(n270) );
  OR2XL U86 ( .A(n328), .B(n299), .Y(n271) );
  NAND2XL U92 ( .A(n384), .B(n319), .Y(n385) );
  INVX1 U93 ( .A(n311), .Y(n328) );
  OAI21XL U95 ( .A0(n369), .A1(n360), .B0(n370), .Y(SUM[12]) );
  OAI2BB1XL U96 ( .A0N(n395), .A1N(n371), .B0(n372), .Y(n370) );
  XNOR2X1 U97 ( .A(n276), .B(n277), .Y(SUM[9]) );
  NAND2X1 U99 ( .A(n368), .B(n278), .Y(n276) );
  XNOR2XL U100 ( .A(n309), .B(n310), .Y(SUM[2]) );
  NAND2XL U101 ( .A(n311), .B(n312), .Y(n309) );
  XOR2X1 U102 ( .A(n294), .B(n295), .Y(SUM[4]) );
  NOR2BX1 U103 ( .AN(n293), .B(n296), .Y(n295) );
  OR2XL U104 ( .A(n374), .B(n377), .Y(n381) );
  INVX1 U105 ( .A(B[7]), .Y(n373) );
  INVX1 U106 ( .A(n369), .Y(n395) );
  INVX1 U107 ( .A(n366), .Y(n394) );
  INVX1 U108 ( .A(n361), .Y(n393) );
  INVX1 U110 ( .A(n359), .Y(n322) );
  XNOR2XL U111 ( .A(n273), .B(n326), .Y(n272) );
  XOR2X1 U113 ( .A(A[24]), .B(B[24]), .Y(n273) );
  AOI2BB2X2 U114 ( .B0(A[30]), .B1(n305), .A0N(n274), .A1N(n275), .Y(n303) );
  NOR2X2 U115 ( .A(A[30]), .B(n305), .Y(n275) );
  XOR2X1 U116 ( .A(B[30]), .B(A[30]), .Y(n306) );
  XOR2X1 U118 ( .A(A[25]), .B(B[25]), .Y(n283) );
  XNOR2X1 U119 ( .A(A[23]), .B(B[23]), .Y(n331) );
  XNOR2X1 U120 ( .A(A[29]), .B(B[29]), .Y(n313) );
  XNOR2X4 U121 ( .A(n282), .B(n297), .Y(SUM[7]) );
  XOR2XL U122 ( .A(n373), .B(A[7]), .Y(n297) );
  XOR2X1 U124 ( .A(n298), .B(n317), .Y(SUM[27]) );
  XOR2X1 U126 ( .A(A[27]), .B(B[27]), .Y(n298) );
  AOI21XL U131 ( .A0(n396), .A1(n304), .B0(n343), .Y(SUM[0]) );
  XNOR2XL U136 ( .A(n340), .B(n338), .Y(SUM[20]) );
  XNOR2X1 U137 ( .A(A[20]), .B(B[20]), .Y(n340) );
  XNOR2X1 U138 ( .A(A[19]), .B(B[19]), .Y(n345) );
  XNOR2XL U140 ( .A(n348), .B(n346), .Y(SUM[18]) );
  XNOR2X1 U143 ( .A(A[18]), .B(B[18]), .Y(n348) );
  XNOR2XL U144 ( .A(n337), .B(n335), .Y(SUM[21]) );
  XNOR2X1 U146 ( .A(A[21]), .B(B[21]), .Y(n337) );
  XOR2XL U149 ( .A(n279), .B(n280), .Y(SUM[8]) );
  OAI21XL U151 ( .A0(B[8]), .A1(A[8]), .B0(n281), .Y(n279) );
  XNOR2X1 U152 ( .A(A[15]), .B(B[15]), .Y(n362) );
  NAND2X1 U153 ( .A(B[4]), .B(A[4]), .Y(n293) );
  XOR2X1 U154 ( .A(n352), .B(n354), .Y(SUM[16]) );
  XOR2X1 U155 ( .A(B[16]), .B(A[16]), .Y(n354) );
  XNOR2X1 U156 ( .A(n290), .B(n291), .Y(SUM[5]) );
  OAI21XL U157 ( .A0(A[5]), .A1(B[5]), .B0(n289), .Y(n291) );
  XNOR2XL U158 ( .A(n351), .B(n349), .Y(SUM[17]) );
  XNOR2X1 U159 ( .A(A[17]), .B(B[17]), .Y(n351) );
  XOR2X1 U160 ( .A(n343), .B(n344), .Y(SUM[1]) );
  XOR2X1 U161 ( .A(B[1]), .B(A[1]), .Y(n344) );
  NOR2X1 U162 ( .A(B[14]), .B(A[14]), .Y(n357) );
  XNOR2X1 U163 ( .A(B[31]), .B(A[31]), .Y(n302) );
  CLKINVX4 U164 ( .A(A[0]), .Y(n304) );
  CLKINVX4 U165 ( .A(n384), .Y(n316) );
  CLKINVX4 U166 ( .A(n379), .Y(n319) );
endmodule


module hash_core_DW01_add_27 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n587, n588, n589, n590, n591, n414, n416, n417, n419, n420, n421,
         n422, n423, n424, n425, n426, n428, n429, n430, n431, n432, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n452, n453, n455, n456, n458, n459, n460, n461, n462,
         n465, n466, n468, n469, n470, n471, n472, n473, n475, n477, n478,
         n479, n480, n481, n482, n483, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n528, n529, n530, n531, n532, n533, n396, n397, n398, n399,
         n400, n401, n402, n404, n405, n407, n408, n409, n410, n411, n412,
         n413, n415, n418, n427, n433, n434, n435, n450, n451, n454, n457,
         n463, n464, n467, n474, n476, n484, n485, n496, n527, n534, n535,
         n537, n539, n540, n541, n542, n544, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586;

  XOR2X4 U20 ( .A(n437), .B(n438), .Y(SUM[31]) );
  XOR2X4 U21 ( .A(B[31]), .B(A[31]), .Y(n438) );
  NOR2BX4 U24 ( .AN(n441), .B(n439), .Y(n442) );
  NAND2X4 U26 ( .A(B[30]), .B(A[30]), .Y(n441) );
  OAI21X4 U40 ( .A0(n455), .A1(n401), .B0(B[27]), .Y(n456) );
  OAI21X4 U43 ( .A0(n459), .A1(n458), .B0(n460), .Y(n455) );
  NAND2BX4 U47 ( .AN(n458), .B(n460), .Y(n461) );
  NOR2X4 U49 ( .A(B[26]), .B(A[26]), .Y(n458) );
  OAI2BB1X4 U52 ( .A0N(n402), .A1N(n465), .B0(n466), .Y(n462) );
  OAI21X4 U53 ( .A0(n465), .A1(n402), .B0(B[24]), .Y(n466) );
  OAI2BB1X4 U56 ( .A0N(A[23]), .A1N(n468), .B0(n469), .Y(n465) );
  OAI21X4 U57 ( .A0(n468), .A1(A[23]), .B0(B[23]), .Y(n469) );
  OAI21X4 U60 ( .A0(n472), .A1(n471), .B0(n473), .Y(n468) );
  OAI2BB1X4 U68 ( .A0N(A[20]), .A1N(n478), .B0(n479), .Y(n475) );
  OAI21X4 U69 ( .A0(n478), .A1(A[20]), .B0(B[20]), .Y(n479) );
  XNOR2X4 U70 ( .A(A[21]), .B(B[21]), .Y(n477) );
  OAI2BB1X4 U72 ( .A0N(A[19]), .A1N(n481), .B0(n482), .Y(n478) );
  OAI21X4 U73 ( .A0(n481), .A1(A[19]), .B0(B[19]), .Y(n482) );
  XNOR2X4 U74 ( .A(A[20]), .B(B[20]), .Y(n480) );
  OAI21X4 U78 ( .A0(n464), .A1(n486), .B0(n488), .Y(n481) );
  NOR2X4 U82 ( .A(n400), .B(A[18]), .Y(n486) );
  XOR2X4 U87 ( .A(n494), .B(n495), .Y(SUM[17]) );
  XOR2X4 U91 ( .A(n396), .B(n497), .Y(SUM[16]) );
  NOR2X4 U93 ( .A(n579), .B(n582), .Y(n490) );
  OAI31X2 U94 ( .A0(n498), .A1(n499), .A2(n500), .B0(n501), .Y(n492) );
  AOI211X2 U96 ( .A0(n504), .A1(n505), .B0(n506), .C0(n507), .Y(n503) );
  XOR2X4 U97 ( .A(n509), .B(n510), .Y(SUM[15]) );
  NOR2X4 U99 ( .A(B[15]), .B(A[15]), .Y(n500) );
  XOR2X4 U102 ( .A(n407), .B(n512), .Y(SUM[14]) );
  NAND2BX4 U104 ( .AN(n499), .B(n508), .Y(n512) );
  NAND2X4 U105 ( .A(B[14]), .B(A[14]), .Y(n508) );
  XOR2X4 U107 ( .A(n513), .B(n514), .Y(n589) );
  NOR2X4 U110 ( .A(A[13]), .B(B[13]), .Y(n506) );
  AOI2BB1X4 U113 ( .A0N(n516), .A1N(n517), .B0(n518), .Y(n504) );
  AOI211X2 U116 ( .A0(n525), .A1(n524), .B0(n520), .C0(n416), .Y(n522) );
  NOR2X4 U122 ( .A(A[11]), .B(B[11]), .Y(n517) );
  AOI2BB1X4 U126 ( .A0N(n414), .A1N(n467), .B0(n576), .Y(n528) );
  NAND2X4 U127 ( .A(B[9]), .B(A[9]), .Y(n525) );
  NOR2X4 U128 ( .A(B[9]), .B(A[9]), .Y(n416) );
  NOR2X4 U129 ( .A(n519), .B(n580), .Y(n414) );
  NAND2X4 U130 ( .A(B[8]), .B(A[8]), .Y(n524) );
  NOR2BX4 U131 ( .AN(n417), .B(n419), .Y(n519) );
  NOR2X4 U132 ( .A(B[8]), .B(A[8]), .Y(n419) );
  AOI31X2 U133 ( .A0(n422), .A1(n426), .A2(n530), .B0(n423), .Y(n417) );
  NOR2X4 U134 ( .A(B[7]), .B(A[7]), .Y(n423) );
  NAND2X4 U135 ( .A(B[7]), .B(A[7]), .Y(n422) );
  OAI221X2 U137 ( .A0(n428), .A1(n485), .B0(A[5]), .B1(n476), .C0(n584), .Y(
        n530) );
  NOR2X4 U138 ( .A(B[6]), .B(A[6]), .Y(n424) );
  OAI2BB1X4 U140 ( .A0N(A[4]), .A1N(n432), .B0(n531), .Y(n428) );
  OAI21X4 U141 ( .A0(n432), .A1(A[4]), .B0(B[4]), .Y(n531) );
  OAI2BB1X4 U142 ( .A0N(A[3]), .A1N(n451), .B0(n532), .Y(n432) );
  OAI2BB1X4 U147 ( .A0N(n537), .A1N(A[1]), .B0(n533), .Y(n449) );
  NOR2X4 U151 ( .A(B[10]), .B(A[10]), .Y(n520) );
  NOR2X4 U153 ( .A(n585), .B(n581), .Y(n483) );
  CLKBUFX8 U2 ( .A(B[2]), .Y(n484) );
  NAND2BX2 U3 ( .AN(n520), .B(n523), .Y(n529) );
  CLKINVX4 U4 ( .A(n548), .Y(n396) );
  INVX4 U5 ( .A(n572), .Y(n548) );
  OAI31X2 U6 ( .A0(n498), .A1(n499), .A2(n500), .B0(n501), .Y(n572) );
  NOR3BX4 U7 ( .AN(n508), .B(n503), .C(n502), .Y(n498) );
  BUFX20 U8 ( .A(n590), .Y(SUM[10]) );
  BUFX16 U9 ( .A(n591), .Y(SUM[9]) );
  OAI21X4 U10 ( .A0(n463), .A1(n527), .B0(n523), .Y(n526) );
  NOR2X2 U11 ( .A(n564), .B(n534), .Y(n397) );
  BUFX8 U12 ( .A(n520), .Y(n527) );
  BUFX8 U13 ( .A(A[27]), .Y(n398) );
  NAND2X4 U14 ( .A(B[10]), .B(A[10]), .Y(n523) );
  NAND4BBX4 U15 ( .AN(n412), .BN(n517), .C(n399), .D(n413), .Y(n415) );
  AND2X4 U16 ( .A(n475), .B(A[21]), .Y(n534) );
  BUFX16 U17 ( .A(n587), .Y(SUM[29]) );
  BUFX8 U18 ( .A(n546), .Y(SUM[4]) );
  INVX4 U19 ( .A(n450), .Y(n451) );
  CLKINVX4 U22 ( .A(n443), .Y(n573) );
  XOR2X2 U23 ( .A(n451), .B(A[3]), .Y(n554) );
  DLY1X1 U25 ( .A(n428), .Y(n496) );
  INVX1 U27 ( .A(n506), .Y(n577) );
  INVX4 U28 ( .A(n415), .Y(n518) );
  INVX4 U29 ( .A(A[5]), .Y(n583) );
  INVX4 U30 ( .A(n424), .Y(n584) );
  AND2X2 U31 ( .A(n462), .B(A[25]), .Y(n535) );
  NAND2X1 U32 ( .A(B[22]), .B(A[22]), .Y(n473) );
  NOR2X2 U33 ( .A(B[22]), .B(A[22]), .Y(n471) );
  CLKINVX3 U34 ( .A(n409), .Y(SUM[20]) );
  BUFX16 U35 ( .A(n483), .Y(n537) );
  INVX3 U36 ( .A(B[3]), .Y(n450) );
  INVX1 U37 ( .A(n416), .Y(n413) );
  BUFX8 U38 ( .A(n416), .Y(n467) );
  INVXL U39 ( .A(n519), .Y(n412) );
  INVX2 U41 ( .A(B[29]), .Y(n405) );
  INVX4 U42 ( .A(n527), .Y(n399) );
  INVX8 U44 ( .A(n568), .Y(SUM[27]) );
  XOR2X4 U45 ( .A(n455), .B(n569), .Y(n568) );
  OAI21X1 U46 ( .A0(n439), .A1(n440), .B0(n441), .Y(n437) );
  AOI21X2 U48 ( .A0(n513), .A1(n577), .B0(n502), .Y(n511) );
  XOR2X1 U50 ( .A(n478), .B(n480), .Y(n409) );
  INVX3 U51 ( .A(n523), .Y(n575) );
  AND2X4 U54 ( .A(n408), .B(n426), .Y(n551) );
  BUFX8 U55 ( .A(B[18]), .Y(n400) );
  BUFX8 U58 ( .A(n398), .Y(n401) );
  BUFX8 U59 ( .A(A[24]), .Y(n402) );
  XNOR2X4 U61 ( .A(n487), .B(n489), .Y(SUM[18]) );
  NAND2BX4 U62 ( .AN(n504), .B(n404), .Y(n542) );
  CLKINVX20 U63 ( .A(n507), .Y(n404) );
  INVX4 U64 ( .A(n421), .Y(n454) );
  XOR2X4 U65 ( .A(A[29]), .B(n405), .Y(n567) );
  INVX8 U66 ( .A(B[0]), .Y(n585) );
  NAND2X2 U67 ( .A(n583), .B(n586), .Y(n429) );
  AND2X4 U71 ( .A(B[5]), .B(A[5]), .Y(n485) );
  BUFX12 U75 ( .A(n589), .Y(SUM[13]) );
  AND2X4 U76 ( .A(B[13]), .B(A[13]), .Y(n502) );
  AOI21X4 U77 ( .A0(n577), .A1(n513), .B0(n502), .Y(n407) );
  NOR2X4 U79 ( .A(A[2]), .B(n484), .Y(n446) );
  XOR2X4 U80 ( .A(n414), .B(n552), .Y(n591) );
  NOR2BX4 U81 ( .AN(n501), .B(n500), .Y(n510) );
  NAND2X4 U83 ( .A(B[15]), .B(A[15]), .Y(n501) );
  CLKINVX3 U84 ( .A(n584), .Y(n427) );
  OR2X2 U85 ( .A(n448), .B(n449), .Y(n436) );
  AOI21X2 U86 ( .A0(n585), .A1(n581), .B0(n537), .Y(SUM[0]) );
  INVX8 U88 ( .A(A[0]), .Y(n581) );
  INVX2 U89 ( .A(n427), .Y(n408) );
  INVX2 U90 ( .A(A[2]), .Y(n433) );
  NOR3X2 U92 ( .A(n522), .B(n521), .C(n575), .Y(n516) );
  INVX8 U95 ( .A(n411), .Y(n444) );
  INVX12 U98 ( .A(n557), .Y(SUM[19]) );
  INVX4 U100 ( .A(A[29]), .Y(n474) );
  XNOR2XL U101 ( .A(n558), .B(n481), .Y(n557) );
  INVX2 U103 ( .A(n586), .Y(n476) );
  OAI21X2 U106 ( .A0(n446), .A1(n448), .B0(n449), .Y(n447) );
  OR2X4 U108 ( .A(n419), .B(n580), .Y(n540) );
  INVX4 U109 ( .A(n524), .Y(n580) );
  NAND2X4 U111 ( .A(n452), .B(n410), .Y(n411) );
  INVX4 U112 ( .A(n453), .Y(n410) );
  OAI21X4 U114 ( .A0(n436), .A1(n446), .B0(n447), .Y(SUM[2]) );
  XNOR3X4 U115 ( .A(A[22]), .B(B[22]), .C(n397), .Y(SUM[22]) );
  XNOR2X4 U117 ( .A(n459), .B(n461), .Y(n418) );
  INVX8 U118 ( .A(n418), .Y(SUM[26]) );
  OAI2BB1X4 U119 ( .A0N(n401), .A1N(n455), .B0(n456), .Y(n452) );
  OAI221X2 U120 ( .A0(B[3]), .A1(A[3]), .B0(n448), .B1(n449), .C0(n457), .Y(
        n532) );
  OAI21X2 U121 ( .A0(n490), .A1(A[17]), .B0(B[17]), .Y(n493) );
  NOR2X1 U123 ( .A(n586), .B(n583), .Y(n430) );
  NAND2BX4 U124 ( .AN(n484), .B(n433), .Y(n457) );
  XOR2X2 U125 ( .A(n468), .B(n470), .Y(n588) );
  INVX8 U136 ( .A(A[16]), .Y(n582) );
  INVX4 U139 ( .A(n493), .Y(n578) );
  INVXL U143 ( .A(n432), .Y(n434) );
  INVX2 U144 ( .A(n434), .Y(n435) );
  AOI211X2 U145 ( .A0(A[29]), .A1(B[29]), .B0(n444), .C0(n445), .Y(n443) );
  XOR2X2 U146 ( .A(B[1]), .B(A[1]), .Y(n550) );
  XOR2X1 U148 ( .A(A[19]), .B(B[19]), .Y(n558) );
  NOR2X2 U149 ( .A(n506), .B(n502), .Y(n514) );
  XNOR2X4 U150 ( .A(n420), .B(n454), .Y(SUM[7]) );
  AOI2BB1X4 U152 ( .A0N(n549), .A1N(n548), .B0(n490), .Y(n495) );
  AOI211X4 U154 ( .A0(n490), .A1(A[17]), .B0(n578), .C0(n574), .Y(n487) );
  AOI21X2 U155 ( .A0(n583), .A1(n586), .B0(n430), .Y(n431) );
  XOR2X4 U156 ( .A(n496), .B(n431), .Y(SUM[5]) );
  NAND2X4 U157 ( .A(n400), .B(A[18]), .Y(n488) );
  AOI2BB1X2 U158 ( .A0N(n414), .A1N(n467), .B0(n576), .Y(n463) );
  AOI211X2 U159 ( .A0(n490), .A1(A[17]), .B0(n574), .C0(n578), .Y(n464) );
  OAI2BB1X4 U160 ( .A0N(n405), .A1N(n474), .B0(n573), .Y(n440) );
  OR2X1 U161 ( .A(n521), .B(n517), .Y(n555) );
  INVX8 U162 ( .A(n525), .Y(n576) );
  NOR2BX4 U163 ( .AN(n422), .B(n423), .Y(n421) );
  XNOR2X2 U164 ( .A(n504), .B(n515), .Y(n541) );
  INVX8 U165 ( .A(n541), .Y(SUM[12]) );
  XNOR2X1 U166 ( .A(B[17]), .B(A[17]), .Y(n494) );
  INVX4 U167 ( .A(n491), .Y(n574) );
  OAI21X4 U168 ( .A0(n511), .A1(n499), .B0(n508), .Y(n509) );
  NOR2X4 U169 ( .A(n564), .B(n534), .Y(n472) );
  NOR2X4 U170 ( .A(n562), .B(n535), .Y(n459) );
  AND2X1 U171 ( .A(n457), .B(n436), .Y(n553) );
  BUFX12 U172 ( .A(n588), .Y(SUM[23]) );
  XNOR2X2 U173 ( .A(B[27]), .B(A[27]), .Y(n569) );
  XOR2X2 U174 ( .A(B[23]), .B(A[23]), .Y(n470) );
  AOI21X2 U175 ( .A0(n582), .A1(n579), .B0(n490), .Y(n497) );
  INVX8 U176 ( .A(B[16]), .Y(n579) );
  AOI21X2 U177 ( .A0(n429), .A1(n428), .B0(n485), .Y(n425) );
  OR2X4 U178 ( .A(n576), .B(n416), .Y(n552) );
  OAI21X4 U179 ( .A0(n537), .A1(A[1]), .B0(B[1]), .Y(n533) );
  OAI221X2 U180 ( .A0(B[16]), .A1(A[16]), .B0(A[17]), .B1(B[17]), .C0(n492), 
        .Y(n491) );
  INVXL U181 ( .A(n417), .Y(n539) );
  XOR2X4 U182 ( .A(n539), .B(n540), .Y(SUM[8]) );
  OAI21X2 U183 ( .A0(n425), .A1(n427), .B0(n426), .Y(n420) );
  NOR2BX4 U184 ( .AN(n488), .B(n486), .Y(n489) );
  NAND2X4 U185 ( .A(B[26]), .B(A[26]), .Y(n460) );
  XOR2X4 U186 ( .A(n452), .B(n544), .Y(SUM[28]) );
  INVX8 U187 ( .A(n560), .Y(SUM[24]) );
  NOR2X4 U188 ( .A(n444), .B(n445), .Y(n566) );
  NAND2X4 U189 ( .A(n542), .B(n505), .Y(n513) );
  NAND2X4 U190 ( .A(B[12]), .B(A[12]), .Y(n505) );
  NOR2X4 U191 ( .A(B[12]), .B(A[12]), .Y(n507) );
  NOR2X4 U192 ( .A(A[14]), .B(B[14]), .Y(n499) );
  NOR2X4 U193 ( .A(n453), .B(n445), .Y(n544) );
  XOR2X1 U194 ( .A(n435), .B(n547), .Y(n546) );
  XOR2X1 U195 ( .A(B[4]), .B(A[4]), .Y(n547) );
  INVXL U196 ( .A(B[25]), .Y(n563) );
  INVX2 U197 ( .A(B[21]), .Y(n565) );
  AND2X1 U198 ( .A(n579), .B(n582), .Y(n549) );
  NOR2X4 U199 ( .A(B[30]), .B(A[30]), .Y(n439) );
  XOR2X4 U200 ( .A(n550), .B(n537), .Y(SUM[1]) );
  XNOR2X4 U201 ( .A(n551), .B(n425), .Y(SUM[6]) );
  NAND2BX1 U202 ( .AN(n507), .B(n505), .Y(n515) );
  XOR2X4 U203 ( .A(n553), .B(n554), .Y(SUM[3]) );
  XNOR2X4 U204 ( .A(n526), .B(n555), .Y(SUM[11]) );
  XOR2X4 U205 ( .A(n440), .B(n442), .Y(n556) );
  INVX8 U206 ( .A(n556), .Y(SUM[30]) );
  XNOR2X4 U207 ( .A(n462), .B(n559), .Y(SUM[25]) );
  XNOR2X4 U208 ( .A(B[25]), .B(A[25]), .Y(n559) );
  XOR2X2 U209 ( .A(n465), .B(n561), .Y(n560) );
  XNOR2X4 U210 ( .A(B[24]), .B(A[24]), .Y(n561) );
  AOI2BB1X4 U211 ( .A0N(A[25]), .A1N(n462), .B0(n563), .Y(n562) );
  AOI2BB1X4 U212 ( .A0N(n475), .A1N(A[21]), .B0(n565), .Y(n564) );
  XOR2X4 U213 ( .A(n566), .B(n567), .Y(n587) );
  NOR2X2 U214 ( .A(B[28]), .B(A[28]), .Y(n453) );
  AND2X4 U215 ( .A(B[28]), .B(A[28]), .Y(n445) );
  XOR2X4 U216 ( .A(n528), .B(n529), .Y(n590) );
  INVX8 U217 ( .A(B[5]), .Y(n586) );
  NAND2X2 U218 ( .A(B[6]), .B(A[6]), .Y(n426) );
  AND2X4 U219 ( .A(B[2]), .B(A[2]), .Y(n448) );
  AND2X4 U220 ( .A(B[11]), .B(A[11]), .Y(n521) );
  XNOR2X2 U221 ( .A(n477), .B(n475), .Y(SUM[21]) );
endmodule


module hash_core_DW01_add_28 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n514, n515, n516, n517, n518, n519, n520, n521, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n388, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n406, n407, n408,
         n409, n410, n411, n412, n413, n415, n416, n418, n419, n420, n421,
         n422, n424, n425, n427, n428, n430, n431, n433, n434, n435, n438,
         n439, n441, n442, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n355, n356, n357, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n387, n389,
         n390, n405, n414, n417, n423, n426, n429, n432, n436, n469, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513;

  XOR2X4 U6 ( .A(n375), .B(n376), .Y(SUM[7]) );
  AOI21X4 U7 ( .A0(n377), .A1(n508), .B0(n378), .Y(n376) );
  XOR2X4 U9 ( .A(n377), .B(n379), .Y(SUM[6]) );
  OAI21X4 U11 ( .A0(n381), .A1(n382), .B0(n383), .Y(n377) );
  XOR2X4 U12 ( .A(n384), .B(n382), .Y(SUM[5]) );
  XNOR2X4 U20 ( .A(n394), .B(n395), .Y(SUM[31]) );
  XNOR2X4 U24 ( .A(n396), .B(n398), .Y(SUM[30]) );
  OAI2BB1X4 U25 ( .A0N(A[29]), .A1N(n399), .B0(n400), .Y(n396) );
  OAI21X4 U26 ( .A0(A[29]), .A1(n399), .B0(B[29]), .Y(n400) );
  OAI2BB1X4 U31 ( .A0N(A[28]), .A1N(n406), .B0(n407), .Y(n399) );
  OAI21X4 U32 ( .A0(n406), .A1(A[28]), .B0(B[28]), .Y(n407) );
  XNOR2X4 U34 ( .A(n406), .B(n408), .Y(SUM[28]) );
  OAI2BB1X4 U35 ( .A0N(A[27]), .A1N(n409), .B0(n410), .Y(n406) );
  OAI21X4 U36 ( .A0(n409), .A1(A[27]), .B0(B[27]), .Y(n410) );
  OAI2BB1X4 U39 ( .A0N(A[26]), .A1N(n412), .B0(n413), .Y(n409) );
  OAI21X4 U40 ( .A0(n412), .A1(A[26]), .B0(B[26]), .Y(n413) );
  OAI2BB1X4 U43 ( .A0N(A[25]), .A1N(n415), .B0(n416), .Y(n412) );
  OAI21X4 U44 ( .A0(n415), .A1(A[25]), .B0(B[25]), .Y(n416) );
  OAI2BB1X4 U47 ( .A0N(A[24]), .A1N(n418), .B0(n419), .Y(n415) );
  OAI21X4 U48 ( .A0(n418), .A1(A[24]), .B0(B[24]), .Y(n419) );
  OAI2BB1X4 U51 ( .A0N(A[23]), .A1N(n421), .B0(n422), .Y(n418) );
  OAI21X4 U52 ( .A0(n421), .A1(A[23]), .B0(B[23]), .Y(n422) );
  OAI2BB1X4 U55 ( .A0N(A[22]), .A1N(n424), .B0(n425), .Y(n421) );
  OAI21X4 U56 ( .A0(n424), .A1(A[22]), .B0(B[22]), .Y(n425) );
  OAI2BB1X4 U59 ( .A0N(n427), .A1N(A[21]), .B0(n428), .Y(n424) );
  OAI21X4 U60 ( .A0(A[21]), .A1(n427), .B0(B[21]), .Y(n428) );
  OAI2BB1X4 U63 ( .A0N(n430), .A1N(A[20]), .B0(n431), .Y(n427) );
  OAI21X4 U64 ( .A0(n430), .A1(A[20]), .B0(B[20]), .Y(n431) );
  OAI2BB1X4 U67 ( .A0N(A[19]), .A1N(n433), .B0(n434), .Y(n430) );
  OAI21X4 U68 ( .A0(n433), .A1(A[19]), .B0(B[19]), .Y(n434) );
  OAI2BB1X4 U73 ( .A0N(A[18]), .A1N(n438), .B0(n439), .Y(n433) );
  OAI21X4 U74 ( .A0(A[18]), .A1(n438), .B0(B[18]), .Y(n439) );
  OAI2BB1X4 U77 ( .A0N(A[17]), .A1N(n441), .B0(n442), .Y(n438) );
  AOI2BB1X4 U82 ( .A0N(A[16]), .A1N(n417), .B0(n445), .Y(n441) );
  AOI21X4 U83 ( .A0(n444), .A1(A[16]), .B0(B[16]), .Y(n445) );
  OAI2BB1X4 U85 ( .A0N(n448), .A1N(n447), .B0(n449), .Y(n444) );
  XOR2X4 U89 ( .A(n455), .B(n456), .Y(SUM[15]) );
  OR2X4 U93 ( .A(A[15]), .B(B[15]), .Y(n448) );
  NOR2X4 U96 ( .A(A[14]), .B(B[14]), .Y(n450) );
  NAND2X4 U101 ( .A(B[13]), .B(A[13]), .Y(n454) );
  NAND2BX4 U106 ( .AN(n465), .B(n464), .Y(n453) );
  OAI2BB1X4 U108 ( .A0N(n466), .A1N(A[11]), .B0(n467), .Y(n465) );
  XOR2X4 U112 ( .A(n471), .B(n472), .Y(SUM[11]) );
  OAI21X4 U114 ( .A0(n468), .A1(n473), .B0(n470), .Y(n471) );
  XNOR2X4 U115 ( .A(n473), .B(n474), .Y(SUM[10]) );
  NAND2BX4 U119 ( .AN(n369), .B(n365), .Y(n473) );
  OAI2BB1X4 U122 ( .A0N(n426), .A1N(A[8]), .B0(n475), .Y(n372) );
  OAI21X4 U123 ( .A0(n373), .A1(A[8]), .B0(B[8]), .Y(n475) );
  OAI211X2 U124 ( .A0(n476), .A1(n513), .B0(n478), .C0(n477), .Y(n373) );
  AOI2BB1X4 U126 ( .A0N(A[7]), .A1N(B[7]), .B0(n386), .Y(n479) );
  NOR2X4 U127 ( .A(B[4]), .B(A[4]), .Y(n386) );
  OR2X4 U130 ( .A(A[3]), .B(B[3]), .Y(n392) );
  OR2X4 U133 ( .A(B[2]), .B(A[2]), .Y(n404) );
  OAI2BB1X4 U134 ( .A0N(A[1]), .A1N(n423), .B0(n481), .Y(n402) );
  OAI21X4 U135 ( .A0(n435), .A1(A[1]), .B0(B[1]), .Y(n481) );
  OAI2BB1X4 U137 ( .A0N(n513), .A1N(n476), .B0(B[7]), .Y(n477) );
  AOI21X4 U138 ( .A0(n508), .A1(n482), .B0(n378), .Y(n476) );
  AND2X2 U139 ( .A(B[6]), .B(A[6]), .Y(n378) );
  OAI21X4 U140 ( .A0(n388), .A1(n381), .B0(n383), .Y(n482) );
  NAND2X4 U141 ( .A(B[5]), .B(A[5]), .Y(n383) );
  NOR2X4 U142 ( .A(A[5]), .B(B[5]), .Y(n381) );
  NAND2X4 U143 ( .A(B[4]), .B(A[4]), .Y(n388) );
  NOR2X4 U144 ( .A(A[6]), .B(B[6]), .Y(n380) );
  NOR2X4 U147 ( .A(n360), .B(n512), .Y(n435) );
  NAND2BX4 U2 ( .AN(n372), .B(n355), .Y(n359) );
  CLKINVX20 U3 ( .A(n371), .Y(n355) );
  NAND2X4 U4 ( .A(n393), .B(n480), .Y(n385) );
  NAND2X2 U5 ( .A(n436), .B(n470), .Y(n466) );
  INVX2 U8 ( .A(n372), .Y(n387) );
  XNOR2X4 U10 ( .A(n409), .B(n411), .Y(SUM[27]) );
  INVX2 U13 ( .A(n414), .Y(n389) );
  NAND2X4 U14 ( .A(n389), .B(n480), .Y(n356) );
  XNOR2X4 U15 ( .A(n401), .B(n402), .Y(SUM[2]) );
  NAND4X4 U16 ( .A(n385), .B(n509), .C(n508), .D(n479), .Y(n478) );
  AOI21X4 U17 ( .A0(n511), .A1(n356), .B0(n510), .Y(n382) );
  NAND2X1 U18 ( .A(n453), .B(n502), .Y(n460) );
  BUFX8 U19 ( .A(n517), .Y(SUM[17]) );
  XOR2X1 U21 ( .A(n441), .B(n494), .Y(n517) );
  NOR2X2 U22 ( .A(A[12]), .B(B[12]), .Y(n462) );
  NAND2X2 U23 ( .A(B[12]), .B(A[12]), .Y(n464) );
  CLKINVX3 U27 ( .A(n454), .Y(n506) );
  XOR2X1 U28 ( .A(B[11]), .B(A[11]), .Y(n472) );
  NOR2X2 U29 ( .A(A[13]), .B(B[13]), .Y(n459) );
  BUFX3 U30 ( .A(n519), .Y(SUM[12]) );
  INVX1 U33 ( .A(n393), .Y(n414) );
  XNOR2X1 U37 ( .A(A[16]), .B(B[16]), .Y(n446) );
  XOR2X1 U38 ( .A(B[17]), .B(A[17]), .Y(n494) );
  AND2X2 U41 ( .A(n432), .B(n429), .Y(n357) );
  XOR2X4 U42 ( .A(n415), .B(n496), .Y(SUM[25]) );
  OR2X4 U45 ( .A(n363), .B(n371), .Y(n365) );
  INVX4 U46 ( .A(n387), .Y(n363) );
  CLKINVX8 U49 ( .A(B[0]), .Y(n360) );
  INVX4 U50 ( .A(B[0]), .Y(n501) );
  INVX8 U53 ( .A(n491), .Y(SUM[20]) );
  XOR2X1 U54 ( .A(n492), .B(n430), .Y(n491) );
  BUFX2 U57 ( .A(n426), .Y(n361) );
  XOR2XL U58 ( .A(n362), .B(n438), .Y(n516) );
  XOR2X1 U61 ( .A(A[18]), .B(B[18]), .Y(n362) );
  XOR2X4 U62 ( .A(B[1]), .B(A[1]), .Y(n495) );
  OAI21XL U65 ( .A0(n462), .A1(n453), .B0(n463), .Y(n519) );
  XOR2X1 U66 ( .A(n433), .B(n364), .Y(n515) );
  XOR2X1 U69 ( .A(A[19]), .B(B[19]), .Y(n364) );
  AOI21XL U70 ( .A0(n501), .A1(n512), .B0(n435), .Y(n521) );
  XOR2X2 U71 ( .A(n356), .B(n487), .Y(SUM[4]) );
  AND2X4 U72 ( .A(B[9]), .B(A[9]), .Y(n371) );
  AOI31X2 U75 ( .A0(n436), .A1(n470), .A2(n366), .B0(n367), .Y(n368) );
  INVX1 U76 ( .A(A[11]), .Y(n366) );
  INVXL U78 ( .A(B[11]), .Y(n367) );
  INVX4 U79 ( .A(n368), .Y(n467) );
  NAND2X4 U80 ( .A(B[3]), .B(A[3]), .Y(n393) );
  NAND2X4 U81 ( .A(n359), .B(n357), .Y(n436) );
  OR2X2 U84 ( .A(n391), .B(n507), .Y(n405) );
  OAI21X4 U86 ( .A0(n369), .A1(n365), .B0(n370), .Y(SUM[9]) );
  XOR2X4 U87 ( .A(n390), .B(n405), .Y(SUM[3]) );
  AND2X1 U88 ( .A(n392), .B(n393), .Y(n390) );
  BUFX8 U90 ( .A(n516), .Y(SUM[18]) );
  BUFX8 U91 ( .A(n521), .Y(SUM[0]) );
  BUFX8 U92 ( .A(n520), .Y(SUM[1]) );
  XOR2X2 U94 ( .A(n421), .B(n497), .Y(n514) );
  OAI2BB1X4 U95 ( .A0N(n448), .A1N(n447), .B0(n449), .Y(n417) );
  OAI21X4 U97 ( .A0(n451), .A1(n450), .B0(n452), .Y(n447) );
  OAI2BB1X2 U98 ( .A0N(A[30]), .A1N(n396), .B0(n397), .Y(n395) );
  OAI21X4 U99 ( .A0(n396), .A1(A[30]), .B0(B[30]), .Y(n397) );
  OAI21X4 U100 ( .A0(n441), .A1(A[17]), .B0(B[17]), .Y(n442) );
  XNOR2X2 U102 ( .A(n412), .B(n493), .Y(SUM[26]) );
  NOR2X4 U103 ( .A(n501), .B(n512), .Y(n423) );
  OAI211X2 U104 ( .A0(n476), .A1(n513), .B0(n478), .C0(n477), .Y(n426) );
  INVX8 U105 ( .A(n489), .Y(SUM[21]) );
  INVXL U107 ( .A(n468), .Y(n429) );
  INVXL U109 ( .A(n369), .Y(n432) );
  NOR2X1 U110 ( .A(B[10]), .B(A[10]), .Y(n468) );
  NOR2X4 U111 ( .A(A[9]), .B(B[9]), .Y(n369) );
  NAND2X4 U113 ( .A(B[10]), .B(A[10]), .Y(n470) );
  AOI31X2 U116 ( .A0(n505), .A1(n502), .A2(n453), .B0(n506), .Y(n451) );
  BUFX4 U117 ( .A(n518), .Y(SUM[16]) );
  XNOR2X1 U118 ( .A(n417), .B(n446), .Y(n518) );
  BUFX8 U120 ( .A(n515), .Y(SUM[19]) );
  INVX4 U121 ( .A(n514), .Y(n469) );
  INVX8 U125 ( .A(n469), .Y(SUM[23]) );
  XOR2X4 U128 ( .A(n460), .B(n461), .Y(SUM[13]) );
  CLKINVX2 U129 ( .A(n452), .Y(n503) );
  XOR2X4 U131 ( .A(n457), .B(n488), .Y(SUM[14]) );
  NAND2X2 U132 ( .A(B[2]), .B(A[2]), .Y(n403) );
  NOR2XL U136 ( .A(n503), .B(n450), .Y(n488) );
  NAND2XL U145 ( .A(n505), .B(n454), .Y(n461) );
  INVX1 U146 ( .A(n381), .Y(n509) );
  INVXL U148 ( .A(n388), .Y(n510) );
  OAI21X4 U149 ( .A0(n459), .A1(n460), .B0(n454), .Y(n457) );
  NOR2XL U150 ( .A(n386), .B(n510), .Y(n487) );
  NAND2XL U151 ( .A(n403), .B(n404), .Y(n401) );
  XOR2X1 U152 ( .A(n490), .B(n427), .Y(n489) );
  XNOR2X1 U153 ( .A(A[21]), .B(B[21]), .Y(n490) );
  XNOR2X1 U154 ( .A(A[20]), .B(B[20]), .Y(n492) );
  XNOR2X1 U155 ( .A(A[26]), .B(B[26]), .Y(n493) );
  XOR2X1 U156 ( .A(n423), .B(n495), .Y(n520) );
  NAND2X2 U157 ( .A(B[15]), .B(A[15]), .Y(n449) );
  INVXL U158 ( .A(n386), .Y(n511) );
  NOR2BX1 U159 ( .AN(n470), .B(n468), .Y(n474) );
  NAND2XL U160 ( .A(n509), .B(n383), .Y(n384) );
  XOR2X1 U161 ( .A(B[7]), .B(n513), .Y(n375) );
  NAND2X1 U162 ( .A(n448), .B(n449), .Y(n455) );
  AOI21X2 U163 ( .A0(n457), .A1(n504), .B0(n503), .Y(n456) );
  INVXL U164 ( .A(n450), .Y(n504) );
  NOR2XL U165 ( .A(n378), .B(n380), .Y(n379) );
  INVX1 U166 ( .A(n403), .Y(n507) );
  XOR2X1 U167 ( .A(B[8]), .B(A[8]), .Y(n374) );
  XNOR2X1 U168 ( .A(A[24]), .B(B[24]), .Y(n420) );
  XOR2X1 U169 ( .A(A[25]), .B(B[25]), .Y(n496) );
  XNOR2X1 U170 ( .A(A[27]), .B(B[27]), .Y(n411) );
  XOR2X1 U171 ( .A(A[23]), .B(B[23]), .Y(n497) );
  XOR2X1 U172 ( .A(n424), .B(n498), .Y(SUM[22]) );
  XOR2X1 U173 ( .A(A[22]), .B(B[22]), .Y(n498) );
  XNOR2X1 U174 ( .A(A[30]), .B(B[30]), .Y(n398) );
  XNOR2X1 U175 ( .A(A[28]), .B(B[28]), .Y(n408) );
  XNOR2X1 U176 ( .A(B[31]), .B(A[31]), .Y(n394) );
  XNOR2X4 U177 ( .A(n399), .B(n500), .Y(n499) );
  INVX8 U178 ( .A(n499), .Y(SUM[29]) );
  XOR2X1 U179 ( .A(A[29]), .B(B[29]), .Y(n500) );
  NAND2X2 U180 ( .A(B[14]), .B(A[14]), .Y(n452) );
  OAI2BB1XL U181 ( .A0N(n502), .A1N(n464), .B0(n465), .Y(n463) );
  OAI21XL U182 ( .A0(n369), .A1(n371), .B0(n363), .Y(n370) );
  OAI21X4 U183 ( .A0(n391), .A1(n507), .B0(n392), .Y(n480) );
  XOR2X1 U184 ( .A(n361), .B(n374), .Y(SUM[8]) );
  XNOR2X2 U185 ( .A(n418), .B(n420), .Y(SUM[24]) );
  AND2X4 U186 ( .A(n402), .B(n404), .Y(n391) );
  CLKINVX4 U187 ( .A(n462), .Y(n502) );
  CLKINVX4 U188 ( .A(n459), .Y(n505) );
  CLKINVX4 U189 ( .A(n380), .Y(n508) );
  CLKINVX4 U190 ( .A(A[0]), .Y(n512) );
  CLKINVX4 U191 ( .A(A[7]), .Y(n513) );
endmodule


module hash_core_DW01_add_7 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n301, n336, n373, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411;

  NAND2BX4 U25 ( .AN(n287), .B(n288), .Y(n290) );
  NOR2X4 U32 ( .A(B[29]), .B(A[29]), .Y(n291) );
  NAND2X4 U51 ( .A(B[26]), .B(A[26]), .Y(n310) );
  AND2X2 U56 ( .A(B[25]), .B(A[25]), .Y(n309) );
  NAND4X2 U62 ( .A(n325), .B(n255), .C(n229), .D(n326), .Y(n324) );
  AOI21X4 U64 ( .A0(n328), .A1(n253), .B0(n254), .Y(n322) );
  OAI2BB1X4 U65 ( .A0N(n229), .A1N(n329), .B0(n330), .Y(n328) );
  NOR2X4 U70 ( .A(B[23]), .B(A[23]), .Y(n321) );
  NOR2X4 U75 ( .A(B[22]), .B(A[22]), .Y(n327) );
  NOR2X4 U84 ( .A(n403), .B(n252), .Y(n329) );
  NAND3X4 U85 ( .A(n341), .B(n342), .C(n343), .Y(n325) );
  OAI211X2 U86 ( .A0(B[17]), .A1(A[17]), .B0(n344), .C0(n345), .Y(n343) );
  AOI2BB1X4 U88 ( .A0N(B[18]), .A1N(A[18]), .B0(n347), .Y(n345) );
  OAI2BB1X4 U105 ( .A0N(n358), .A1N(A[16]), .B0(n359), .Y(n344) );
  OAI21X4 U106 ( .A0(A[16]), .A1(n358), .B0(B[16]), .Y(n359) );
  AOI31X2 U110 ( .A0(n365), .A1(n366), .A2(n367), .B0(n368), .Y(n364) );
  AOI211X2 U113 ( .A0(n370), .A1(n247), .B0(n248), .C0(n371), .Y(n361) );
  AND2X2 U117 ( .A(B[15]), .B(A[15]), .Y(n368) );
  NOR2X4 U118 ( .A(B[15]), .B(A[15]), .Y(n362) );
  AND2X2 U123 ( .A(B[14]), .B(A[14]), .Y(n371) );
  NOR2X4 U132 ( .A(n408), .B(n246), .Y(n370) );
  OAI211X2 U133 ( .A0(n243), .A1(n245), .B0(n381), .C0(n382), .Y(n366) );
  NOR2X4 U145 ( .A(A[10]), .B(B[10]), .Y(n385) );
  NOR2X4 U148 ( .A(B[9]), .B(A[9]), .Y(n388) );
  OAI211X2 U152 ( .A0(n394), .A1(n262), .B0(n395), .C0(n396), .Y(n266) );
  OAI2BB1X4 U155 ( .A0N(n283), .A1N(A[3]), .B0(n398), .Y(n279) );
  AOI21X4 U163 ( .A0(n401), .A1(n400), .B0(n272), .Y(n394) );
  AND2X2 U164 ( .A(B[6]), .B(A[6]), .Y(n272) );
  NOR2X4 U167 ( .A(B[5]), .B(A[5]), .Y(n275) );
  AOI21X4 U2 ( .A0(n257), .A1(n317), .B0(n309), .Y(n315) );
  OAI21X2 U3 ( .A0(n305), .A1(n315), .B0(n310), .Y(n313) );
  NOR2BX4 U4 ( .AN(n307), .B(n306), .Y(n314) );
  XOR2X4 U5 ( .A(n313), .B(n314), .Y(SUM[27]) );
  OR2X4 U6 ( .A(A[28]), .B(B[28]), .Y(n226) );
  NAND2X2 U7 ( .A(A[28]), .B(B[28]), .Y(n292) );
  NOR2BX2 U8 ( .AN(n292), .B(n228), .Y(n303) );
  XOR2X4 U9 ( .A(n303), .B(n302), .Y(SUM[28]) );
  NOR2BX4 U10 ( .AN(n227), .B(A[30]), .Y(n287) );
  CLKINVX20 U11 ( .A(B[30]), .Y(n227) );
  NOR2XL U12 ( .A(B[28]), .B(A[28]), .Y(n228) );
  NAND3X1 U13 ( .A(n238), .B(n239), .C(n294), .Y(n289) );
  NAND2XL U14 ( .A(n293), .B(n292), .Y(n299) );
  INVX1 U15 ( .A(B[29]), .Y(n232) );
  CLKINVX3 U16 ( .A(n310), .Y(n258) );
  INVX1 U17 ( .A(B[27]), .Y(n233) );
  INVXL U18 ( .A(n329), .Y(n231) );
  XOR2X2 U19 ( .A(n299), .B(n300), .Y(SUM[29]) );
  OAI21X2 U20 ( .A0(n385), .A1(n386), .B0(n387), .Y(n384) );
  INVXL U21 ( .A(n230), .Y(n337) );
  OR2X4 U22 ( .A(B[21]), .B(A[21]), .Y(n229) );
  OAI2BB1X1 U23 ( .A0N(n325), .A1N(n339), .B0(n231), .Y(n230) );
  OAI2BB1X4 U24 ( .A0N(n229), .A1N(n230), .B0(n330), .Y(n333) );
  XOR2X1 U26 ( .A(n338), .B(n337), .Y(SUM[21]) );
  AOI21X1 U27 ( .A0(n333), .A1(n253), .B0(n254), .Y(n332) );
  XNOR2X1 U28 ( .A(n335), .B(n333), .Y(SUM[22]) );
  INVX8 U29 ( .A(n321), .Y(n255) );
  NAND2X4 U30 ( .A(n240), .B(n312), .Y(n317) );
  OAI31X4 U31 ( .A0(n361), .A1(n362), .A2(n363), .B0(n364), .Y(n358) );
  NAND2X4 U33 ( .A(B[30]), .B(A[30]), .Y(n288) );
  NAND2BX4 U34 ( .AN(n232), .B(A[29]), .Y(n294) );
  NOR2BX4 U35 ( .AN(n233), .B(A[27]), .Y(n306) );
  NOR2BX2 U36 ( .AN(n294), .B(n291), .Y(n300) );
  NAND2X4 U37 ( .A(n226), .B(n236), .Y(n293) );
  OAI221X2 U38 ( .A0(n321), .A1(n322), .B0(n234), .B1(n235), .C0(n324), .Y(
        n319) );
  INVXL U39 ( .A(A[23]), .Y(n234) );
  INVX1 U40 ( .A(B[23]), .Y(n235) );
  XOR2X4 U41 ( .A(A[31]), .B(B[31]), .Y(n286) );
  NAND2X1 U42 ( .A(B[18]), .B(A[18]), .Y(n348) );
  XOR2X1 U43 ( .A(n355), .B(n353), .Y(SUM[18]) );
  NAND2X2 U44 ( .A(B[27]), .B(A[27]), .Y(n307) );
  XNOR2X4 U45 ( .A(n290), .B(n289), .Y(SUM[30]) );
  OAI31X2 U46 ( .A0(n304), .A1(n305), .A2(n306), .B0(n307), .Y(n236) );
  AND3X4 U47 ( .A(n238), .B(n239), .C(n294), .Y(n237) );
  OAI31X4 U48 ( .A0(n304), .A1(n305), .A2(n306), .B0(n307), .Y(n302) );
  OR2X4 U49 ( .A(n291), .B(n292), .Y(n238) );
  OR2X4 U50 ( .A(n291), .B(n293), .Y(n239) );
  OAI21X4 U52 ( .A0(n237), .A1(n287), .B0(n288), .Y(n285) );
  XOR2X4 U53 ( .A(n285), .B(n286), .Y(SUM[31]) );
  NOR3X4 U54 ( .A(n308), .B(n258), .C(n309), .Y(n304) );
  INVX4 U55 ( .A(n348), .Y(n251) );
  OAI21X2 U57 ( .A0(n251), .A1(n346), .B0(n345), .Y(n341) );
  NOR2X4 U58 ( .A(B[13]), .B(A[13]), .Y(n369) );
  NAND2XL U59 ( .A(B[13]), .B(A[13]), .Y(n372) );
  INVX4 U60 ( .A(A[24]), .Y(n256) );
  INVX1 U61 ( .A(B[24]), .Y(n404) );
  OAI21X4 U63 ( .A0(B[24]), .A1(A[24]), .B0(n319), .Y(n312) );
  OR2X2 U66 ( .A(n256), .B(n404), .Y(n240) );
  INVXL U67 ( .A(n311), .Y(n257) );
  NOR2XL U68 ( .A(n309), .B(n311), .Y(n318) );
  OAI21X2 U69 ( .A0(A[3]), .A1(n283), .B0(B[3]), .Y(n398) );
  NOR2X4 U71 ( .A(A[25]), .B(B[25]), .Y(n311) );
  OAI2BB1X4 U72 ( .A0N(n262), .A1N(n394), .B0(B[7]), .Y(n395) );
  NAND4X1 U73 ( .A(n279), .B(n401), .C(n373), .D(n397), .Y(n396) );
  AOI22X4 U74 ( .A0(n245), .A1(n409), .B0(n261), .B1(n411), .Y(n383) );
  NAND2X2 U76 ( .A(B[5]), .B(A[5]), .Y(n277) );
  NAND2X1 U77 ( .A(B[2]), .B(A[2]), .Y(n298) );
  INVX4 U78 ( .A(A[7]), .Y(n262) );
  AOI21X4 U79 ( .A0(n252), .A1(n403), .B0(n327), .Y(n326) );
  AOI21X2 U80 ( .A0(n268), .A1(n259), .B0(n260), .Y(n386) );
  NOR2X4 U81 ( .A(n411), .B(n261), .Y(n268) );
  INVX4 U82 ( .A(A[17]), .Y(n250) );
  NOR2X4 U83 ( .A(n362), .B(n369), .Y(n365) );
  OAI21X4 U87 ( .A0(n297), .A1(n296), .B0(n298), .Y(n283) );
  NOR2X2 U89 ( .A(n406), .B(n336), .Y(n349) );
  CLKINVX4 U90 ( .A(n274), .Y(n401) );
  INVX4 U91 ( .A(A[4]), .Y(n402) );
  CLKINVX4 U92 ( .A(n275), .Y(n373) );
  OAI21X1 U93 ( .A0(n369), .A1(n377), .B0(n372), .Y(n375) );
  XNOR2X1 U94 ( .A(n241), .B(n374), .Y(SUM[15]) );
  NOR2XL U95 ( .A(n362), .B(n368), .Y(n241) );
  AOI21XL U96 ( .A0(n250), .A1(n405), .B0(n346), .Y(n357) );
  XOR2XL U97 ( .A(n263), .B(n264), .Y(SUM[9]) );
  XOR2XL U98 ( .A(n295), .B(n296), .Y(SUM[2]) );
  NAND2BXL U99 ( .AN(n297), .B(n298), .Y(n295) );
  AOI21XL U100 ( .A0(n406), .A1(n336), .B0(n349), .Y(SUM[0]) );
  NOR2X4 U101 ( .A(B[14]), .B(A[14]), .Y(n363) );
  NAND2X4 U102 ( .A(B[9]), .B(A[9]), .Y(n265) );
  NAND2X1 U103 ( .A(B[10]), .B(A[10]), .Y(n387) );
  CLKINVX2 U104 ( .A(n399), .Y(n301) );
  INVX1 U107 ( .A(A[8]), .Y(n261) );
  INVX2 U108 ( .A(A[11]), .Y(n245) );
  INVX4 U109 ( .A(A[20]), .Y(n252) );
  INVX1 U111 ( .A(A[0]), .Y(n336) );
  AOI21XL U112 ( .A0(n246), .A1(n408), .B0(n363), .Y(n367) );
  INVX1 U114 ( .A(n265), .Y(n260) );
  INVX1 U115 ( .A(n369), .Y(n247) );
  NOR2X1 U116 ( .A(n405), .B(n250), .Y(n346) );
  INVXL U119 ( .A(n385), .Y(n242) );
  OAI2BB1X2 U120 ( .A0N(n281), .A1N(n373), .B0(n277), .Y(n400) );
  XOR2X1 U121 ( .A(n319), .B(n320), .Y(SUM[24]) );
  XNOR2XL U122 ( .A(n404), .B(A[24]), .Y(n320) );
  XOR2X1 U124 ( .A(n317), .B(n318), .Y(SUM[25]) );
  XOR2X1 U125 ( .A(n316), .B(n315), .Y(SUM[26]) );
  NAND2BXL U126 ( .AN(n305), .B(n310), .Y(n316) );
  INVX1 U127 ( .A(n372), .Y(n248) );
  AOI21XL U128 ( .A0(n344), .A1(n356), .B0(n346), .Y(n353) );
  NAND2X1 U129 ( .A(n250), .B(n405), .Y(n356) );
  NAND2XL U130 ( .A(n252), .B(n403), .Y(n339) );
  NOR2X1 U131 ( .A(n407), .B(n402), .Y(n281) );
  XOR2X1 U134 ( .A(n331), .B(n332), .Y(SUM[23]) );
  NAND2XL U135 ( .A(n255), .B(n323), .Y(n331) );
  XNOR2X1 U136 ( .A(n376), .B(n375), .Y(SUM[14]) );
  NAND2BXL U137 ( .AN(n371), .B(n249), .Y(n376) );
  NAND2XL U138 ( .A(n253), .B(n334), .Y(n335) );
  XOR2X1 U139 ( .A(n325), .B(n340), .Y(SUM[20]) );
  AOI21XL U140 ( .A0(n252), .A1(n403), .B0(n329), .Y(n340) );
  XOR2X1 U141 ( .A(n344), .B(n357), .Y(SUM[17]) );
  NAND2XL U142 ( .A(n229), .B(n330), .Y(n338) );
  AOI21XL U143 ( .A0(n375), .A1(n249), .B0(n371), .Y(n374) );
  OAI21XL U144 ( .A0(n264), .A1(n388), .B0(n265), .Y(n391) );
  INVX1 U146 ( .A(n363), .Y(n249) );
  XOR2X1 U147 ( .A(n391), .B(n392), .Y(SUM[10]) );
  NOR2XL U149 ( .A(n385), .B(n244), .Y(n392) );
  XOR2X1 U150 ( .A(n378), .B(n377), .Y(SUM[13]) );
  NAND2XL U151 ( .A(n247), .B(n372), .Y(n378) );
  XOR2X1 U153 ( .A(n366), .B(n380), .Y(SUM[12]) );
  AOI21XL U154 ( .A0(n246), .A1(n408), .B0(n370), .Y(n380) );
  AOI21XL U156 ( .A0(n279), .A1(n280), .B0(n281), .Y(n276) );
  NAND2XL U157 ( .A(n402), .B(n407), .Y(n280) );
  OAI21XL U158 ( .A0(n275), .A1(n276), .B0(n277), .Y(n271) );
  INVX1 U159 ( .A(n387), .Y(n244) );
  XOR2X1 U160 ( .A(n266), .B(n267), .Y(SUM[8]) );
  AOI21XL U161 ( .A0(n261), .A1(n411), .B0(n268), .Y(n267) );
  XOR2X1 U162 ( .A(n271), .B(n273), .Y(SUM[6]) );
  NOR2XL U165 ( .A(n274), .B(n272), .Y(n273) );
  NAND2XL U166 ( .A(n259), .B(n265), .Y(n263) );
  XOR2X1 U168 ( .A(n279), .B(n282), .Y(SUM[4]) );
  AOI21XL U169 ( .A0(n402), .A1(n407), .B0(n281), .Y(n282) );
  XOR2X1 U170 ( .A(n278), .B(n276), .Y(SUM[5]) );
  NAND2XL U171 ( .A(n373), .B(n277), .Y(n278) );
  OAI21XL U172 ( .A0(A[11]), .A1(n384), .B0(B[11]), .Y(n381) );
  NAND4X1 U173 ( .A(n266), .B(n242), .C(n259), .D(n383), .Y(n382) );
  INVX1 U174 ( .A(n384), .Y(n243) );
  NOR2X2 U175 ( .A(B[26]), .B(A[26]), .Y(n305) );
  NOR2X1 U176 ( .A(B[19]), .B(A[19]), .Y(n347) );
  NAND2X1 U177 ( .A(B[21]), .B(A[21]), .Y(n330) );
  INVX1 U178 ( .A(B[11]), .Y(n409) );
  NAND2XL U179 ( .A(B[23]), .B(A[23]), .Y(n323) );
  NOR2X2 U180 ( .A(B[2]), .B(A[2]), .Y(n297) );
  NOR2X2 U181 ( .A(A[6]), .B(B[6]), .Y(n274) );
  AOI22X1 U182 ( .A0(n402), .A1(n407), .B0(n262), .B1(n410), .Y(n397) );
  INVX1 U183 ( .A(B[7]), .Y(n410) );
  NAND2XL U184 ( .A(B[19]), .B(A[19]), .Y(n342) );
  NOR2BXL U185 ( .AN(n379), .B(n370), .Y(n377) );
  OAI21XL U186 ( .A0(A[12]), .A1(B[12]), .B0(n366), .Y(n379) );
  XOR2X1 U187 ( .A(n358), .B(n360), .Y(SUM[16]) );
  XOR2XL U188 ( .A(B[16]), .B(A[16]), .Y(n360) );
  OAI21XL U189 ( .A0(B[18]), .A1(A[18]), .B0(n348), .Y(n355) );
  XOR2X2 U190 ( .A(n351), .B(n352), .Y(SUM[19]) );
  NOR2BXL U191 ( .AN(n342), .B(n347), .Y(n352) );
  OAI21XL U192 ( .A0(n353), .A1(n354), .B0(n348), .Y(n351) );
  NOR2XL U193 ( .A(A[18]), .B(B[18]), .Y(n354) );
  AOI21X1 U194 ( .A0(n349), .A1(A[1]), .B0(n301), .Y(n296) );
  OAI21X1 U195 ( .A0(n349), .A1(A[1]), .B0(B[1]), .Y(n399) );
  NOR2BXL U196 ( .AN(n393), .B(n268), .Y(n264) );
  OAI21XL U197 ( .A0(A[8]), .A1(B[8]), .B0(n266), .Y(n393) );
  XOR2X1 U198 ( .A(n389), .B(n390), .Y(SUM[11]) );
  XNOR2XL U199 ( .A(B[11]), .B(A[11]), .Y(n389) );
  AOI21XL U200 ( .A0(n391), .A1(n242), .B0(n244), .Y(n390) );
  INVX1 U201 ( .A(B[4]), .Y(n407) );
  INVX1 U202 ( .A(B[0]), .Y(n406) );
  XOR2X1 U203 ( .A(n269), .B(n270), .Y(SUM[7]) );
  XNOR2XL U204 ( .A(B[7]), .B(A[7]), .Y(n269) );
  AOI21XL U205 ( .A0(n271), .A1(n401), .B0(n272), .Y(n270) );
  INVX1 U206 ( .A(B[8]), .Y(n411) );
  XOR2X1 U207 ( .A(n283), .B(n284), .Y(SUM[3]) );
  XOR2XL U208 ( .A(B[3]), .B(A[3]), .Y(n284) );
  INVX1 U209 ( .A(B[12]), .Y(n408) );
  XOR2X1 U210 ( .A(n349), .B(n350), .Y(SUM[1]) );
  XOR2XL U211 ( .A(B[1]), .B(A[1]), .Y(n350) );
  INVX1 U212 ( .A(B[20]), .Y(n403) );
  INVX1 U213 ( .A(B[17]), .Y(n405) );
  OAI32X2 U214 ( .A0(n404), .A1(n311), .A2(n256), .B0(n311), .B1(n312), .Y(
        n308) );
  NAND2X2 U215 ( .A(B[22]), .B(A[22]), .Y(n334) );
  CLKINVX4 U216 ( .A(A[12]), .Y(n246) );
  CLKINVX4 U217 ( .A(n327), .Y(n253) );
  CLKINVX4 U218 ( .A(n334), .Y(n254) );
  CLKINVX4 U219 ( .A(n388), .Y(n259) );
endmodule


module hash_core_DW01_add_9 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n449, n271, n272, n273, n274, n275, n276, n277, n278, n279, n282,
         n283, n285, n286, n287, n288, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n327, n328, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n368, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n383, n384, n385, n386, n388, n389, n390, n391,
         n392, n394, n396, n398, n399, n401, n402, n403, n404, n405, n406,
         n407, n408, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n280,
         n281, n284, n289, n311, n326, n329, n330, n367, n369, n382, n387,
         n393, n395, n397, n400, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448;

  XOR2X4 U6 ( .A(n275), .B(n276), .Y(SUM[7]) );
  AOI21X4 U14 ( .A0(n285), .A1(n442), .B0(n286), .Y(n282) );
  XOR2X4 U19 ( .A(n291), .B(n292), .Y(SUM[31]) );
  XNOR2X4 U22 ( .A(B[31]), .B(A[31]), .Y(n291) );
  OAI211X2 U24 ( .A0(n264), .A1(n298), .B0(n299), .C0(n300), .Y(n293) );
  OAI21X4 U27 ( .A0(B[30]), .A1(A[30]), .B0(n295), .Y(n296) );
  NAND2X4 U28 ( .A(B[30]), .B(A[30]), .Y(n295) );
  AOI21X4 U32 ( .A0(n313), .A1(n302), .B0(n434), .Y(n312) );
  NOR2X4 U35 ( .A(A[29]), .B(B[29]), .Y(n297) );
  XNOR2X4 U36 ( .A(n314), .B(n313), .Y(SUM[28]) );
  NAND2X4 U37 ( .A(n304), .B(n315), .Y(n313) );
  OAI211X2 U41 ( .A0(B[24]), .A1(A[24]), .B0(n253), .C0(n317), .Y(n305) );
  NOR2X4 U42 ( .A(n321), .B(n281), .Y(n317) );
  XOR2X4 U46 ( .A(n323), .B(n324), .Y(SUM[27]) );
  AOI21X4 U47 ( .A0(n325), .A1(n433), .B0(n240), .Y(n324) );
  NOR2X4 U53 ( .A(B[26]), .B(A[26]), .Y(n321) );
  OAI21X4 U55 ( .A0(n281), .A1(n327), .B0(n319), .Y(n325) );
  XOR2X4 U56 ( .A(n327), .B(n328), .Y(SUM[25]) );
  XOR2X4 U69 ( .A(n340), .B(n341), .Y(SUM[23]) );
  NAND2X4 U75 ( .A(n431), .B(n446), .Y(n336) );
  XOR2X4 U77 ( .A(n245), .B(n346), .Y(SUM[21]) );
  AOI21X4 U78 ( .A0(n334), .A1(n347), .B0(n337), .Y(n345) );
  NOR2X4 U82 ( .A(B[21]), .B(A[21]), .Y(n344) );
  XOR2X4 U83 ( .A(n334), .B(n348), .Y(SUM[20]) );
  OAI2BB1X4 U84 ( .A0N(n243), .A1N(A[19]), .B0(n350), .Y(n334) );
  AOI211X2 U87 ( .A0(n355), .A1(n356), .B0(n357), .C0(n427), .Y(n351) );
  NOR2X4 U89 ( .A(n428), .B(n445), .Y(n337) );
  XOR2X4 U92 ( .A(n362), .B(n363), .Y(SUM[19]) );
  OAI21X4 U94 ( .A0(n353), .A1(n364), .B0(n354), .Y(n362) );
  XOR2X4 U95 ( .A(n365), .B(n364), .Y(SUM[18]) );
  AOI2BB1X4 U96 ( .A0N(n366), .A1N(n352), .B0(n357), .Y(n364) );
  AND2X2 U103 ( .A(B[17]), .B(A[17]), .Y(n357) );
  OAI211X2 U108 ( .A0(n422), .A1(n376), .B0(n377), .C0(n378), .Y(n374) );
  XOR2X4 U112 ( .A(n379), .B(n380), .Y(SUM[15]) );
  AND2X2 U120 ( .A(B[14]), .B(A[14]), .Y(n375) );
  OAI21X4 U121 ( .A0(n383), .A1(n384), .B0(n378), .Y(n381) );
  XOR2X4 U122 ( .A(n385), .B(n384), .Y(SUM[13]) );
  AOI2BB1X4 U123 ( .A0N(n422), .A1N(n376), .B0(n424), .Y(n384) );
  AOI21X4 U138 ( .A0(n399), .A1(n423), .B0(n409), .Y(n398) );
  OAI21X4 U144 ( .A0(n271), .A1(n280), .B0(n268), .Y(n399) );
  AOI211X2 U150 ( .A0(n402), .A1(A[7]), .B0(n440), .C0(n403), .Y(n401) );
  OAI21X4 U154 ( .A0(n290), .A1(n448), .B0(n405), .Y(n285) );
  AOI21X4 U156 ( .A0(n443), .A1(n307), .B0(n310), .Y(n290) );
  OAI21X4 U163 ( .A0(n407), .A1(n277), .B0(n279), .Y(n402) );
  AOI21X4 U165 ( .A0(n286), .A1(n246), .B0(n283), .Y(n407) );
  AND2X2 U168 ( .A(B[4]), .B(A[4]), .Y(n286) );
  CLKINVX4 U170 ( .A(n408), .Y(SUM[0]) );
  INVX2 U2 ( .A(n356), .Y(n393) );
  INVX8 U3 ( .A(n349), .Y(n266) );
  NAND3X1 U4 ( .A(n304), .B(n306), .C(n305), .Y(n301) );
  CLKINVX4 U5 ( .A(B[5]), .Y(n262) );
  INVX4 U7 ( .A(n262), .Y(n263) );
  BUFX8 U8 ( .A(n318), .Y(n240) );
  NAND3X2 U9 ( .A(n429), .B(n334), .C(n335), .Y(n333) );
  INVX2 U10 ( .A(n439), .Y(n249) );
  XOR2X2 U11 ( .A(n439), .B(n273), .Y(n449) );
  BUFX4 U12 ( .A(n283), .Y(n242) );
  OR2X4 U13 ( .A(n283), .B(n251), .Y(n415) );
  AOI2BB1X4 U15 ( .A0N(n252), .A1N(n241), .B0(n260), .Y(n327) );
  CLKINVX20 U16 ( .A(A[24]), .Y(n241) );
  CLKINVX8 U17 ( .A(n252), .Y(n253) );
  INVX4 U18 ( .A(n320), .Y(n252) );
  CLKINVX4 U20 ( .A(n351), .Y(n289) );
  INVX4 U21 ( .A(n266), .Y(n243) );
  XOR2X4 U23 ( .A(n244), .B(n284), .Y(SUM[22]) );
  CLKINVX20 U25 ( .A(n343), .Y(n244) );
  OAI21X4 U26 ( .A0(B[23]), .A1(A[23]), .B0(n336), .Y(n332) );
  AOI21X2 U29 ( .A0(n423), .A1(n394), .B0(n409), .Y(n388) );
  NOR2X1 U30 ( .A(n395), .B(n409), .Y(n400) );
  OAI2BB1X2 U31 ( .A0N(n444), .A1N(n388), .B0(B[11]), .Y(n389) );
  INVX3 U33 ( .A(n249), .Y(n250) );
  BUFX4 U34 ( .A(n342), .Y(n284) );
  AOI21X2 U38 ( .A0(n334), .A1(n347), .B0(n337), .Y(n245) );
  AOI21X4 U39 ( .A0(n445), .A1(n428), .B0(n332), .Y(n335) );
  AOI211X1 U40 ( .A0(n337), .A1(n429), .B0(n338), .C0(n430), .Y(n331) );
  INVX4 U43 ( .A(B[22]), .Y(n431) );
  INVX2 U44 ( .A(A[22]), .Y(n446) );
  CLKINVX3 U45 ( .A(n259), .Y(n391) );
  INVXL U48 ( .A(B[24]), .Y(n261) );
  OAI21X2 U49 ( .A0(n360), .A1(n358), .B0(n361), .Y(n307) );
  INVX2 U50 ( .A(A[20]), .Y(n445) );
  INVX2 U51 ( .A(n277), .Y(n441) );
  NOR2X2 U52 ( .A(n263), .B(A[5]), .Y(n251) );
  NAND2X2 U54 ( .A(n429), .B(n339), .Y(n346) );
  INVX2 U57 ( .A(n298), .Y(n434) );
  XNOR2X2 U58 ( .A(n410), .B(n393), .Y(SUM[16]) );
  AND2X2 U59 ( .A(n355), .B(n368), .Y(n410) );
  NAND2BX2 U60 ( .AN(n338), .B(n336), .Y(n343) );
  XOR2X2 U61 ( .A(n358), .B(n359), .Y(SUM[1]) );
  INVX2 U62 ( .A(n449), .Y(n269) );
  OR2X4 U63 ( .A(n263), .B(A[5]), .Y(n246) );
  INVX2 U64 ( .A(n254), .Y(n280) );
  AND2X4 U65 ( .A(n303), .B(n302), .Y(n247) );
  XOR2X4 U66 ( .A(n419), .B(n253), .Y(SUM[24]) );
  XNOR2X4 U67 ( .A(n381), .B(n248), .Y(SUM[14]) );
  OR2X2 U68 ( .A(n375), .B(n371), .Y(n248) );
  AOI2BB1X4 U70 ( .A0N(n320), .A1N(A[24]), .B0(n261), .Y(n260) );
  AOI2BB1X1 U71 ( .A0N(A[7]), .A1N(B[7]), .B0(n287), .Y(n404) );
  AND4X2 U72 ( .A(n246), .B(n285), .C(n441), .D(n404), .Y(n403) );
  NAND2X4 U73 ( .A(B[25]), .B(A[25]), .Y(n319) );
  INVX2 U74 ( .A(n321), .Y(n433) );
  OAI221X2 U76 ( .A0(n331), .A1(n332), .B0(n447), .B1(n432), .C0(n333), .Y(
        n320) );
  AOI21X2 U79 ( .A0(n356), .A1(n355), .B0(n427), .Y(n366) );
  OR2X4 U80 ( .A(B[16]), .B(A[16]), .Y(n355) );
  INVX2 U81 ( .A(n295), .Y(n436) );
  NOR2X2 U85 ( .A(B[6]), .B(A[6]), .Y(n277) );
  NAND2X2 U86 ( .A(B[13]), .B(A[13]), .Y(n378) );
  NOR2X2 U88 ( .A(B[13]), .B(A[13]), .Y(n383) );
  INVX8 U90 ( .A(n386), .Y(n422) );
  INVX1 U91 ( .A(n377), .Y(n424) );
  NAND2X2 U93 ( .A(B[12]), .B(A[12]), .Y(n377) );
  OR2X2 U97 ( .A(B[9]), .B(A[9]), .Y(n254) );
  NAND2BX1 U98 ( .AN(B[12]), .B(n255), .Y(n256) );
  INVXL U99 ( .A(A[12]), .Y(n255) );
  INVX4 U100 ( .A(n256), .Y(n376) );
  OR2X4 U101 ( .A(n257), .B(n258), .Y(n396) );
  INVXL U102 ( .A(B[8]), .Y(n257) );
  INVXL U104 ( .A(A[8]), .Y(n258) );
  NAND4X2 U105 ( .A(n437), .B(n250), .C(n254), .D(n391), .Y(n390) );
  AOI21X4 U106 ( .A0(n439), .A1(n437), .B0(n438), .Y(n271) );
  INVX3 U107 ( .A(n396), .Y(n438) );
  OAI21X4 U109 ( .A0(A[11]), .A1(B[11]), .B0(n423), .Y(n259) );
  BUFX4 U110 ( .A(n392), .Y(n395) );
  INVX8 U111 ( .A(n395), .Y(n423) );
  XOR2X2 U113 ( .A(n422), .B(n397), .Y(SUM[12]) );
  AND2X4 U114 ( .A(n263), .B(A[5]), .Y(n283) );
  INVX4 U115 ( .A(n406), .Y(n440) );
  BUFX3 U116 ( .A(n272), .Y(n268) );
  OAI21X2 U117 ( .A0(n396), .A1(n280), .B0(n268), .Y(n394) );
  NAND2X2 U118 ( .A(B[27]), .B(A[27]), .Y(n304) );
  NOR2XL U119 ( .A(B[10]), .B(A[10]), .Y(n392) );
  OAI2BB1X4 U124 ( .A0N(n305), .A1N(n306), .B0(n303), .Y(n315) );
  OAI211X2 U125 ( .A0(n388), .A1(n444), .B0(n389), .C0(n390), .Y(n386) );
  NOR2X2 U126 ( .A(B[2]), .B(A[2]), .Y(n309) );
  INVX4 U127 ( .A(n342), .Y(n330) );
  AOI21X4 U128 ( .A0(n421), .A1(n294), .B0(n436), .Y(n292) );
  INVX8 U129 ( .A(n420), .Y(SUM[30]) );
  NAND2X2 U130 ( .A(B[29]), .B(A[29]), .Y(n299) );
  NAND2X4 U131 ( .A(B[28]), .B(A[28]), .Y(n298) );
  NOR2X2 U132 ( .A(B[25]), .B(A[25]), .Y(n322) );
  INVX4 U133 ( .A(n274), .Y(n437) );
  NOR2X1 U134 ( .A(n274), .B(n438), .Y(n273) );
  NOR2X2 U135 ( .A(B[8]), .B(A[8]), .Y(n274) );
  INVXL U136 ( .A(n339), .Y(n430) );
  NAND2X2 U137 ( .A(B[21]), .B(A[21]), .Y(n339) );
  OAI21X4 U139 ( .A0(n345), .A1(n344), .B0(n339), .Y(n342) );
  INVX2 U140 ( .A(n435), .Y(n264) );
  INVX8 U141 ( .A(n297), .Y(n435) );
  OR2X4 U142 ( .A(A[30]), .B(B[30]), .Y(n294) );
  OAI2BB1X2 U143 ( .A0N(n448), .A1N(n290), .B0(B[3]), .Y(n405) );
  NAND3X4 U145 ( .A(n247), .B(n435), .C(n301), .Y(n300) );
  OR2X4 U146 ( .A(B[28]), .B(A[28]), .Y(n302) );
  AND2X1 U147 ( .A(B[2]), .B(A[2]), .Y(n310) );
  AOI21X4 U148 ( .A0(n316), .A1(n317), .B0(n240), .Y(n306) );
  OR2X4 U149 ( .A(n318), .B(n321), .Y(n414) );
  AND2X4 U151 ( .A(B[26]), .B(A[26]), .Y(n318) );
  OAI21X2 U152 ( .A0(A[7]), .A1(n402), .B0(B[7]), .Y(n406) );
  NAND2X4 U153 ( .A(n265), .B(n266), .Y(n267) );
  NAND2X4 U155 ( .A(n267), .B(B[19]), .Y(n350) );
  INVX12 U157 ( .A(A[19]), .Y(n265) );
  OR2X4 U158 ( .A(A[27]), .B(B[27]), .Y(n303) );
  INVX4 U159 ( .A(n269), .Y(SUM[8]) );
  OAI2BB1X2 U160 ( .A0N(B[24]), .A1N(A[24]), .B0(n319), .Y(n316) );
  OR2X4 U161 ( .A(n286), .B(n287), .Y(n288) );
  INVX4 U162 ( .A(n287), .Y(n442) );
  NOR2X4 U164 ( .A(B[4]), .B(A[4]), .Y(n287) );
  NAND2X4 U166 ( .A(n303), .B(n304), .Y(n323) );
  AOI21X2 U167 ( .A0(n428), .A1(n445), .B0(n337), .Y(n348) );
  INVX12 U169 ( .A(B[20]), .Y(n428) );
  BUFX4 U171 ( .A(n322), .Y(n281) );
  NAND2X4 U172 ( .A(B[6]), .B(A[6]), .Y(n279) );
  NOR2X4 U173 ( .A(n431), .B(n446), .Y(n338) );
  NAND3X4 U174 ( .A(n289), .B(n311), .C(n326), .Y(n329) );
  NAND2X4 U175 ( .A(n329), .B(n354), .Y(n349) );
  CLKINVXL U176 ( .A(n352), .Y(n311) );
  INVXL U177 ( .A(n353), .Y(n326) );
  NOR2X4 U178 ( .A(B[17]), .B(A[17]), .Y(n352) );
  NOR2X4 U179 ( .A(B[18]), .B(A[18]), .Y(n353) );
  NAND2X4 U180 ( .A(B[18]), .B(A[18]), .Y(n354) );
  NOR2X1 U181 ( .A(n277), .B(n278), .Y(n382) );
  NOR2X4 U182 ( .A(n330), .B(n367), .Y(n369) );
  NOR2X4 U183 ( .A(n369), .B(n338), .Y(n341) );
  INVXL U184 ( .A(n336), .Y(n367) );
  INVXL U185 ( .A(n279), .Y(n387) );
  OR2X4 U186 ( .A(n382), .B(n387), .Y(n275) );
  AOI2BB1X4 U187 ( .A0N(n251), .A1N(n282), .B0(n242), .Y(n278) );
  NAND2X2 U188 ( .A(n445), .B(n428), .Y(n347) );
  AND2X2 U189 ( .A(n254), .B(n268), .Y(n412) );
  INVX4 U190 ( .A(n368), .Y(n427) );
  NAND2X2 U191 ( .A(n298), .B(n302), .Y(n314) );
  OR2X1 U192 ( .A(n376), .B(n424), .Y(n397) );
  XNOR2X4 U193 ( .A(n288), .B(n285), .Y(SUM[4]) );
  NOR2XL U194 ( .A(B[1]), .B(A[1]), .Y(n360) );
  XOR2X4 U195 ( .A(n399), .B(n400), .Y(SUM[10]) );
  XNOR2X4 U196 ( .A(n271), .B(n412), .Y(SUM[9]) );
  AND2X2 U197 ( .A(n435), .B(n299), .Y(n416) );
  NAND2BX4 U198 ( .AN(n281), .B(n319), .Y(n328) );
  NOR2XL U199 ( .A(B[14]), .B(A[14]), .Y(n371) );
  AND2X1 U200 ( .A(B[10]), .B(A[10]), .Y(n409) );
  NAND2XL U201 ( .A(B[9]), .B(A[9]), .Y(n272) );
  INVXL U202 ( .A(n371), .Y(n426) );
  NAND2BXL U203 ( .AN(n372), .B(n373), .Y(n379) );
  XOR2X4 U204 ( .A(n398), .B(n411), .Y(SUM[11]) );
  XOR2X1 U205 ( .A(B[11]), .B(n444), .Y(n411) );
  XNOR2XL U206 ( .A(n448), .B(B[3]), .Y(n418) );
  NAND2X1 U207 ( .A(n425), .B(n378), .Y(n385) );
  INVX1 U208 ( .A(n309), .Y(n443) );
  XNOR2X2 U209 ( .A(n413), .B(n278), .Y(SUM[6]) );
  AND2X1 U210 ( .A(n441), .B(n279), .Y(n413) );
  INVX1 U211 ( .A(n383), .Y(n425) );
  XOR2X1 U212 ( .A(n307), .B(n308), .Y(SUM[2]) );
  NOR2XL U213 ( .A(n309), .B(n310), .Y(n308) );
  XNOR2X4 U214 ( .A(n325), .B(n414), .Y(SUM[26]) );
  AOI21X2 U215 ( .A0(n381), .A1(n426), .B0(n375), .Y(n380) );
  XOR2X2 U216 ( .A(n282), .B(n415), .Y(SUM[5]) );
  XNOR2X4 U217 ( .A(n416), .B(n312), .Y(SUM[29]) );
  XOR2X2 U218 ( .A(n366), .B(n417), .Y(SUM[17]) );
  OR2X4 U219 ( .A(n357), .B(n352), .Y(n417) );
  NAND2BX1 U220 ( .AN(n353), .B(n354), .Y(n365) );
  XNOR2XL U221 ( .A(n418), .B(n290), .Y(SUM[3]) );
  NAND2BXL U222 ( .AN(n360), .B(n361), .Y(n359) );
  XOR2X1 U223 ( .A(A[24]), .B(B[24]), .Y(n419) );
  XOR2XL U224 ( .A(n447), .B(B[23]), .Y(n340) );
  XOR2X1 U225 ( .A(B[19]), .B(A[19]), .Y(n363) );
  INVXL U226 ( .A(B[23]), .Y(n432) );
  NAND2XL U227 ( .A(B[0]), .B(A[0]), .Y(n358) );
  XOR2X1 U228 ( .A(B[7]), .B(A[7]), .Y(n276) );
  NOR2XL U229 ( .A(B[15]), .B(A[15]), .Y(n372) );
  NAND2XL U230 ( .A(B[16]), .B(A[16]), .Y(n368) );
  INVX1 U231 ( .A(A[23]), .Y(n447) );
  XOR2X4 U232 ( .A(n421), .B(n296), .Y(n420) );
  OAI21XL U233 ( .A0(B[0]), .A1(A[0]), .B0(n358), .Y(n408) );
  NAND2XL U234 ( .A(B[15]), .B(A[15]), .Y(n373) );
  BUFX8 U235 ( .A(n293), .Y(n421) );
  NAND2X1 U236 ( .A(B[1]), .B(A[1]), .Y(n361) );
  OAI31X4 U237 ( .A0(n370), .A1(n371), .A2(n372), .B0(n373), .Y(n356) );
  AOI21X2 U238 ( .A0(n374), .A1(n425), .B0(n375), .Y(n370) );
  INVX4 U239 ( .A(n401), .Y(n439) );
  CLKINVX4 U240 ( .A(n344), .Y(n429) );
  CLKINVX4 U241 ( .A(A[11]), .Y(n444) );
  CLKINVX4 U242 ( .A(A[3]), .Y(n448) );
endmodule


module hash_core_DW01_add_19 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n429, n270, n272, n273, n275, n276, n277, n278, n279, n280, n281,
         n282, n284, n285, n287, n288, n289, n290, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n381, n383, n384, n385, n386,
         n387, n388, n389, n390, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n271, n274, n283, n286, n291, n292, n380,
         n382, n391, n402, n403, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428;

  XOR2X4 U6 ( .A(n279), .B(n278), .Y(SUM[7]) );
  AOI2BB1X4 U11 ( .A0N(n424), .A1N(n284), .B0(n285), .Y(n280) );
  OAI2BB1X4 U14 ( .A0N(n289), .A1N(n288), .B0(n290), .Y(n284) );
  XNOR2X4 U23 ( .A(n303), .B(n302), .Y(SUM[30]) );
  OAI21X4 U24 ( .A0(n304), .A1(n428), .B0(n305), .Y(n302) );
  OAI2BB1X4 U25 ( .A0N(n428), .A1N(n304), .B0(B[29]), .Y(n305) );
  NOR2X4 U30 ( .A(n295), .B(n307), .Y(n306) );
  XOR2X4 U36 ( .A(n312), .B(n315), .Y(SUM[28]) );
  AND2X2 U38 ( .A(B[28]), .B(A[28]), .Y(n313) );
  OAI21X4 U40 ( .A0(n316), .A1(n317), .B0(n318), .Y(n312) );
  AOI21X4 U42 ( .A0(n320), .A1(n407), .B0(n321), .Y(n317) );
  XOR2X4 U46 ( .A(n320), .B(n323), .Y(SUM[26]) );
  AND2X2 U48 ( .A(B[26]), .B(A[26]), .Y(n321) );
  OAI21X4 U50 ( .A0(n324), .A1(n325), .B0(n326), .Y(n320) );
  XOR2X4 U51 ( .A(n327), .B(n324), .Y(SUM[25]) );
  XOR2X4 U56 ( .A(n328), .B(n331), .Y(SUM[24]) );
  AND2X2 U58 ( .A(B[24]), .B(A[24]), .Y(n329) );
  OAI21X4 U60 ( .A0(n332), .A1(n333), .B0(n334), .Y(n328) );
  XOR2X4 U61 ( .A(n335), .B(n333), .Y(SUM[23]) );
  XOR2X4 U66 ( .A(n336), .B(n339), .Y(SUM[22]) );
  AND2X2 U68 ( .A(B[22]), .B(A[22]), .Y(n337) );
  OAI21X4 U70 ( .A0(n340), .A1(n341), .B0(n342), .Y(n336) );
  XOR2X4 U76 ( .A(n344), .B(n347), .Y(SUM[20]) );
  OAI21X4 U80 ( .A0(n348), .A1(n349), .B0(n350), .Y(n344) );
  XOR2X4 U81 ( .A(n351), .B(n248), .Y(SUM[1]) );
  XOR2X4 U83 ( .A(n352), .B(n349), .Y(SUM[19]) );
  XOR2X4 U88 ( .A(n353), .B(n356), .Y(SUM[18]) );
  OAI21X4 U92 ( .A0(n357), .A1(n358), .B0(n359), .Y(n353) );
  XOR2X4 U98 ( .A(n361), .B(n364), .Y(SUM[16]) );
  AND2X2 U100 ( .A(B[16]), .B(A[16]), .Y(n362) );
  OAI2BB1X4 U105 ( .A0N(n426), .A1N(n365), .B0(B[15]), .Y(n366) );
  XOR2X4 U108 ( .A(n376), .B(n377), .Y(SUM[15]) );
  AND2X2 U113 ( .A(B[14]), .B(A[14]), .Y(n372) );
  NOR2X4 U120 ( .A(B[13]), .B(A[13]), .Y(n374) );
  NOR2X4 U124 ( .A(B[12]), .B(A[12]), .Y(n370) );
  OAI21X4 U132 ( .A0(n393), .A1(n387), .B0(n390), .Y(n392) );
  XOR2X4 U134 ( .A(n394), .B(n393), .Y(SUM[10]) );
  AOI2BB1X4 U135 ( .A0N(n270), .A1N(n273), .B0(n272), .Y(n393) );
  AOI21X4 U138 ( .A0(n275), .A1(n277), .B0(n418), .Y(n270) );
  NAND2X4 U139 ( .A(B[8]), .B(A[8]), .Y(n276) );
  OR2X4 U140 ( .A(B[8]), .B(A[8]), .Y(n277) );
  OAI21X4 U141 ( .A0(n395), .A1(n396), .B0(n397), .Y(n275) );
  OAI2BB1X4 U143 ( .A0N(n297), .A1N(n295), .B0(n399), .Y(n288) );
  NAND2X4 U148 ( .A(n250), .B(A[1]), .Y(n310) );
  NOR2X4 U149 ( .A(B[2]), .B(A[2]), .Y(n307) );
  OR2X4 U151 ( .A(A[3]), .B(B[3]), .Y(n297) );
  OR2X4 U152 ( .A(B[4]), .B(A[4]), .Y(n289) );
  NOR2X4 U153 ( .A(A[7]), .B(B[7]), .Y(n396) );
  AOI211X2 U154 ( .A0(B[7]), .A1(A[7]), .B0(n401), .C0(n281), .Y(n395) );
  AND2X2 U155 ( .A(B[6]), .B(A[6]), .Y(n281) );
  AOI21X4 U156 ( .A0(n253), .A1(n290), .B0(n422), .Y(n401) );
  NOR2X4 U158 ( .A(B[6]), .B(A[6]), .Y(n282) );
  NOR2X4 U159 ( .A(B[5]), .B(A[5]), .Y(n285) );
  NAND2X4 U160 ( .A(B[4]), .B(A[4]), .Y(n290) );
  NAND2X4 U2 ( .A(n283), .B(n375), .Y(n378) );
  OR2X4 U3 ( .A(n374), .B(n381), .Y(n283) );
  XNOR2X4 U4 ( .A(n280), .B(n246), .Y(SUM[6]) );
  OR2XL U5 ( .A(n281), .B(n282), .Y(n246) );
  NAND2X1 U7 ( .A(n288), .B(n258), .Y(n397) );
  OAI21X2 U8 ( .A0(A[11]), .A1(n388), .B0(B[11]), .Y(n384) );
  INVXL U9 ( .A(A[15]), .Y(n426) );
  NOR2X2 U10 ( .A(B[16]), .B(A[16]), .Y(n363) );
  INVXL U12 ( .A(n281), .Y(n251) );
  INVXL U13 ( .A(n282), .Y(n421) );
  NAND2BX1 U15 ( .AN(n358), .B(n359), .Y(n360) );
  INVX2 U16 ( .A(n263), .Y(SUM[8]) );
  AND2X2 U17 ( .A(n253), .B(n262), .Y(n286) );
  NAND2X2 U18 ( .A(n414), .B(n375), .Y(n292) );
  INVX1 U19 ( .A(n355), .Y(n411) );
  NOR2X1 U20 ( .A(n355), .B(n354), .Y(n356) );
  NOR2X2 U21 ( .A(n363), .B(n362), .Y(n364) );
  XOR2X2 U22 ( .A(n311), .B(n304), .Y(SUM[29]) );
  INVX1 U26 ( .A(B[4]), .Y(n249) );
  OAI211X4 U27 ( .A0(n365), .A1(n426), .B0(n366), .C0(n367), .Y(n361) );
  NAND2X2 U28 ( .A(n296), .B(n297), .Y(n247) );
  XOR2X4 U29 ( .A(n293), .B(n247), .Y(SUM[3]) );
  XNOR2X2 U31 ( .A(n275), .B(n264), .Y(n263) );
  OAI2BB1X4 U32 ( .A0N(n250), .A1N(A[1]), .B0(n256), .Y(n351) );
  NAND2X4 U33 ( .A(n254), .B(n266), .Y(n267) );
  INVX4 U34 ( .A(n265), .Y(n254) );
  AOI21X2 U35 ( .A0(n418), .A1(n419), .B0(n272), .Y(n389) );
  AND2X4 U37 ( .A(B[9]), .B(A[9]), .Y(n272) );
  AOI21X2 U39 ( .A0(n294), .A1(n423), .B0(n295), .Y(n293) );
  NAND2X1 U41 ( .A(A[0]), .B(B[0]), .Y(n248) );
  XNOR3X4 U43 ( .A(A[4]), .B(n249), .C(n288), .Y(n429) );
  BUFX16 U44 ( .A(B[1]), .Y(n250) );
  BUFX12 U45 ( .A(n429), .Y(SUM[4]) );
  XOR2X4 U47 ( .A(n294), .B(n306), .Y(SUM[2]) );
  XOR2X2 U49 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  OAI2BB2X4 U52 ( .B0(n308), .B1(n309), .A0N(n250), .A1N(A[1]), .Y(n294) );
  AOI31X2 U53 ( .A0(n400), .A1(n423), .A2(n297), .B0(n425), .Y(n399) );
  INVX4 U54 ( .A(n307), .Y(n423) );
  INVXL U55 ( .A(n296), .Y(n425) );
  OAI2BB1X4 U57 ( .A0N(n421), .A1N(n280), .B0(n251), .Y(n252) );
  INVX4 U59 ( .A(n252), .Y(n279) );
  BUFX8 U62 ( .A(n287), .Y(n253) );
  INVX1 U63 ( .A(n368), .Y(n265) );
  NAND2X1 U64 ( .A(n261), .B(n275), .Y(n385) );
  NAND3X1 U65 ( .A(n289), .B(n398), .C(n420), .Y(n257) );
  NOR2X4 U67 ( .A(n285), .B(n282), .Y(n398) );
  OAI2BB1X4 U69 ( .A0N(n289), .A1N(n288), .B0(n290), .Y(n255) );
  INVX4 U71 ( .A(n291), .Y(SUM[13]) );
  OR2X4 U72 ( .A(n250), .B(A[1]), .Y(n256) );
  NOR2X4 U73 ( .A(n250), .B(A[1]), .Y(n308) );
  NAND2X4 U74 ( .A(B[0]), .B(A[0]), .Y(n309) );
  INVX1 U75 ( .A(n257), .Y(n258) );
  INVX4 U77 ( .A(n396), .Y(n420) );
  NAND2X1 U78 ( .A(B[5]), .B(A[5]), .Y(n287) );
  NAND2X4 U79 ( .A(B[3]), .B(A[3]), .Y(n296) );
  XNOR2XL U82 ( .A(n292), .B(n381), .Y(n291) );
  AOI21X4 U84 ( .A0(n378), .A1(n413), .B0(n372), .Y(n377) );
  AOI2BB1XL U85 ( .A0N(A[11]), .A1N(B[11]), .B0(n387), .Y(n386) );
  NAND3XL U86 ( .A(n277), .B(n386), .C(n419), .Y(n260) );
  INVX2 U87 ( .A(n260), .Y(n261) );
  INVX4 U89 ( .A(n273), .Y(n419) );
  XNOR2X1 U90 ( .A(B[15]), .B(A[15]), .Y(n376) );
  NAND2X2 U91 ( .A(n274), .B(n390), .Y(n388) );
  INVX4 U93 ( .A(n387), .Y(n269) );
  INVX2 U94 ( .A(n389), .Y(n271) );
  INVXL U95 ( .A(n285), .Y(n262) );
  NOR2X1 U96 ( .A(n370), .B(n416), .Y(n383) );
  INVXL U97 ( .A(n253), .Y(n424) );
  INVX2 U99 ( .A(n388), .Y(n417) );
  NAND2X2 U101 ( .A(B[13]), .B(A[13]), .Y(n375) );
  NAND2X2 U102 ( .A(n265), .B(n383), .Y(n268) );
  NAND2X4 U103 ( .A(n267), .B(n268), .Y(SUM[12]) );
  AOI21X4 U104 ( .A0(n328), .A1(n408), .B0(n329), .Y(n324) );
  XOR2X2 U106 ( .A(n298), .B(n299), .Y(SUM[31]) );
  AND2X1 U107 ( .A(n276), .B(n277), .Y(n264) );
  AOI21X4 U109 ( .A0(n344), .A1(n410), .B0(n345), .Y(n340) );
  INVX4 U110 ( .A(n370), .Y(n415) );
  AOI21X4 U111 ( .A0(n368), .A1(n415), .B0(n416), .Y(n381) );
  NAND2X1 U112 ( .A(n269), .B(n271), .Y(n274) );
  OAI211X2 U114 ( .A0(n417), .A1(n427), .B0(n384), .C0(n385), .Y(n368) );
  AND2X1 U115 ( .A(B[20]), .B(A[20]), .Y(n345) );
  INVX1 U116 ( .A(n383), .Y(n266) );
  NOR2X2 U117 ( .A(B[10]), .B(A[10]), .Y(n387) );
  XOR2X4 U118 ( .A(n360), .B(n357), .Y(SUM[17]) );
  INVX1 U119 ( .A(n319), .Y(n382) );
  NAND2X4 U121 ( .A(B[10]), .B(A[10]), .Y(n390) );
  XOR2X4 U122 ( .A(n255), .B(n286), .Y(SUM[5]) );
  XOR2X4 U123 ( .A(n270), .B(n402), .Y(SUM[9]) );
  OR2XL U125 ( .A(n272), .B(n273), .Y(n402) );
  XOR2X4 U126 ( .A(n378), .B(n380), .Y(SUM[14]) );
  NOR2X2 U127 ( .A(n379), .B(n372), .Y(n380) );
  AOI21X4 U128 ( .A0(n361), .A1(n412), .B0(n362), .Y(n357) );
  AOI21X4 U129 ( .A0(n353), .A1(n411), .B0(n354), .Y(n349) );
  AOI21X4 U130 ( .A0(n336), .A1(n409), .B0(n337), .Y(n333) );
  XNOR2X4 U131 ( .A(n382), .B(n317), .Y(SUM[27]) );
  NOR2X4 U133 ( .A(B[9]), .B(A[9]), .Y(n273) );
  XNOR2X4 U136 ( .A(n391), .B(n392), .Y(SUM[11]) );
  XNOR2XL U137 ( .A(B[11]), .B(A[11]), .Y(n391) );
  NAND2X4 U142 ( .A(B[12]), .B(A[12]), .Y(n373) );
  NOR2X4 U144 ( .A(A[14]), .B(B[14]), .Y(n379) );
  AND2X1 U145 ( .A(B[18]), .B(A[18]), .Y(n354) );
  NAND2BXL U146 ( .AN(n387), .B(n390), .Y(n394) );
  INVX1 U147 ( .A(n363), .Y(n412) );
  INVX1 U150 ( .A(n346), .Y(n410) );
  INVX1 U157 ( .A(n338), .Y(n409) );
  XOR2X2 U161 ( .A(n343), .B(n340), .Y(SUM[21]) );
  NAND2BX1 U162 ( .AN(n341), .B(n342), .Y(n343) );
  NAND2BX1 U163 ( .AN(n348), .B(n350), .Y(n352) );
  NAND2BX1 U164 ( .AN(n332), .B(n334), .Y(n335) );
  NOR2X1 U165 ( .A(n346), .B(n345), .Y(n347) );
  NOR2X1 U166 ( .A(n330), .B(n329), .Y(n331) );
  NOR2X1 U167 ( .A(n338), .B(n337), .Y(n339) );
  AOI21X2 U168 ( .A0(n406), .A1(n312), .B0(n313), .Y(n304) );
  INVX1 U169 ( .A(n314), .Y(n406) );
  INVX1 U170 ( .A(n330), .Y(n408) );
  INVX1 U171 ( .A(n322), .Y(n407) );
  NAND2BX1 U172 ( .AN(n300), .B(n301), .Y(n303) );
  INVX1 U173 ( .A(n379), .Y(n413) );
  NAND2BX1 U174 ( .AN(n325), .B(n326), .Y(n327) );
  NAND2BX1 U175 ( .AN(n316), .B(n318), .Y(n319) );
  OAI21XL U176 ( .A0(n373), .A1(n374), .B0(n375), .Y(n371) );
  OAI21XL U177 ( .A0(n300), .A1(n405), .B0(n301), .Y(n298) );
  INVXL U178 ( .A(n302), .Y(n405) );
  NOR2X1 U179 ( .A(n314), .B(n313), .Y(n315) );
  NOR2X1 U180 ( .A(n322), .B(n321), .Y(n323) );
  INVX1 U181 ( .A(n373), .Y(n416) );
  INVXL U182 ( .A(A[11]), .Y(n427) );
  AOI21X2 U183 ( .A0(n413), .A1(n371), .B0(n372), .Y(n365) );
  NAND4XL U184 ( .A(n254), .B(n413), .C(n414), .D(n369), .Y(n367) );
  OAI2BB1X1 U185 ( .A0N(A[7]), .A1N(B[7]), .B0(n420), .Y(n278) );
  XNOR2X1 U186 ( .A(A[29]), .B(B[29]), .Y(n311) );
  NOR2X1 U187 ( .A(B[17]), .B(A[17]), .Y(n358) );
  NAND2X1 U188 ( .A(B[17]), .B(A[17]), .Y(n359) );
  AOI2BB1XL U189 ( .A0N(A[15]), .A1N(B[15]), .B0(n370), .Y(n369) );
  XOR2X1 U190 ( .A(B[31]), .B(A[31]), .Y(n299) );
  NOR2X1 U191 ( .A(B[18]), .B(A[18]), .Y(n355) );
  NOR2X1 U192 ( .A(B[20]), .B(A[20]), .Y(n346) );
  NOR2X1 U193 ( .A(B[19]), .B(A[19]), .Y(n348) );
  NAND2X1 U194 ( .A(B[19]), .B(A[19]), .Y(n350) );
  NOR2X1 U195 ( .A(A[22]), .B(B[22]), .Y(n338) );
  NOR2X1 U196 ( .A(B[23]), .B(A[23]), .Y(n332) );
  NOR2X1 U197 ( .A(B[21]), .B(A[21]), .Y(n341) );
  NAND2X1 U198 ( .A(B[21]), .B(A[21]), .Y(n342) );
  NAND2X1 U199 ( .A(B[23]), .B(A[23]), .Y(n334) );
  NOR2X1 U200 ( .A(A[26]), .B(B[26]), .Y(n322) );
  NOR2X1 U201 ( .A(B[24]), .B(A[24]), .Y(n330) );
  NOR2X1 U202 ( .A(B[25]), .B(A[25]), .Y(n325) );
  NAND2X1 U203 ( .A(B[25]), .B(A[25]), .Y(n326) );
  NOR2X1 U204 ( .A(B[28]), .B(A[28]), .Y(n314) );
  NOR2X1 U205 ( .A(B[27]), .B(A[27]), .Y(n316) );
  NAND2X1 U206 ( .A(B[27]), .B(A[27]), .Y(n318) );
  NOR2X1 U207 ( .A(B[30]), .B(A[30]), .Y(n300) );
  NAND2X1 U208 ( .A(B[30]), .B(A[30]), .Y(n301) );
  AOI2BB2X4 U209 ( .B0(n310), .B1(n403), .A0N(A[1]), .A1N(n250), .Y(n400) );
  NAND2X4 U210 ( .A(A[0]), .B(B[0]), .Y(n403) );
  AND2X4 U211 ( .A(B[2]), .B(A[2]), .Y(n295) );
  CLKINVX4 U212 ( .A(n374), .Y(n414) );
  CLKINVX4 U213 ( .A(n276), .Y(n418) );
  CLKINVX4 U214 ( .A(n398), .Y(n422) );
  CLKINVX4 U215 ( .A(A[29]), .Y(n428) );
endmodule


module hash_core_DW01_add_24 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n297,
         n298, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n333,
         n334, n335, n336, n337, n338, n339, n341, n342, n343, n344, n345,
         n346, n347, n349, n350, n351, n352, n353, n354, n355, n357, n358,
         n359, n360, n361, n362, n363, n365, n366, n367, n369, n370, n371,
         n372, n374, n375, n376, n377, n378, n379, n380, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n394, n395, n396,
         n397, n398, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n410, n411, n412, n414, n415, n416, n417, n418, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n296, n299, n312, n332, n340,
         n348, n356, n364, n368, n373, n381, n393, n399, n409, n413, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459;

  NAND3BX4 U11 ( .AN(n262), .B(n300), .C(n301), .Y(n293) );
  XOR2X4 U14 ( .A(n306), .B(n307), .Y(SUM[5]) );
  XOR2X4 U19 ( .A(n313), .B(n314), .Y(SUM[3]) );
  XNOR2X4 U26 ( .A(n322), .B(n320), .Y(SUM[30]) );
  OAI21X4 U27 ( .A0(n323), .A1(n447), .B0(n324), .Y(n320) );
  OAI2BB1X4 U28 ( .A0N(n447), .A1N(n323), .B0(B[29]), .Y(n324) );
  XOR2X4 U30 ( .A(n325), .B(n316), .Y(SUM[2]) );
  AOI21X4 U31 ( .A0(n450), .A1(n266), .B0(n326), .Y(n316) );
  AOI21X4 U35 ( .A0(n435), .A1(n329), .B0(n330), .Y(n323) );
  XNOR2X4 U36 ( .A(A[29]), .B(B[29]), .Y(n328) );
  AND2X2 U39 ( .A(B[28]), .B(A[28]), .Y(n330) );
  OAI21X4 U41 ( .A0(n333), .A1(n334), .B0(n335), .Y(n329) );
  AOI21X4 U43 ( .A0(n337), .A1(n434), .B0(n338), .Y(n334) );
  AND2X2 U49 ( .A(B[26]), .B(A[26]), .Y(n338) );
  OAI21X4 U51 ( .A0(n341), .A1(n342), .B0(n343), .Y(n337) );
  AOI21X4 U53 ( .A0(n345), .A1(n436), .B0(n346), .Y(n341) );
  NOR2X4 U56 ( .A(B[25]), .B(A[25]), .Y(n342) );
  AND2X2 U59 ( .A(B[24]), .B(A[24]), .Y(n346) );
  XOR2X4 U62 ( .A(n352), .B(n350), .Y(SUM[23]) );
  AOI21X4 U63 ( .A0(n353), .A1(n437), .B0(n354), .Y(n350) );
  NAND2BX4 U64 ( .AN(n349), .B(n351), .Y(n352) );
  NOR2X4 U66 ( .A(B[23]), .B(A[23]), .Y(n349) );
  AND2X2 U69 ( .A(B[22]), .B(A[22]), .Y(n354) );
  OAI21X4 U71 ( .A0(n357), .A1(n358), .B0(n359), .Y(n353) );
  XOR2X4 U72 ( .A(n360), .B(n357), .Y(SUM[21]) );
  AOI21X4 U73 ( .A0(n361), .A1(n438), .B0(n362), .Y(n357) );
  AND2X2 U79 ( .A(B[20]), .B(A[20]), .Y(n362) );
  OAI21X4 U81 ( .A0(n365), .A1(n366), .B0(n367), .Y(n361) );
  NOR2X4 U88 ( .A(B[19]), .B(A[19]), .Y(n365) );
  AND2X2 U91 ( .A(B[18]), .B(A[18]), .Y(n371) );
  AND2X2 U101 ( .A(B[16]), .B(A[16]), .Y(n379) );
  OAI211X2 U103 ( .A0(n382), .A1(n445), .B0(n383), .C0(n384), .Y(n378) );
  AOI2BB1X4 U105 ( .A0N(A[15]), .A1N(B[15]), .B0(n388), .Y(n387) );
  AOI21X4 U107 ( .A0(n386), .A1(n389), .B0(n448), .Y(n382) );
  XNOR2X4 U112 ( .A(n397), .B(n395), .Y(SUM[14]) );
  OAI21X4 U113 ( .A0(n391), .A1(n398), .B0(n392), .Y(n395) );
  AOI21X4 U118 ( .A0(n385), .A1(n443), .B0(n442), .Y(n398) );
  AOI21X4 U127 ( .A0(n444), .A1(n406), .B0(n407), .Y(n401) );
  AOI21X4 U133 ( .A0(n411), .A1(n444), .B0(n407), .Y(n410) );
  NOR2X4 U138 ( .A(B[10]), .B(A[10]), .Y(n412) );
  OAI21X4 U139 ( .A0(n286), .A1(n405), .B0(n287), .Y(n411) );
  AOI21X4 U142 ( .A0(n288), .A1(n451), .B0(n296), .Y(n286) );
  OR2X4 U145 ( .A(B[7]), .B(A[7]), .Y(n294) );
  NAND2X4 U147 ( .A(A[6]), .B(B[6]), .Y(n298) );
  NAND2X4 U148 ( .A(A[7]), .B(B[7]), .Y(n295) );
  NAND2X4 U152 ( .A(n258), .B(n304), .Y(n310) );
  OR2X4 U153 ( .A(B[3]), .B(A[3]), .Y(n303) );
  NAND3BX4 U154 ( .AN(n417), .B(n279), .C(n418), .Y(n304) );
  NOR2X4 U158 ( .A(B[2]), .B(A[2]), .Y(n315) );
  NOR2X4 U159 ( .A(B[4]), .B(A[4]), .Y(n309) );
  NOR2X4 U161 ( .A(B[6]), .B(A[6]), .Y(n297) );
  AOI2BB1X4 U166 ( .A0N(n265), .A1N(A[0]), .B0(n450), .Y(SUM[0]) );
  NAND2X4 U167 ( .A(A[0]), .B(B[0]), .Y(n327) );
  INVXL U2 ( .A(n457), .Y(n285) );
  NAND3X4 U3 ( .A(n269), .B(n270), .C(n271), .Y(n255) );
  XNOR2X4 U4 ( .A(n400), .B(n255), .Y(SUM[12]) );
  OAI21X1 U5 ( .A0(B[11]), .A1(A[11]), .B0(n288), .Y(n404) );
  INVX8 U6 ( .A(n273), .Y(n288) );
  OAI2BB1X4 U7 ( .A0N(n445), .A1N(n382), .B0(B[15]), .Y(n383) );
  INVX8 U8 ( .A(n298), .Y(n456) );
  INVX8 U9 ( .A(n405), .Y(n299) );
  INVX1 U10 ( .A(n374), .Y(n340) );
  INVX2 U12 ( .A(n396), .Y(n448) );
  INVX1 U13 ( .A(n459), .Y(n263) );
  NAND2X2 U15 ( .A(n390), .B(n443), .Y(n400) );
  XNOR2X2 U16 ( .A(A[30]), .B(B[30]), .Y(n322) );
  NAND2BX2 U17 ( .AN(n365), .B(n367), .Y(n369) );
  XOR2X2 U18 ( .A(n328), .B(n323), .Y(SUM[29]) );
  INVX4 U20 ( .A(n377), .Y(n332) );
  NAND2X2 U21 ( .A(n377), .B(n340), .Y(n348) );
  NAND2BX4 U22 ( .AN(n375), .B(n376), .Y(n377) );
  INVX4 U23 ( .A(n456), .Y(n256) );
  XNOR2X4 U24 ( .A(n410), .B(n257), .Y(SUM[11]) );
  XOR2X1 U25 ( .A(B[11]), .B(A[11]), .Y(n257) );
  CLKINVX3 U29 ( .A(n264), .Y(n265) );
  CLKINVX2 U32 ( .A(B[0]), .Y(n264) );
  XOR2X4 U33 ( .A(n288), .B(n289), .Y(SUM[8]) );
  CLKBUFX2 U34 ( .A(n303), .Y(n258) );
  NAND3X2 U37 ( .A(n283), .B(n266), .C(n285), .Y(n418) );
  INVX1 U38 ( .A(n305), .Y(n427) );
  INVX8 U40 ( .A(n450), .Y(n259) );
  CLKINVX8 U42 ( .A(n327), .Y(n450) );
  BUFX2 U44 ( .A(n283), .Y(n260) );
  INVX8 U45 ( .A(n412), .Y(n444) );
  AOI21X4 U46 ( .A0(n395), .A1(n386), .B0(n448), .Y(n394) );
  NAND3BX4 U47 ( .AN(n278), .B(n453), .C(n302), .Y(n261) );
  OR2X4 U48 ( .A(n304), .B(n427), .Y(n302) );
  AND3X4 U50 ( .A(n263), .B(B[4]), .C(n454), .Y(n262) );
  NAND2X2 U52 ( .A(n454), .B(n453), .Y(n280) );
  NAND2X2 U54 ( .A(n310), .B(n305), .Y(n311) );
  NAND2X2 U55 ( .A(n428), .B(n292), .Y(n431) );
  INVX3 U57 ( .A(n292), .Y(n429) );
  NAND3BX2 U58 ( .AN(n262), .B(n261), .C(n301), .Y(n267) );
  INVX4 U60 ( .A(n458), .Y(n266) );
  CLKINVX8 U61 ( .A(A[1]), .Y(n458) );
  NOR2X2 U65 ( .A(n412), .B(n407), .Y(n422) );
  INVX4 U67 ( .A(n388), .Y(n443) );
  OAI2BB1X4 U68 ( .A0N(n268), .A1N(n301), .B0(n455), .Y(n415) );
  NAND3X1 U70 ( .A(A[4]), .B(B[4]), .C(n454), .Y(n268) );
  NAND3BX4 U74 ( .AN(n280), .B(n311), .C(n455), .Y(n416) );
  INVX2 U75 ( .A(n316), .Y(n282) );
  OR2X4 U76 ( .A(n401), .B(n446), .Y(n269) );
  OR2X4 U77 ( .A(n402), .B(n449), .Y(n270) );
  OR2X4 U78 ( .A(n403), .B(n404), .Y(n271) );
  NAND3X4 U80 ( .A(n269), .B(n270), .C(n271), .Y(n385) );
  INVXL U82 ( .A(A[11]), .Y(n446) );
  AND2X2 U83 ( .A(n401), .B(n446), .Y(n402) );
  INVXL U84 ( .A(B[11]), .Y(n449) );
  BUFX8 U85 ( .A(n317), .Y(n279) );
  INVX4 U86 ( .A(n277), .Y(n301) );
  NAND2X4 U87 ( .A(n284), .B(n279), .Y(n313) );
  NAND2X4 U89 ( .A(n260), .B(n282), .Y(n284) );
  XNOR2X4 U90 ( .A(n293), .B(n272), .Y(n421) );
  NOR2X4 U92 ( .A(n456), .B(n297), .Y(n272) );
  INVX4 U93 ( .A(A[4]), .Y(n459) );
  OAI2BB1X4 U94 ( .A0N(n274), .A1N(n275), .B0(n454), .Y(n278) );
  NAND2X4 U95 ( .A(n414), .B(n294), .Y(n273) );
  INVXL U96 ( .A(B[3]), .Y(n274) );
  INVXL U97 ( .A(A[3]), .Y(n275) );
  NAND2BX2 U98 ( .AN(n277), .B(n454), .Y(n381) );
  XNOR2X2 U99 ( .A(n369), .B(n366), .Y(n276) );
  CLKINVX8 U100 ( .A(n276), .Y(SUM[19]) );
  AOI21X4 U102 ( .A0(n458), .A1(n327), .B0(n457), .Y(n326) );
  AOI21X4 U104 ( .A0(n451), .A1(n288), .B0(n296), .Y(n281) );
  INVX4 U106 ( .A(n290), .Y(n451) );
  INVX8 U108 ( .A(n408), .Y(n296) );
  AOI211X2 U109 ( .A0(n458), .A1(n457), .B0(n315), .C0(n259), .Y(n417) );
  XOR2X4 U110 ( .A(n378), .B(n424), .Y(SUM[16]) );
  CLKINVX4 U111 ( .A(n381), .Y(n307) );
  INVX3 U114 ( .A(B[4]), .Y(n452) );
  NAND2X1 U115 ( .A(B[4]), .B(A[4]), .Y(n364) );
  INVX4 U116 ( .A(n291), .Y(n428) );
  NAND2X4 U117 ( .A(n294), .B(n295), .Y(n291) );
  AND2X4 U119 ( .A(B[5]), .B(A[5]), .Y(n277) );
  NAND3BX4 U120 ( .AN(n278), .B(n453), .C(n302), .Y(n300) );
  XNOR2X4 U121 ( .A(n311), .B(n368), .Y(SUM[4]) );
  NAND2X4 U122 ( .A(n364), .B(n453), .Y(n368) );
  INVX8 U123 ( .A(n308), .Y(n454) );
  XOR2X4 U124 ( .A(n457), .B(n433), .Y(n432) );
  INVX8 U125 ( .A(n315), .Y(n283) );
  NAND2X4 U126 ( .A(B[13]), .B(A[13]), .Y(n392) );
  NAND4X4 U128 ( .A(n416), .B(n415), .C(n295), .D(n256), .Y(n414) );
  OAI222X2 U129 ( .A0(n459), .A1(n452), .B0(n309), .B1(n305), .C0(n310), .C1(
        n309), .Y(n306) );
  NAND2X4 U130 ( .A(n291), .B(n429), .Y(n430) );
  AND2X4 U131 ( .A(n303), .B(n305), .Y(n314) );
  INVX8 U132 ( .A(n421), .Y(SUM[6]) );
  NAND2X4 U134 ( .A(n348), .B(n356), .Y(SUM[17]) );
  BUFX8 U135 ( .A(A[1]), .Y(n433) );
  NAND4X1 U136 ( .A(n255), .B(n386), .C(n441), .D(n387), .Y(n384) );
  NAND2X2 U137 ( .A(n441), .B(n392), .Y(n399) );
  INVX3 U140 ( .A(n391), .Y(n441) );
  INVX4 U141 ( .A(n309), .Y(n453) );
  XOR2X4 U143 ( .A(n259), .B(n432), .Y(SUM[1]) );
  XOR2X4 U144 ( .A(n281), .B(n393), .Y(SUM[9]) );
  NAND2X2 U146 ( .A(n296), .B(n299), .Y(n312) );
  NAND2X2 U149 ( .A(n312), .B(n287), .Y(n406) );
  NAND2X2 U150 ( .A(B[9]), .B(A[9]), .Y(n287) );
  NAND2XL U151 ( .A(n332), .B(n374), .Y(n356) );
  OAI21X4 U155 ( .A0(n390), .A1(n391), .B0(n392), .Y(n389) );
  NOR2X4 U156 ( .A(B[21]), .B(A[21]), .Y(n358) );
  NAND2XL U157 ( .A(B[21]), .B(A[21]), .Y(n359) );
  NOR2X4 U160 ( .A(B[5]), .B(A[5]), .Y(n308) );
  AOI21X4 U162 ( .A0(n370), .A1(n439), .B0(n371), .Y(n366) );
  NAND2X4 U163 ( .A(n373), .B(n376), .Y(n370) );
  XOR2X1 U164 ( .A(n370), .B(n419), .Y(SUM[18]) );
  NOR2X4 U165 ( .A(B[16]), .B(A[16]), .Y(n380) );
  AOI21X4 U168 ( .A0(n378), .A1(n440), .B0(n379), .Y(n374) );
  NAND2X4 U169 ( .A(B[12]), .B(A[12]), .Y(n390) );
  OR2X2 U170 ( .A(n374), .B(n375), .Y(n373) );
  NOR2X4 U171 ( .A(B[17]), .B(A[17]), .Y(n375) );
  NAND2X4 U172 ( .A(B[17]), .B(A[17]), .Y(n376) );
  NOR2X4 U173 ( .A(B[9]), .B(A[9]), .Y(n405) );
  OR2X4 U174 ( .A(A[14]), .B(B[14]), .Y(n386) );
  XOR2X2 U175 ( .A(n337), .B(n423), .Y(SUM[26]) );
  NOR2X2 U176 ( .A(B[8]), .B(A[8]), .Y(n290) );
  NOR2X2 U177 ( .A(B[24]), .B(A[24]), .Y(n347) );
  NAND2X2 U178 ( .A(n299), .B(n287), .Y(n393) );
  NOR2X4 U179 ( .A(B[13]), .B(A[13]), .Y(n391) );
  NOR2X4 U180 ( .A(B[20]), .B(A[20]), .Y(n363) );
  NAND2X4 U181 ( .A(B[25]), .B(A[25]), .Y(n343) );
  NOR2X4 U182 ( .A(B[12]), .B(A[12]), .Y(n388) );
  XOR2X4 U183 ( .A(n361), .B(n409), .Y(SUM[20]) );
  NOR2X4 U184 ( .A(n363), .B(n362), .Y(n409) );
  XOR2X4 U185 ( .A(n345), .B(n413), .Y(SUM[24]) );
  NOR2X4 U186 ( .A(n347), .B(n346), .Y(n413) );
  NAND2X2 U187 ( .A(B[8]), .B(A[8]), .Y(n408) );
  AOI21X4 U188 ( .A0(n320), .A1(A[30]), .B0(B[30]), .Y(n321) );
  NAND2X2 U189 ( .A(B[19]), .B(A[19]), .Y(n367) );
  NOR2X1 U190 ( .A(A[22]), .B(B[22]), .Y(n355) );
  XOR2X4 U191 ( .A(n344), .B(n341), .Y(SUM[25]) );
  NAND2BX4 U192 ( .AN(n342), .B(n343), .Y(n344) );
  OAI21X4 U193 ( .A0(n349), .A1(n350), .B0(n351), .Y(n345) );
  AOI21X4 U194 ( .A0(n267), .A1(n455), .B0(n456), .Y(n292) );
  XOR2X4 U195 ( .A(n398), .B(n399), .Y(SUM[13]) );
  NOR2XL U196 ( .A(n372), .B(n371), .Y(n419) );
  XOR2X1 U197 ( .A(n353), .B(n420), .Y(SUM[22]) );
  NOR2XL U198 ( .A(n355), .B(n354), .Y(n420) );
  XOR2X4 U199 ( .A(n411), .B(n422), .Y(SUM[10]) );
  INVXL U200 ( .A(n331), .Y(n435) );
  INVX4 U201 ( .A(n339), .Y(n434) );
  NOR2X4 U202 ( .A(n339), .B(n338), .Y(n423) );
  NAND2X4 U203 ( .A(A[3]), .B(B[3]), .Y(n305) );
  NAND2X4 U204 ( .A(B[14]), .B(A[14]), .Y(n396) );
  NOR2X2 U205 ( .A(n380), .B(n379), .Y(n424) );
  INVXL U206 ( .A(n390), .Y(n442) );
  NOR2X4 U207 ( .A(B[18]), .B(A[18]), .Y(n372) );
  INVXL U208 ( .A(A[15]), .Y(n445) );
  XNOR2X2 U209 ( .A(n318), .B(n319), .Y(SUM[31]) );
  NOR2X1 U210 ( .A(n296), .B(n290), .Y(n289) );
  NAND2X1 U211 ( .A(n396), .B(n386), .Y(n397) );
  INVX1 U212 ( .A(n363), .Y(n438) );
  INVX1 U213 ( .A(n347), .Y(n436) );
  INVX1 U214 ( .A(n372), .Y(n439) );
  INVX1 U215 ( .A(n355), .Y(n437) );
  NAND2BX1 U216 ( .AN(n358), .B(n359), .Y(n360) );
  XOR2X2 U217 ( .A(n336), .B(n334), .Y(SUM[27]) );
  NAND2BX1 U218 ( .AN(n333), .B(n335), .Y(n336) );
  XNOR2X4 U219 ( .A(n329), .B(n425), .Y(SUM[28]) );
  OR2X4 U220 ( .A(n331), .B(n330), .Y(n425) );
  INVX1 U221 ( .A(n380), .Y(n440) );
  NOR2X2 U222 ( .A(A[26]), .B(B[26]), .Y(n339) );
  NOR2X2 U223 ( .A(B[28]), .B(A[28]), .Y(n331) );
  NOR2X1 U224 ( .A(B[27]), .B(A[27]), .Y(n333) );
  NAND2X1 U225 ( .A(B[27]), .B(A[27]), .Y(n335) );
  NAND2X2 U226 ( .A(B[23]), .B(A[23]), .Y(n351) );
  AOI2BB1XL U227 ( .A0N(A[30]), .A1N(n320), .B0(n321), .Y(n318) );
  NAND3XL U228 ( .A(n299), .B(n451), .C(n444), .Y(n403) );
  XNOR2X4 U229 ( .A(n426), .B(n394), .Y(SUM[15]) );
  XOR2X1 U230 ( .A(B[15]), .B(A[15]), .Y(n426) );
  INVX1 U231 ( .A(A[29]), .Y(n447) );
  XNOR2X2 U232 ( .A(B[31]), .B(A[31]), .Y(n319) );
  NAND2X4 U233 ( .A(n430), .B(n431), .Y(SUM[7]) );
  NAND2X4 U234 ( .A(n283), .B(n317), .Y(n325) );
  NAND2X2 U235 ( .A(B[2]), .B(A[2]), .Y(n317) );
  AND2X4 U236 ( .A(B[10]), .B(A[10]), .Y(n407) );
  INVX8 U237 ( .A(n297), .Y(n455) );
  INVX8 U238 ( .A(B[1]), .Y(n457) );
endmodule


module hash_core ( clk, reset, Wt, inner_busy, first_block, output_enable, 
        digest );
  input [31:0] Wt;
  output [31:0] digest;
  input clk, reset, inner_busy, first_block, output_enable;
  wire   N121, N122, N123, N124, N125, N126, N127, N795, N796, N797, N798,
         N799, N800, N801, N802, N803, N804, N805, N806, N807, N808, N809,
         N810, N811, N812, N813, N814, N815, N816, N817, N818, N819, N820,
         N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831,
         N832, N833, N834, N835, N836, N837, N838, N839, N840, N841, N842,
         N843, N844, N845, N846, N847, N848, N849, N850, N851, N852, N853,
         N854, N855, N856, N857, N858, N859, N860, N861, N862, N863, N864,
         N865, N866, N867, N868, N869, N870, N871, N872, N873, N874, N875,
         N876, N877, N878, N879, N880, N881, N882, N883, N884, N885, N886,
         N887, N888, N889, N890, N891, N892, N893, N894, N895, N896, N897,
         N898, N899, N900, N901, N902, N903, N904, N905, N906, N907, N908,
         N909, N910, N911, N912, N913, N914, N915, N916, N917, N918, N919,
         N920, N921, N922, N923, N924, N925, N926, N927, N928, N929, N930,
         N931, N932, N933, N934, N935, N936, N937, N938, N939, N940, N941,
         N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952,
         N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963,
         N964, N965, N966, N967, N968, N969, N970, N971, N972, N973, N974,
         N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985,
         N986, N987, N988, N989, N990, N991, N992, N993, N994, N995, N996,
         N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006,
         N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016,
         N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026,
         N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036,
         N1037, N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046,
         N1047, N1048, N1049, N1050, N2946, N2947, N2948, N2949, N2950, N2951,
         N2952, N2953, N2954, N2955, N2956, N2957, N2958, N2959, N2960, N2961,
         N2962, N2963, N2964, N2965, N2966, N2967, N2968, N2969, N2970, N2971,
         N2972, N2973, N2974, N2975, N2976, N2977, N3047, N3048, N3049, N3050,
         N3051, N3052, N3053, N3054, N3055, N3056, N3057, N3058, N3059, N3060,
         N3061, N3062, N3063, N3064, N3065, N3066, N3067, N3068, N3069, N3070,
         N3071, N3072, N3073, N3074, N3075, N3076, N3077, N3078, N3079, N3080,
         N3081, n1140, n1141, n1142, n1143, n1144, n1145, n1151, n1152, n1153,
         n1154, n1156, n1157, n1161, n1163, n1165, n1167, n1168, n1434, n2417,
         n2419, n2420, n2422, n2423, n2424, n2425, n2426, n2432, n2433, n2436,
         n2437, n2439, n2443, n2444, n2447, n2449, n2451, n2452, n2454, n2455,
         n2456, n2457, n2458, n2464, n2465, n2468, n2469, n2471, n2475, n2476,
         n2479, n2483, n2484, n2485, n2486, n2487, n2488, n2494, n2495, n2496,
         n2497, n2499, n2500, n2503, n2504, n2506, n2508, n2510, n2514, n2515,
         n2516, n2517, n2518, n2519, n2525, n2526, n2527, n2528, n2530, n2531,
         n2534, n2535, n2537, n2539, n2541, n2542, n2543, n2546, n2547, n2548,
         n2549, n2553, n2554, n2556, n2557, n2558, n2560, n2561, n2562, n2563,
         n2566, n2567, n2569, n2570, n2571, n2574, n2575, n2577, n2580, n2582,
         n2584, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2596,
         n2598, n2601, n2602, n2603, n2605, n2608, n2610, n2614, n2619, n2620,
         n2621, n2624, n2626, n2629, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2642, n2643, n2645, n2646, n2652, n2654, n2656, n2657,
         n2659, n2663, n2667, n2668, n2671, n2674, n2675, n2677, n2678, n2684,
         n2686, n2688, n2689, n2691, n2695, n2699, n2700, n2704, n2706, n2710,
         n2715, n2716, n2717, n2720, n2722, n2725, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2737, n2740, n2742, n2744, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2756, n2758, n2761, n2762,
         n2763, n2765, n2769, n2770, n2771, n2772, n2776, n2777, n2779, n2780,
         n2781, n2783, n2784, n2785, n2786, n2789, n2790, n2792, n2793, n2794,
         n2797, n2800, n2802, n2803, n2804, n2806, n2807, n2809, n2810, n2813,
         n2814, n2815, n2816, n2818, n2820, n2821, n2822, n2824, n2829, n2831,
         n2832, n2834, n2835, n2836, n2838, n2839, n2841, n2842, n2845, n2846,
         n2847, n2848, n2850, n2852, n2853, n2854, n2856, n2861, n2863, n2865,
         n2866, n2868, n2870, n2876, n2879, n2880, n2881, n2882, n2885, n2886,
         n2889, n2890, n2893, n2894, n2895, n2897, n2898, n2900, n2902, n2908,
         n2911, n2912, n2913, n2914, n2917, n2918, n2921, n2922, n2925, n2926,
         n2927, n40, n259, n321, n353, n995, n996, n1048, n1049, n1050,
         T2_32_9_, T2_32_8_, T2_32_7_, T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_,
         T2_32_31_, T2_32_30_, T2_32_2_, T2_32_29_, T2_32_28_, T2_32_27_,
         T2_32_26_, T2_32_25_, T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_,
         T2_32_20_, T2_32_1_, T2_32_19_, T2_32_18_, T2_32_17_, T2_32_16_,
         T2_32_15_, T2_32_14_, T2_32_13_, T2_32_12_, T2_32_11_, T2_32_10_,
         T2_32_0_, T1_32_9_, T1_32_8_, T1_32_7_, T1_32_6_, T1_32_5_, T1_32_4_,
         T1_32_3_, T1_32_31_, T1_32_30_, T1_32_2_, T1_32_29_, T1_32_28_,
         T1_32_27_, T1_32_26_, T1_32_25_, T1_32_24_, T1_32_23_, T1_32_22_,
         T1_32_21_, T1_32_20_, T1_32_1_, T1_32_19_, T1_32_18_, T1_32_17_,
         T1_32_16_, T1_32_15_, T1_32_14_, T1_32_13_, T1_32_12_, T1_32_11_,
         T1_32_10_, T1_32_0_, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90,
         N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76,
         N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62,
         N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48,
         N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34,
         N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N119, N118, N117,
         N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106,
         N105, N104, N103, N102, N101, N100, n265, n287, n330, n365, n418,
         n447, n450, n452, n453, n454, n466, n468, n469, n470, n473, n474,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n536, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n656, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n677, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n969, n970, n972, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1092, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1146, n1147, n1148, n1149, n1150, n1155, n1158, n1159, n1162,
         n1164, n1166, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1246, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1263, n1265, n1266, n1270, n1271, n1272, n1273, n1274,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2680, n2681, n2682, n2683, n2685, n2687,
         n2690, n2692, n2693, n2694, n2696, n2697, n2698, n2701, n2702, n2703,
         n2705, n2707, n2708, n2709, n2711, n2712, n2713, n2714, n2718, n2719,
         n2721, n2723, n2724, n2726, n2727, n2736, n2738, n2739, n2741, n2743,
         n2745, n2746, n2755, n2757, n2759, n2760, n2764, n2766, n2767, n2768,
         n2773, n2774, n2775, n2778, n2782, n2787, n2788, n2791, n2795, n2796,
         n2798, n2799, n2801, n2805, n2808, n2811, n2812, n2817, n2819, n2823,
         n2825, n2826, n2827, n2828, n2830, n2833, n2837, n2840, n2843, n2844,
         n2849, n2851, n2855, n2857, n2858, n2859, n2860, n2862, n2864, n2867,
         n2869, n2871, n2872, n2873, n2874, n2875, n2877, n2878, n2883, n2884,
         n2887, n2888, n2891, n2892, n2896, n2899, n2901, n2903, n2904, n2905,
         n2906, n2907, n2909, n2910, n2915, n2916, n2919, n2920, n2923, n2924,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860;
  wire   [31:0] f1_EFG_32;
  wire   [31:0] f2_ABC_32;
  wire   [31:0] f3_A_32;
  wire   [31:0] f4_E_32;
  wire   [31:0] Kt;
  wire   [31:0] next_E;
  wire   [31:0] next_A;
  wire   [255:0] SHA256_result;
  wire   [6:0] round;
  wire   [31:0] H0;
  wire   [31:0] H1;
  wire   [31:0] H2;
  wire   [31:0] H3;
  wire   [31:0] H4;
  wire   [31:0] H5;
  wire   [31:0] H6;
  wire   [31:0] H7;
  wire   [2:0] read_counter;

  CLKINVX8 U2005 ( .A(reset), .Y(n1434) );
  DFFHQX4 E_reg_0_ ( .D(n2734), .CK(clk), .Q(SHA256_result[96]) );
  DFFHQX4 B_reg_0_ ( .D(n2831), .CK(clk), .Q(SHA256_result[192]) );
  DFFHQX4 A_reg_0_ ( .D(n2895), .CK(clk), .Q(SHA256_result[224]) );
  DFFHQX4 C_reg_0_ ( .D(n1622), .CK(clk), .Q(SHA256_result[160]) );
  DFFHQX4 C_reg_1_ ( .D(n2797), .CK(clk), .Q(SHA256_result[161]) );
  DFFX4 F_reg_1_ ( .D(n1568), .CK(clk), .Q(SHA256_result[65]), .QN(n1167) );
  DFFHQX4 B_reg_1_ ( .D(n1582), .CK(clk), .Q(SHA256_result[193]) );
  DFFHQX4 D_reg_0_ ( .D(n1595), .CK(clk), .Q(SHA256_result[128]) );
  DFFHQX4 A_reg_4_ ( .D(n3584), .CK(clk), .Q(SHA256_result[228]) );
  DFFHQX4 A_reg_5_ ( .D(n2890), .CK(clk), .Q(SHA256_result[229]) );
  DFFHQX4 A_reg_6_ ( .D(n2889), .CK(clk), .Q(SHA256_result[230]) );
  DFFHQX4 A_reg_7_ ( .D(n3583), .CK(clk), .Q(SHA256_result[231]) );
  DFFHQX4 A_reg_8_ ( .D(n3582), .CK(clk), .Q(SHA256_result[232]) );
  DFFHQX4 A_reg_11_ ( .D(n3581), .CK(clk), .Q(SHA256_result[235]) );
  DFFHQX4 A_reg_17_ ( .D(n3579), .CK(clk), .Q(SHA256_result[241]) );
  DFFHQX4 A_reg_20_ ( .D(n3577), .CK(clk), .Q(SHA256_result[244]) );
  DFFHQX4 A_reg_26_ ( .D(n3572), .CK(clk), .Q(SHA256_result[250]) );
  DFFHQX4 E_reg_18_ ( .D(n2716), .CK(clk), .Q(SHA256_result[114]) );
  DFFHQX4 E_reg_21_ ( .D(n3561), .CK(clk), .Q(SHA256_result[117]) );
  DFFHQX4 E_reg_22_ ( .D(n3560), .CK(clk), .Q(SHA256_result[118]) );
  DFFHQX4 A_reg_9_ ( .D(n2886), .CK(clk), .Q(SHA256_result[233]) );
  DFFHQX4 A_reg_10_ ( .D(n2885), .CK(clk), .Q(SHA256_result[234]) );
  DFFX4 F_reg_12_ ( .D(n1561), .CK(clk), .Q(SHA256_result[76]), .QN(n1156) );
  DFFHQX4 Kt_reg_15_ ( .D(N2961), .CK(clk), .Q(Kt[15]) );
  DFFHQX4 Kt_reg_14_ ( .D(N2960), .CK(clk), .Q(Kt[14]) );
  DFFHQX4 Kt_reg_13_ ( .D(N2959), .CK(clk), .Q(Kt[13]) );
  DFFHQX4 Kt_reg_12_ ( .D(N2958), .CK(clk), .Q(Kt[12]) );
  DFFHQX4 Kt_reg_11_ ( .D(N2957), .CK(clk), .Q(Kt[11]) );
  DFFHQX4 Kt_reg_10_ ( .D(N2956), .CK(clk), .Q(Kt[10]) );
  DFFX4 F_reg_11_ ( .D(n2691), .CK(clk), .Q(SHA256_result[75]), .QN(n1157) );
  DFFHQX4 F_reg_9_ ( .D(n1563), .CK(clk), .Q(SHA256_result[73]) );
  DFFHQX4 F_reg_10_ ( .D(n1562), .CK(clk), .Q(SHA256_result[74]) );
  DFFHQX4 G_reg_9_ ( .D(n1632), .CK(clk), .Q(SHA256_result[41]) );
  DFFHQX4 G_reg_13_ ( .D(n1630), .CK(clk), .Q(SHA256_result[45]) );
  DFFHQX4 H_reg_9_ ( .D(n1605), .CK(clk), .Q(SHA256_result[9]) );
  DFFHQX4 G_reg_12_ ( .D(n2499), .CK(clk), .Q(SHA256_result[44]) );
  DFFHQX4 C_reg_7_ ( .D(n1619), .CK(clk), .Q(SHA256_result[167]) );
  DFFHQX4 G_reg_10_ ( .D(n1631), .CK(clk), .Q(SHA256_result[42]) );
  DFFHQX4 B_reg_3_ ( .D(n1581), .CK(clk), .Q(SHA256_result[195]) );
  DFFHQX4 C_reg_2_ ( .D(n1621), .CK(clk), .Q(SHA256_result[162]) );
  DFFHQX4 H_reg_10_ ( .D(n2469), .CK(clk), .Q(SHA256_result[10]) );
  DFFHQX4 B_reg_7_ ( .D(n2824), .CK(clk), .Q(SHA256_result[199]) );
  DFFHQX4 B_reg_4_ ( .D(n1580), .CK(clk), .Q(SHA256_result[196]) );
  DFFHQX4 B_reg_6_ ( .D(n1578), .CK(clk), .Q(SHA256_result[198]) );
  DFFHQX4 C_reg_3_ ( .D(n1620), .CK(clk), .Q(SHA256_result[163]) );
  DFFHQX4 C_reg_9_ ( .D(n2789), .CK(clk), .Q(SHA256_result[169]) );
  DFFHQX4 B_reg_13_ ( .D(n2818), .CK(clk), .Q(SHA256_result[205]) );
  DFFHQX4 C_reg_13_ ( .D(n2785), .CK(clk), .Q(SHA256_result[173]) );
  DFFHQX4 B_reg_8_ ( .D(n1577), .CK(clk), .Q(SHA256_result[200]) );
  DFFHQX4 C_reg_5_ ( .D(n2793), .CK(clk), .Q(SHA256_result[165]) );
  DFFHQX4 C_reg_8_ ( .D(n2790), .CK(clk), .Q(SHA256_result[168]) );
  DFFHQX4 G_reg_11_ ( .D(n2500), .CK(clk), .Q(SHA256_result[43]) );
  DFFHQX4 B_reg_5_ ( .D(n1579), .CK(clk), .Q(SHA256_result[197]) );
  DFFHQX4 B_reg_9_ ( .D(n2822), .CK(clk), .Q(SHA256_result[201]) );
  DFFHQX4 C_reg_4_ ( .D(n2794), .CK(clk), .Q(SHA256_result[164]) );
  DFFHQX4 Kt_reg_0_ ( .D(N2946), .CK(clk), .Q(Kt[0]) );
  DFFHQX4 A_reg_1_ ( .D(n2894), .CK(clk), .Q(SHA256_result[225]) );
  DFFHQX4 A_reg_3_ ( .D(n3585), .CK(clk), .Q(SHA256_result[227]) );
  DFFHQX4 A_reg_12_ ( .D(n3580), .CK(clk), .Q(SHA256_result[236]) );
  DFFHQX4 A_reg_18_ ( .D(n3578), .CK(clk), .Q(SHA256_result[242]) );
  DFFHQX4 A_reg_23_ ( .D(n3574), .CK(clk), .Q(SHA256_result[247]) );
  DFFHQX4 A_reg_22_ ( .D(n3575), .CK(clk), .Q(SHA256_result[246]) );
  DFFHQX4 E_reg_17_ ( .D(n2717), .CK(clk), .Q(SHA256_result[113]) );
  DFFHQX4 E_reg_20_ ( .D(n3562), .CK(clk), .Q(SHA256_result[116]) );
  DFFHQX4 A_reg_2_ ( .D(n2893), .CK(clk), .Q(SHA256_result[226]) );
  DFFHQX4 A_reg_24_ ( .D(n3573), .CK(clk), .Q(SHA256_result[248]) );
  DFFHQX4 E_reg_19_ ( .D(n2715), .CK(clk), .Q(SHA256_result[115]) );
  DFFHQX4 E_reg_25_ ( .D(n3558), .CK(clk), .Q(SHA256_result[121]) );
  DFFHQX4 E_reg_14_ ( .D(n2720), .CK(clk), .Q(SHA256_result[110]) );
  DFFHQX4 E_reg_26_ ( .D(n3557), .CK(clk), .Q(SHA256_result[122]) );
  DFFHQX4 E_reg_16_ ( .D(n3563), .CK(clk), .Q(SHA256_result[112]) );
  DFFHQX4 E_reg_28_ ( .D(n2706), .CK(clk), .Q(SHA256_result[124]) );
  DFFHQX4 E_reg_13_ ( .D(n3565), .CK(clk), .Q(SHA256_result[109]) );
  DFFHQX4 E_reg_15_ ( .D(n3564), .CK(clk), .Q(SHA256_result[111]) );
  DFFHQX4 E_reg_9_ ( .D(n2725), .CK(clk), .Q(SHA256_result[105]) );
  DFFHQX4 E_reg_8_ ( .D(n3568), .CK(clk), .Q(SHA256_result[104]) );
  DFFHQX4 E_reg_10_ ( .D(n3567), .CK(clk), .Q(SHA256_result[106]) );
  DFFHQX4 E_reg_27_ ( .D(n3556), .CK(clk), .Q(SHA256_result[123]) );
  DFFHQX4 E_reg_12_ ( .D(n2722), .CK(clk), .Q(SHA256_result[108]) );
  DFFHQX4 E_reg_11_ ( .D(n3566), .CK(clk), .Q(SHA256_result[107]) );
  DFFX4 F_reg_0_ ( .D(n1569), .CK(clk), .Q(SHA256_result[64]), .QN(n1168) );
  DFFHQX4 Kt_reg_8_ ( .D(N2954), .CK(clk), .Q(Kt[8]) );
  DFFHQX4 Kt_reg_9_ ( .D(N2955), .CK(clk), .Q(Kt[9]) );
  DFFHQX4 Kt_reg_7_ ( .D(N2953), .CK(clk), .Q(Kt[7]) );
  DFFHQX4 Kt_reg_6_ ( .D(N2952), .CK(clk), .Q(Kt[6]) );
  DFFHQX4 Kt_reg_4_ ( .D(N2950), .CK(clk), .Q(Kt[4]) );
  DFFHQX4 Kt_reg_2_ ( .D(N2948), .CK(clk), .Q(Kt[2]) );
  DFFHQX4 Kt_reg_5_ ( .D(N2951), .CK(clk), .Q(Kt[5]) );
  DFFHQX4 H_reg_2_ ( .D(n1609), .CK(clk), .Q(SHA256_result[2]) );
  DFFHQX4 H_reg_6_ ( .D(n1607), .CK(clk), .Q(SHA256_result[6]) );
  DFFHQX4 H_reg_5_ ( .D(n1608), .CK(clk), .Q(SHA256_result[5]) );
  DFFHQX4 H_reg_1_ ( .D(n1610), .CK(clk), .Q(SHA256_result[1]) );
  DFFHQX4 F_reg_2_ ( .D(n2700), .CK(clk), .Q(SHA256_result[66]) );
  DFFHQX4 G_reg_7_ ( .D(n2504), .CK(clk), .Q(SHA256_result[39]) );
  DFFHQX4 H_reg_3_ ( .D(n2476), .CK(clk), .Q(SHA256_result[3]) );
  DFFHQX4 G_reg_8_ ( .D(n2503), .CK(clk), .Q(SHA256_result[40]) );
  DFFHQX4 H_reg_4_ ( .D(n2475), .CK(clk), .Q(SHA256_result[4]) );
  DFFHQX4 H_reg_0_ ( .D(n2479), .CK(clk), .Q(SHA256_result[0]) );
  DFFHQX4 H_reg_7_ ( .D(n1606), .CK(clk), .Q(SHA256_result[7]) );
  DFFHQX4 A_reg_25_ ( .D(n2870), .CK(clk), .Q(SHA256_result[249]) );
  DFFHQX4 A_reg_27_ ( .D(n2868), .CK(clk), .Q(SHA256_result[251]) );
  DFFHQX4 A_reg_14_ ( .D(n2881), .CK(clk), .Q(SHA256_result[238]) );
  DFFHQX4 A_reg_19_ ( .D(n2876), .CK(clk), .Q(SHA256_result[243]) );
  DFFHQX4 A_reg_15_ ( .D(n2880), .CK(clk), .Q(SHA256_result[239]) );
  DFFHQX4 A_reg_13_ ( .D(n2882), .CK(clk), .Q(SHA256_result[237]) );
  DFFHQX4 G_reg_3_ ( .D(n2508), .CK(clk), .Q(SHA256_result[35]) );
  DFFHQX4 E_reg_1_ ( .D(n2733), .CK(clk), .Q(SHA256_result[97]) );
  DFFHQX4 F_reg_6_ ( .D(n1565), .CK(clk), .Q(SHA256_result[70]) );
  DFFX4 F_reg_5_ ( .D(n1566), .CK(clk), .Q(SHA256_result[69]), .QN(n1163) );
  DFFHQX4 G_reg_6_ ( .D(n1633), .CK(clk), .Q(SHA256_result[38]) );
  DFFHQX4 F_reg_4_ ( .D(n1567), .CK(clk), .Q(SHA256_result[68]) );
  DFFHQX4 Kt_reg_1_ ( .D(N2947), .CK(clk), .Q(Kt[1]) );
  DFFHQX4 E_reg_2_ ( .D(n2732), .CK(clk), .Q(SHA256_result[98]) );
  DFFHQX4 E_reg_3_ ( .D(n2731), .CK(clk), .Q(SHA256_result[99]) );
  DFFHQX4 G_reg_5_ ( .D(n2506), .CK(clk), .Q(SHA256_result[37]) );
  DFFHQX4 A_reg_16_ ( .D(n2879), .CK(clk), .Q(SHA256_result[240]) );
  DFFHQX4 G_reg_4_ ( .D(n1634), .CK(clk), .Q(SHA256_result[36]) );
  DFFHQX4 Kt_reg_3_ ( .D(N2949), .CK(clk), .Q(Kt[3]) );
  DFFHQX4 E_reg_5_ ( .D(n2729), .CK(clk), .Q(SHA256_result[101]) );
  DFFHQX4 E_reg_4_ ( .D(n2730), .CK(clk), .Q(SHA256_result[100]) );
  DFFHQX4 G_reg_0_ ( .D(n2543), .CK(clk), .Q(SHA256_result[32]) );
  DFFHQX4 E_reg_6_ ( .D(n2728), .CK(clk), .Q(SHA256_result[102]) );
  DFFHQX4 E_reg_7_ ( .D(n3569), .CK(clk), .Q(SHA256_result[103]) );
  DFFHQX4 G_reg_1_ ( .D(n2510), .CK(clk), .Q(SHA256_result[33]) );
  DFFHQX4 C_reg_6_ ( .D(n2792), .CK(clk), .Q(SHA256_result[166]) );
  DFFHQX4 G_reg_2_ ( .D(n1635), .CK(clk), .Q(SHA256_result[34]) );
  DFFHQX4 B_reg_2_ ( .D(n2829), .CK(clk), .Q(SHA256_result[194]) );
  AND2X2 U879 ( .A(first_block), .B(n3013), .Y(n660) );
  AND2X2 U1288 ( .A(n1078), .B(n3724), .Y(n1237) );
  AND2X2 U1289 ( .A(output_enable), .B(n1434), .Y(n1078) );
  AND2X2 U1520 ( .A(n1399), .B(n3762), .Y(n1332) );
  hash_core_DW01_add_0 add_317 ( .A({SHA256_result[63:33], n2827}), .B(H7), 
        .SUM({N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, 
        N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, 
        N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, 
        N1021, N1020, N1019}) );
  hash_core_DW01_add_1 add_316 ( .A({SHA256_result[95:82], n3807, 
        SHA256_result[80], n3808, SHA256_result[78:64]}), .B(H6), .SUM({N1018, 
        N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, 
        N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, 
        N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987}) );
  hash_core_DW01_add_2 add_315 ( .A({n2682, n2871, n2860, n2874, n2864, n2877, 
        n2883, n2930, n2909, n2910, n2915, n2896, n2884, SHA256_result[114], 
        n2899, n2875, n2872, n2878, n2873, n2859, n2858, n2867, n2869, 
        SHA256_result[104], n2830, n2833, n2840, n2837, n2843, n2844, n2851, 
        n2934}), .B(H5), .SUM({N986, N985, N984, N983, N982, N981, N980, N979, 
        N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, 
        N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955}) );
  hash_core_DW01_add_4 add_313 ( .A(SHA256_result[191:160]), .B(H3), .SUM({
        N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, 
        N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, 
        N898, N897, N896, N895, N894, N893, N892, N891}) );
  hash_core_DW01_add_5 add_312 ( .A(SHA256_result[223:192]), .B(H2), .SUM({
        N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, 
        N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, 
        N866, N865, N864, N863, N862, N861, N860, N859}) );
  hash_core_DW01_add_6 add_311 ( .A({n2887, n2855, n2849, n2862, 
        SHA256_result[251], n2916, n2857, n2888, n2903, n2901, n2891, 
        SHA256_result[244:243], n2904, n2919, SHA256_result[240:234], n2907, 
        n2920, n2923, n2924, n2928, n2929, n2905, n2892, n2906, n2933}), .B(H1), .SUM({N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, 
        N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, 
        N834, N833, N832, N831, N830, N829, N828, N827}) );
  hash_core_DW01_inc_0 add_119 ( .A({round[6], n2932, round[4], n2931, n996, 
        round[1:0]}), .SUM({N127, N126, N125, N124, N123, N122, N121}) );
  hash_core_DW01_add_16 add_310 ( .A(next_A), .B(H0), .SUM({N826, N825, N824, 
        N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, 
        N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, 
        N799, N798, N797, N796, N795}) );
  hash_core_DW01_add_25 add_112 ( .A(SHA256_result[159:128]), .B({T1_32_31_, 
        T1_32_30_, T1_32_29_, T1_32_28_, n2694, T1_32_26_, T1_32_25_, 
        T1_32_24_, T1_32_23_, T1_32_22_, T1_32_21_, T1_32_20_, T1_32_19_, 
        T1_32_18_, T1_32_17_, T1_32_16_, T1_32_15_, T1_32_14_, T1_32_13_, 
        T1_32_12_, T1_32_11_, T1_32_10_, T1_32_9_, T1_32_8_, T1_32_7_, 
        T1_32_6_, T1_32_5_, T1_32_4_, T1_32_3_, T1_32_2_, T1_32_1_, T1_32_0_}), 
        .SUM(next_E) );
  hash_core_DW01_add_26 add_1_root_add_0_root_add_113 ( .A(f2_ABC_32), .B(
        f3_A_32), .SUM({T2_32_31_, T2_32_30_, T2_32_29_, T2_32_28_, T2_32_27_, 
        T2_32_26_, T2_32_25_, T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_, 
        T2_32_20_, T2_32_19_, T2_32_18_, T2_32_17_, T2_32_16_, T2_32_15_, 
        T2_32_14_, T2_32_13_, T2_32_12_, T2_32_11_, T2_32_10_, T2_32_9_, 
        T2_32_8_, T2_32_7_, T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_, T2_32_2_, 
        T2_32_1_, T2_32_0_}) );
  hash_core_DW01_add_27 add_0_root_add_0_root_add_108_4 ( .A({N119, N118, N117, 
        N116, N115, N114, N113, N112, N111, n2696, N109, N108, N107, N106, 
        N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, 
        N92, N91, N90, N89, N88}), .B({N87, N86, N85, N84, N83, N82, N81, N80, 
        N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, 
        N65, N64, N63, N62, N61, N60, N59, N58, N57, N56}), .SUM({T1_32_31_, 
        T1_32_30_, T1_32_29_, T1_32_28_, T1_32_27_, T1_32_26_, T1_32_25_, 
        T1_32_24_, T1_32_23_, T1_32_22_, T1_32_21_, T1_32_20_, T1_32_19_, 
        T1_32_18_, T1_32_17_, T1_32_16_, T1_32_15_, T1_32_14_, T1_32_13_, 
        T1_32_12_, T1_32_11_, T1_32_10_, T1_32_9_, T1_32_8_, T1_32_7_, 
        T1_32_6_, T1_32_5_, T1_32_4_, T1_32_3_, T1_32_2_, T1_32_1_, T1_32_0_})
         );
  hash_core_DW01_add_28 add_2_root_add_0_root_add_108_4 ( .A(
        SHA256_result[31:0]), .B({f1_EFG_32[31], n365, f1_EFG_32[29:23], n265, 
        n287, f1_EFG_32[20], n259, f1_EFG_32[18:11], n330, n321, 
        f1_EFG_32[8:7], n353, f1_EFG_32[5], n418, f1_EFG_32[3:0]}), .SUM({N119, 
        N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, 
        N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, 
        N93, N92, N91, N90, N89, N88}) );
  hash_core_DW01_add_7 add_314 ( .A({next_E[31], n2405, next_E[29], n2826, 
        next_E[27:0]}), .B(H4), .SUM({N954, N953, N952, N951, N950, N949, N948, 
        N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, 
        N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, 
        N923}) );
  hash_core_DW01_add_9 add_0_root_add_0_root_add_113 ( .A({T2_32_31_, 
        T2_32_30_, T2_32_29_, T2_32_28_, T2_32_27_, T2_32_26_, T2_32_25_, 
        T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_, T2_32_20_, T2_32_19_, 
        T2_32_18_, T2_32_17_, T2_32_16_, T2_32_15_, T2_32_14_, T2_32_13_, 
        T2_32_12_, T2_32_11_, T2_32_10_, T2_32_9_, T2_32_8_, T2_32_7_, 
        T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_, T2_32_2_, T2_32_1_, T2_32_0_}), 
        .B({T1_32_31_, T1_32_30_, T1_32_29_, T1_32_28_, T1_32_27_, T1_32_26_, 
        T1_32_25_, T1_32_24_, T1_32_23_, T1_32_22_, T1_32_21_, T1_32_20_, 
        T1_32_19_, T1_32_18_, T1_32_17_, n2693, T1_32_15_, n2701, T1_32_13_, 
        T1_32_12_, n2690, T1_32_10_, T1_32_9_, T1_32_8_, T1_32_7_, T1_32_6_, 
        T1_32_5_, T1_32_4_, T1_32_3_, n2697, T1_32_1_, T1_32_0_}), .SUM(next_A) );
  hash_core_DW01_add_19 add_3_root_add_0_root_add_108_4 ( .A(Wt), .B(Kt), 
        .SUM({N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24}) );
  hash_core_DW01_add_24 add_1_root_add_0_root_add_108_4 ( .A(f4_E_32), .B({N55, 
        N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, 
        N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24}), .SUM({N87, N86, N85, N84, N83, N82, N81, N80, N79, 
        N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, 
        N64, N63, N62, N61, N60, N59, N58, N57, N56}) );
  DFFHQXL A_reg_31_ ( .D(n3570), .CK(clk), .Q(SHA256_result[255]) );
  DFFHQX1 H0_reg_31_ ( .D(n3705), .CK(clk), .Q(H0[31]) );
  DFFHQXL H1_reg_31_ ( .D(n2832), .CK(clk), .Q(H1[31]) );
  DFFHQXL H5_reg_31_ ( .D(n2639), .CK(clk), .Q(H5[31]) );
  DFFHQX1 H2_reg_31_ ( .D(n3689), .CK(clk), .Q(H2[31]) );
  DFFHQX1 H6_reg_31_ ( .D(n3688), .CK(clk), .Q(H6[31]) );
  DFFHQXL H4_reg_30_ ( .D(n2608), .CK(clk), .Q(H4[30]) );
  DFFHQXL H7_reg_30_ ( .D(n2417), .CK(clk), .Q(H7[30]) );
  DFFHQXL H1_reg_27_ ( .D(n2836), .CK(clk), .Q(H1[27]) );
  DFFHQXL H1_reg_28_ ( .D(n2835), .CK(clk), .Q(H1[28]) );
  DFFHQXL H1_reg_29_ ( .D(n2834), .CK(clk), .Q(H1[29]) );
  DFFHQXL H2_reg_28_ ( .D(n2547), .CK(clk), .Q(H2[28]) );
  DFFHQXL H2_reg_29_ ( .D(n2546), .CK(clk), .Q(H2[29]) );
  DFFHQXL H5_reg_28_ ( .D(n2642), .CK(clk), .Q(H5[28]) );
  DFFHQXL H7_reg_27_ ( .D(n2420), .CK(clk), .Q(H7[27]) );
  DFFHQXL H7_reg_28_ ( .D(n2419), .CK(clk), .Q(H7[28]) );
  DFFHQX1 read_counter_reg_1_ ( .D(N3080), .CK(clk), .Q(read_counter[1]) );
  DFFHQX1 H6_reg_30_ ( .D(n3695), .CK(clk), .Q(H6[30]) );
  DFFHQX1 H6_reg_29_ ( .D(n3691), .CK(clk), .Q(H6[29]) );
  DFFHQXL H0_reg_29_ ( .D(n2898), .CK(clk), .Q(H0[29]) );
  DFFHQXL H4_reg_28_ ( .D(n2610), .CK(clk), .Q(H4[28]) );
  DFFHQXL H0_reg_27_ ( .D(n2900), .CK(clk), .Q(H0[27]) );
  DFFHQXL D_reg_31_ ( .D(n2735), .CK(clk), .Q(SHA256_result[159]) );
  DFFHQXL D_reg_30_ ( .D(n1583), .CK(clk), .Q(SHA256_result[158]) );
  DFFHQXL H1_reg_24_ ( .D(n2839), .CK(clk), .Q(H1[24]) );
  DFFHQXL H1_reg_25_ ( .D(n2838), .CK(clk), .Q(H1[25]) );
  DFFHQXL H6_reg_23_ ( .D(n2519), .CK(clk), .Q(H6[23]) );
  DFFHQXL H7_reg_24_ ( .D(n2423), .CK(clk), .Q(H7[24]) );
  DFFHQXL H7_reg_25_ ( .D(n2422), .CK(clk), .Q(H7[25]) );
  DFFHQX1 H1_reg_26_ ( .D(n3675), .CK(clk), .Q(H1[26]) );
  DFFHQX1 H1_reg_23_ ( .D(n3673), .CK(clk), .Q(H1[23]) );
  DFFHQX1 H2_reg_24_ ( .D(n3671), .CK(clk), .Q(H2[24]) );
  DFFHQX1 H5_reg_26_ ( .D(n3659), .CK(clk), .Q(H5[26]) );
  DFFHQX1 read_counter_reg_0_ ( .D(N3079), .CK(clk), .Q(read_counter[0]) );
  DFFHQXL H4_reg_24_ ( .D(n2614), .CK(clk), .Q(H4[24]) );
  DFFHQX1 H4_reg_25_ ( .D(n3682), .CK(clk), .Q(H4[25]) );
  DFFHQXL H5_reg_24_ ( .D(n2646), .CK(clk), .Q(H5[24]) );
  DFFHQXL H5_reg_27_ ( .D(n2643), .CK(clk), .Q(H5[27]) );
  DFFHQXL H0_reg_25_ ( .D(n2902), .CK(clk), .Q(H0[25]) );
  DFFHQXL H7_reg_23_ ( .D(n2424), .CK(clk), .Q(H7[23]) );
  DFFHQXL H5_reg_25_ ( .D(n2645), .CK(clk), .Q(H5[25]) );
  DFFHQXL H_reg_31_ ( .D(n1048), .CK(clk), .Q(SHA256_result[31]) );
  DFFHQXL D_reg_29_ ( .D(n2737), .CK(clk), .Q(SHA256_result[157]) );
  DFFHQX1 H4_reg_20_ ( .D(n3681), .CK(clk), .Q(H4[20]) );
  DFFHQXL H1_reg_22_ ( .D(n2841), .CK(clk), .Q(H1[22]) );
  DFFHQXL H1_reg_21_ ( .D(n2842), .CK(clk), .Q(H1[21]) );
  DFFHQX1 Kt_reg_30_ ( .D(N2976), .CK(clk), .Q(Kt[30]) );
  DFFHQXL H4_reg_17_ ( .D(n2621), .CK(clk), .Q(H4[17]) );
  DFFHQX1 H6_reg_22_ ( .D(n3636), .CK(clk), .Q(H6[22]) );
  DFFHQX1 H1_reg_20_ ( .D(n3651), .CK(clk), .Q(H1[20]) );
  DFFHQX1 H2_reg_20_ ( .D(n3655), .CK(clk), .Q(H2[20]) );
  DFFHQX1 H7_reg_19_ ( .D(n3643), .CK(clk), .Q(H7[19]) );
  DFFHQXL H4_reg_19_ ( .D(n2619), .CK(clk), .Q(H4[19]) );
  DFFHQXL H7_reg_22_ ( .D(n2425), .CK(clk), .Q(H7[22]) );
  DFFHQX1 H0_reg_20_ ( .D(n3676), .CK(clk), .Q(H0[20]) );
  DFFHQX1 H4_reg_16_ ( .D(n3667), .CK(clk), .Q(H4[16]) );
  DFFHQX1 H4_reg_21_ ( .D(n3680), .CK(clk), .Q(H4[21]) );
  DFFHQXL H7_reg_21_ ( .D(n2426), .CK(clk), .Q(H7[21]) );
  DFFHQX1 H0_reg_21_ ( .D(n3658), .CK(clk), .Q(H0[21]) );
  DFFHQXL H4_reg_18_ ( .D(n2620), .CK(clk), .Q(H4[18]) );
  DFFHQXL F_reg_31_ ( .D(n2671), .CK(clk), .Q(SHA256_result[95]) );
  DFFHQXL F_reg_30_ ( .D(n1551), .CK(clk), .Q(SHA256_result[94]) );
  DFFHQXL H_reg_30_ ( .D(n2449), .CK(clk), .Q(SHA256_result[30]) );
  DFFTRX1 round_reg_1_ ( .D(N122), .RN(n40), .CK(clk), .Q(round[1]), .QN(n2389) );
  DFFHQX1 Kt_reg_28_ ( .D(N2974), .CK(clk), .Q(Kt[28]) );
  DFFHQXL H5_reg_18_ ( .D(n2652), .CK(clk), .Q(H5[18]) );
  DFFHQXL H6_reg_17_ ( .D(n2525), .CK(clk), .Q(H6[17]) );
  DFFHQXL H0_reg_19_ ( .D(n2908), .CK(clk), .Q(H0[19]) );
  DFFHQXL H4_reg_14_ ( .D(n2624), .CK(clk), .Q(H4[14]) );
  DFFHQX1 H7_reg_16_ ( .D(n3650), .CK(clk), .Q(H7[16]) );
  DFFHQXL H4_reg_12_ ( .D(n2626), .CK(clk), .Q(H4[12]) );
  DFFHQX1 H4_reg_15_ ( .D(n3664), .CK(clk), .Q(H4[15]) );
  DFFHQX1 H0_reg_17_ ( .D(n3660), .CK(clk), .Q(H0[17]) );
  DFFHQXL H0_reg_16_ ( .D(n2911), .CK(clk), .Q(H0[16]) );
  DFFHQXL H6_reg_15_ ( .D(n2527), .CK(clk), .Q(H6[15]) );
  DFFHQX1 H4_reg_13_ ( .D(n3665), .CK(clk), .Q(H4[13]) );
  DFFHQXL H6_reg_16_ ( .D(n2526), .CK(clk), .Q(H6[16]) );
  DFFHQX1 H2_reg_16_ ( .D(n3649), .CK(clk), .Q(H2[16]) );
  DFFHQXL H0_reg_15_ ( .D(n2912), .CK(clk), .Q(H0[15]) );
  DFFTRX1 round_reg_4_ ( .D(N125), .RN(n40), .CK(clk), .Q(round[4]), .QN(n2388) );
  DFFTRX1 round_reg_0_ ( .D(N121), .RN(n40), .CK(clk), .Q(round[0]), .QN(n2398) );
  DFFTRX1 round_reg_5_ ( .D(N126), .RN(n40), .CK(clk), .Q(n995), .QN(n2391) );
  DFFHQX1 Kt_reg_26_ ( .D(N2972), .CK(clk), .Q(Kt[26]) );
  DFFHQXL H5_reg_14_ ( .D(n2656), .CK(clk), .Q(H5[14]) );
  DFFHQXL H5_reg_16_ ( .D(n2654), .CK(clk), .Q(H5[16]) );
  DFFHQXL H5_reg_13_ ( .D(n2657), .CK(clk), .Q(H5[13]) );
  DFFHQXL H6_reg_11_ ( .D(n2531), .CK(clk), .Q(H6[11]) );
  DFFHQXL H4_reg_6_ ( .D(n2632), .CK(clk), .Q(H4[6]) );
  DFFHQXL H0_reg_14_ ( .D(n2913), .CK(clk), .Q(H0[14]) );
  DFFHQXL H4_reg_3_ ( .D(n2635), .CK(clk), .Q(H4[3]) );
  DFFHQXL H4_reg_5_ ( .D(n2633), .CK(clk), .Q(H4[5]) );
  DFFHQXL H4_reg_9_ ( .D(n2629), .CK(clk), .Q(H4[9]) );
  DFFHQX1 H4_reg_8_ ( .D(n3661), .CK(clk), .Q(H4[8]) );
  DFFHQXL H6_reg_14_ ( .D(n2528), .CK(clk), .Q(H6[14]) );
  DFFHQXL H6_reg_12_ ( .D(n2530), .CK(clk), .Q(H6[12]) );
  DFFHQX1 H4_reg_7_ ( .D(n3662), .CK(clk), .Q(H4[7]) );
  DFFHQX1 H4_reg_11_ ( .D(n3663), .CK(clk), .Q(H4[11]) );
  DFFHQXL H0_reg_13_ ( .D(n2914), .CK(clk), .Q(H0[13]) );
  DFFHQXL H4_reg_0_ ( .D(n2638), .CK(clk), .Q(H4[0]) );
  DFFHQXL H4_reg_4_ ( .D(n2634), .CK(clk), .Q(H4[4]) );
  DFFHQXL H5_reg_11_ ( .D(n2659), .CK(clk), .Q(H5[11]) );
  DFFHQXL H6_reg_7_ ( .D(n2535), .CK(clk), .Q(H6[7]) );
  DFFHQXL H6_reg_8_ ( .D(n2534), .CK(clk), .Q(H6[8]) );
  DFFHQX1 H2_reg_10_ ( .D(n3645), .CK(clk), .Q(H2[10]) );
  DFFHQX1 H3_reg_11_ ( .D(n3657), .CK(clk), .Q(H3[11]) );
  DFFHQX1 H6_reg_10_ ( .D(n3635), .CK(clk), .Q(H6[10]) );
  DFFHQXL H0_reg_6_ ( .D(n2921), .CK(clk), .Q(H0[6]) );
  DFFHQXL H4_reg_1_ ( .D(n2637), .CK(clk), .Q(H4[1]) );
  DFFHQXL H4_reg_2_ ( .D(n2636), .CK(clk), .Q(H4[2]) );
  DFFHQXL H0_reg_9_ ( .D(n2918), .CK(clk), .Q(H0[9]) );
  DFFHQXL H0_reg_10_ ( .D(n2917), .CK(clk), .Q(H0[10]) );
  DFFHQXL H0_reg_5_ ( .D(n2922), .CK(clk), .Q(H0[5]) );
  DFFHQXL H1_reg_7_ ( .D(n2856), .CK(clk), .Q(H1[7]) );
  DFFHQXL H6_reg_5_ ( .D(n2537), .CK(clk), .Q(H6[5]) );
  DFFHQXL H7_reg_4_ ( .D(n2443), .CK(clk), .Q(H7[4]) );
  DFFHQXL H6_reg_3_ ( .D(n2539), .CK(clk), .Q(H6[3]) );
  DFFHQX1 H5_reg_7_ ( .D(n2663), .CK(clk), .Q(H5[7]) );
  DFFHQX1 H6_reg_6_ ( .D(n3638), .CK(clk), .Q(H6[6]) );
  DFFHQX1 H7_reg_6_ ( .D(n3597), .CK(clk), .Q(H7[6]) );
  DFFHQX1 H7_reg_7_ ( .D(n3644), .CK(clk), .Q(H7[7]) );
  DFFHQX1 H6_reg_4_ ( .D(n3637), .CK(clk), .Q(H6[4]) );
  DFFHQX1 H7_reg_5_ ( .D(n3617), .CK(clk), .Q(H7[5]) );
  DFFHQXL H2_reg_5_ ( .D(n2570), .CK(clk), .Q(H2[5]) );
  DFFHQX1 H1_reg_5_ ( .D(n3653), .CK(clk), .Q(H1[5]) );
  DFFHQXL H2_reg_4_ ( .D(n2571), .CK(clk), .Q(H2[4]) );
  DFFHQX1 H1_reg_4_ ( .D(n3590), .CK(clk), .Q(H1[4]) );
  DFFHQXL E_reg_23_ ( .D(n3559), .CK(clk), .Q(SHA256_result[119]) );
  DFFHQXL E_reg_24_ ( .D(n2710), .CK(clk), .Q(SHA256_result[120]) );
  DFFHQXL A_reg_30_ ( .D(n2865), .CK(clk), .Q(SHA256_result[254]) );
  DFFX1 F_reg_17_ ( .D(n1559), .CK(clk), .Q(n3807), .QN(n1151) );
  DFFX1 F_reg_15_ ( .D(n1560), .CK(clk), .Q(n3808), .QN(n1153) );
  DFFHQX1 Kt_reg_18_ ( .D(N2964), .CK(clk), .Q(Kt[18]) );
  DFFHQXL H5_reg_3_ ( .D(n2667), .CK(clk), .Q(H5[3]) );
  DFFHQXL H3_reg_5_ ( .D(n2601), .CK(clk), .Q(H3[5]) );
  DFFHQX1 H1_reg_3_ ( .D(n3654), .CK(clk), .Q(H1[3]) );
  DFFHQX1 H2_reg_2_ ( .D(n3626), .CK(clk), .Q(H2[2]) );
  DFFHQX1 H2_reg_3_ ( .D(n3642), .CK(clk), .Q(H2[3]) );
  DFFHQX1 H6_reg_2_ ( .D(n3639), .CK(clk), .Q(H6[2]) );
  DFFHQX1 H7_reg_2_ ( .D(n3620), .CK(clk), .Q(H7[2]) );
  DFFHQX1 H5_reg_2_ ( .D(n2668), .CK(clk), .Q(H5[2]) );
  DFFHQX1 H3_reg_4_ ( .D(n2602), .CK(clk), .Q(H3[4]) );
  DFFHQX1 H3_reg_6_ ( .D(n3594), .CK(clk), .Q(H3[6]) );
  DFFHQX1 H3_reg_3_ ( .D(n2603), .CK(clk), .Q(H3[3]) );
  DFFHQX1 H_reg_14_ ( .D(n2465), .CK(clk), .Q(SHA256_result[14]) );
  DFFHQX1 B_reg_14_ ( .D(n1575), .CK(clk), .Q(SHA256_result[206]) );
  DFFHQXL A_reg_29_ ( .D(n2866), .CK(clk), .Q(SHA256_result[253]) );
  DFFHQXL A_reg_28_ ( .D(n3571), .CK(clk), .Q(SHA256_result[252]) );
  DFFHQXL E_reg_30_ ( .D(n2704), .CK(clk), .Q(SHA256_result[126]) );
  DFFHQXL E_reg_29_ ( .D(n3555), .CK(clk), .Q(SHA256_result[125]) );
  DFFHQX1 digest_reg_31_ ( .D(N3078), .CK(clk), .Q(digest[31]) );
  DFFHQX1 digest_reg_30_ ( .D(N3077), .CK(clk), .Q(digest[30]) );
  DFFHQX1 digest_reg_29_ ( .D(N3076), .CK(clk), .Q(digest[29]) );
  DFFHQX1 digest_reg_28_ ( .D(N3075), .CK(clk), .Q(digest[28]) );
  DFFHQX1 digest_reg_27_ ( .D(N3074), .CK(clk), .Q(digest[27]) );
  DFFHQX1 digest_reg_26_ ( .D(N3073), .CK(clk), .Q(digest[26]) );
  DFFHQX1 digest_reg_25_ ( .D(N3072), .CK(clk), .Q(digest[25]) );
  DFFHQX1 digest_reg_24_ ( .D(N3071), .CK(clk), .Q(digest[24]) );
  DFFHQX1 digest_reg_23_ ( .D(N3070), .CK(clk), .Q(digest[23]) );
  DFFHQX1 digest_reg_22_ ( .D(N3069), .CK(clk), .Q(digest[22]) );
  DFFHQX1 digest_reg_21_ ( .D(N3068), .CK(clk), .Q(digest[21]) );
  DFFHQX1 digest_reg_20_ ( .D(N3067), .CK(clk), .Q(digest[20]) );
  DFFHQX1 digest_reg_19_ ( .D(N3066), .CK(clk), .Q(digest[19]) );
  DFFHQX1 digest_reg_18_ ( .D(N3065), .CK(clk), .Q(digest[18]) );
  DFFHQX1 digest_reg_17_ ( .D(N3064), .CK(clk), .Q(digest[17]) );
  DFFHQX1 digest_reg_16_ ( .D(N3063), .CK(clk), .Q(digest[16]) );
  DFFHQX1 digest_reg_15_ ( .D(N3062), .CK(clk), .Q(digest[15]) );
  DFFHQX1 digest_reg_14_ ( .D(N3061), .CK(clk), .Q(digest[14]) );
  DFFHQX1 digest_reg_13_ ( .D(N3060), .CK(clk), .Q(digest[13]) );
  DFFHQX1 digest_reg_12_ ( .D(N3059), .CK(clk), .Q(digest[12]) );
  DFFHQX1 digest_reg_11_ ( .D(N3058), .CK(clk), .Q(digest[11]) );
  DFFHQX1 digest_reg_10_ ( .D(N3057), .CK(clk), .Q(digest[10]) );
  DFFHQX1 digest_reg_9_ ( .D(N3056), .CK(clk), .Q(digest[9]) );
  DFFHQX1 digest_reg_8_ ( .D(N3055), .CK(clk), .Q(digest[8]) );
  DFFHQX1 digest_reg_7_ ( .D(N3054), .CK(clk), .Q(digest[7]) );
  DFFHQX1 digest_reg_6_ ( .D(N3053), .CK(clk), .Q(digest[6]) );
  DFFHQX1 digest_reg_5_ ( .D(N3052), .CK(clk), .Q(digest[5]) );
  DFFHQX1 digest_reg_4_ ( .D(N3051), .CK(clk), .Q(digest[4]) );
  DFFHQX1 digest_reg_3_ ( .D(N3050), .CK(clk), .Q(digest[3]) );
  DFFHQX1 digest_reg_2_ ( .D(N3049), .CK(clk), .Q(digest[2]) );
  DFFHQX1 digest_reg_1_ ( .D(N3048), .CK(clk), .Q(digest[1]) );
  DFFHQX1 digest_reg_0_ ( .D(N3047), .CK(clk), .Q(digest[0]) );
  DFFHQX1 G_reg_18_ ( .D(n1629), .CK(clk), .Q(SHA256_result[50]) );
  DFFHQX1 Kt_reg_20_ ( .D(N2966), .CK(clk), .Q(Kt[20]) );
  DFFHQX1 Kt_reg_19_ ( .D(N2965), .CK(clk), .Q(Kt[19]) );
  DFFHQXL D_reg_28_ ( .D(n1584), .CK(clk), .Q(SHA256_result[156]) );
  DFFHQXL B_reg_30_ ( .D(n1570), .CK(clk), .Q(SHA256_result[222]) );
  DFFHQXL G_reg_31_ ( .D(n1049), .CK(clk), .Q(SHA256_result[63]) );
  DFFHQXL G_reg_30_ ( .D(n1623), .CK(clk), .Q(SHA256_result[62]) );
  DFFHQXL B_reg_29_ ( .D(n2802), .CK(clk), .Q(SHA256_result[221]) );
  DFFHQXL C_reg_29_ ( .D(n2769), .CK(clk), .Q(SHA256_result[189]) );
  DFFHQXL C_reg_30_ ( .D(n1611), .CK(clk), .Q(SHA256_result[190]) );
  DFFHQXL B_reg_28_ ( .D(n2803), .CK(clk), .Q(SHA256_result[220]) );
  DFFHQXL H_reg_28_ ( .D(n2451), .CK(clk), .Q(SHA256_result[28]) );
  DFFHQXL H_reg_29_ ( .D(n1596), .CK(clk), .Q(SHA256_result[29]) );
  DFFTRX1 round_reg_3_ ( .D(N124), .RN(n40), .CK(clk), .Q(round[3]), .QN(n2390) );
  DFFHQX4 H5_reg_1_ ( .D(n3647), .CK(clk), .Q(H5[1]) );
  DFFHQX4 H3_reg_0_ ( .D(n3615), .CK(clk), .Q(H3[0]) );
  DFFHQXL C_reg_31_ ( .D(n1050), .CK(clk), .Q(SHA256_result[191]) );
  DFFHQX4 H2_reg_1_ ( .D(n2574), .CK(clk), .Q(H2[1]) );
  DFFHQX4 H1_reg_1_ ( .D(n3591), .CK(clk), .Q(H1[1]) );
  DFFHQX4 H2_reg_0_ ( .D(n3623), .CK(clk), .Q(H2[0]) );
  DFFHQX4 H3_reg_1_ ( .D(n2605), .CK(clk), .Q(H3[1]) );
  DFFHQX4 H5_reg_0_ ( .D(n3598), .CK(clk), .Q(H5[0]) );
  DFFHQX4 H6_reg_1_ ( .D(n2541), .CK(clk), .Q(H6[1]) );
  DFFHQX4 H1_reg_0_ ( .D(n2863), .CK(clk), .Q(H1[0]) );
  DFFHQX4 H1_reg_2_ ( .D(n2861), .CK(clk), .Q(H1[2]) );
  DFFHQX4 H7_reg_1_ ( .D(n3648), .CK(clk), .Q(H7[1]) );
  DFFHQX4 H6_reg_0_ ( .D(n2542), .CK(clk), .Q(H6[0]) );
  DFFHQXL B_reg_31_ ( .D(n2800), .CK(clk), .Q(SHA256_result[223]) );
  DFFHQX4 H7_reg_0_ ( .D(n2447), .CK(clk), .Q(H7[0]) );
  DFFX4 E_reg_31_ ( .D(n3554), .CK(clk), .Q(n2682), .QN(n2683) );
  DFFHQX4 H7_reg_3_ ( .D(n2444), .CK(clk), .Q(H7[3]) );
  DFFTRXL round_reg_6_ ( .D(N127), .RN(n40), .CK(clk), .Q(round[6]), .QN(n3553) );
  DFFXL read_counter_reg_2_ ( .D(N3081), .CK(clk), .Q(read_counter[2]), .QN(
        n3723) );
  DFFHQXL Kt_reg_23_ ( .D(N2969), .CK(clk), .Q(Kt[23]) );
  DFFHQXL Kt_reg_21_ ( .D(N2967), .CK(clk), .Q(Kt[21]) );
  DFFHQXL Kt_reg_24_ ( .D(N2970), .CK(clk), .Q(Kt[24]) );
  DFFHQXL Kt_reg_31_ ( .D(N2977), .CK(clk), .Q(Kt[31]) );
  DFFHQXL G_reg_20_ ( .D(n1627), .CK(clk), .Q(SHA256_result[52]) );
  DFFHQXL Kt_reg_22_ ( .D(N2968), .CK(clk), .Q(Kt[22]) );
  DFFHQXL Kt_reg_29_ ( .D(N2975), .CK(clk), .Q(Kt[29]) );
  DFFHQXL Kt_reg_16_ ( .D(N2962), .CK(clk), .Q(Kt[16]) );
  DFFHQXL Kt_reg_25_ ( .D(N2971), .CK(clk), .Q(Kt[25]) );
  DFFHQXL Kt_reg_27_ ( .D(N2973), .CK(clk), .Q(Kt[27]) );
  DFFHQXL H7_reg_12_ ( .D(n3596), .CK(clk), .Q(H7[12]) );
  DFFHQXL H0_reg_7_ ( .D(n3601), .CK(clk), .Q(H0[7]) );
  DFFHQXL F_reg_22_ ( .D(n1555), .CK(clk), .Q(SHA256_result[86]) );
  AND2X1 round_reg_2__U2 ( .A(N123), .B(n40), .Y(n2680) );
  DFFX2 round_reg_2_ ( .D(n2680), .CK(clk), .Q(n996), .QN(n3165) );
  DFFXL D_reg_19_ ( .D(n2747), .CK(clk), .Q(SHA256_result[147]), .QN(n3773) );
  DFFXL D_reg_18_ ( .D(n2748), .CK(clk), .Q(SHA256_result[146]), .QN(n3772) );
  DFFXL D_reg_17_ ( .D(n2749), .CK(clk), .Q(SHA256_result[145]), .QN(n3787) );
  DFFXL D_reg_16_ ( .D(n2750), .CK(clk), .Q(SHA256_result[144]), .QN(n3781) );
  DFFXL H0_reg_1_ ( .D(n2926), .CK(clk), .Q(H0[1]) );
  DFFXL F_reg_21_ ( .D(n1556), .CK(clk), .Q(SHA256_result[85]) );
  DFFXL D_reg_21_ ( .D(n1588), .CK(clk), .Q(SHA256_result[149]) );
  DFFXL D_reg_24_ ( .D(n2742), .CK(clk), .Q(SHA256_result[152]), .QN(n3726) );
  DFFXL D_reg_22_ ( .D(n2744), .CK(clk), .Q(SHA256_result[150]), .QN(n3774) );
  DFFXL H_reg_24_ ( .D(n2455), .CK(clk), .Q(SHA256_result[24]), .QN(n3790) );
  DFFXL H_reg_23_ ( .D(n2456), .CK(clk), .Q(SHA256_result[23]), .QN(n3789) );
  DFFXL H_reg_22_ ( .D(n2457), .CK(clk), .Q(SHA256_result[22]), .QN(n3788) );
  DFFXL H_reg_21_ ( .D(n2458), .CK(clk), .Q(SHA256_result[21]), .QN(n3805) );
  DFFXL B_reg_20_ ( .D(n1573), .CK(clk), .Q(SHA256_result[212]), .QN(n3534) );
  DFFXL H_reg_11_ ( .D(n2468), .CK(clk), .Q(SHA256_result[11]), .QN(n3823) );
  DFFXL D_reg_25_ ( .D(n1586), .CK(clk), .Q(SHA256_result[153]) );
  DFFXL H0_reg_2_ ( .D(n2925), .CK(clk), .Q(H0[2]) );
  DFFXL H0_reg_0_ ( .D(n2927), .CK(clk), .Q(H0[0]) );
  DFFXL H_reg_19_ ( .D(n1599), .CK(clk), .Q(SHA256_result[19]) );
  DFFXL H_reg_20_ ( .D(n1598), .CK(clk), .Q(SHA256_result[20]) );
  DFFXL D_reg_2_ ( .D(n1594), .CK(clk), .Q(SHA256_result[130]) );
  DFFXL H_reg_25_ ( .D(n2454), .CK(clk), .Q(SHA256_result[25]), .QN(n3791) );
  DFFXL D_reg_20_ ( .D(n1589), .CK(clk), .Q(SHA256_result[148]) );
  DFFXL B_reg_11_ ( .D(n2820), .CK(clk), .Q(SHA256_result[203]), .QN(n3827) );
  DFFXL H_reg_18_ ( .D(n1600), .CK(clk), .Q(SHA256_result[18]) );
  DFFXL C_reg_26_ ( .D(n2772), .CK(clk), .Q(SHA256_result[186]), .QN(n3850) );
  DFFXL C_reg_22_ ( .D(n2776), .CK(clk), .Q(SHA256_result[182]), .QN(n3860) );
  DFFXL C_reg_21_ ( .D(n2777), .CK(clk), .Q(SHA256_result[181]), .QN(n3531) );
  DFFXL B_reg_26_ ( .D(n1571), .CK(clk), .Q(SHA256_result[218]) );
  DFFXL H_reg_12_ ( .D(n1604), .CK(clk), .Q(SHA256_result[12]) );
  DFFXL B_reg_10_ ( .D(n2821), .CK(clk), .Q(SHA256_result[202]), .QN(n3826) );
  DFFXL H_reg_13_ ( .D(n1603), .CK(clk), .Q(SHA256_result[13]) );
  DFFXL H2_reg_15_ ( .D(n2560), .CK(clk), .Q(H2[15]) );
  DFFXL H2_reg_14_ ( .D(n2561), .CK(clk), .Q(H2[14]) );
  DFFXL H2_reg_13_ ( .D(n2562), .CK(clk), .Q(H2[13]) );
  DFFXL H2_reg_12_ ( .D(n2563), .CK(clk), .Q(H2[12]) );
  DFFXL C_reg_19_ ( .D(n2779), .CK(clk), .Q(SHA256_result[179]), .QN(n3806) );
  DFFXL H2_reg_17_ ( .D(n2558), .CK(clk), .Q(H2[17]) );
  DFFXL H2_reg_26_ ( .D(n2549), .CK(clk), .Q(H2[26]) );
  DFFXL H2_reg_18_ ( .D(n2557), .CK(clk), .Q(H2[18]) );
  DFFXL H2_reg_9_ ( .D(n2566), .CK(clk), .Q(H2[9]) );
  DFFXL H2_reg_22_ ( .D(n2553), .CK(clk), .Q(H2[22]) );
  DFFXL G_reg_22_ ( .D(n1625), .CK(clk), .Q(SHA256_result[54]) );
  DFFXL G_reg_21_ ( .D(n1626), .CK(clk), .Q(SHA256_result[53]) );
  DFFXL H2_reg_19_ ( .D(n2556), .CK(clk), .Q(H2[19]) );
  DFFXL C_reg_25_ ( .D(n1612), .CK(clk), .Q(SHA256_result[185]), .QN(n3527) );
  DFFXL C_reg_24_ ( .D(n1613), .CK(clk), .Q(SHA256_result[184]) );
  DFFXL C_reg_23_ ( .D(n1614), .CK(clk), .Q(SHA256_result[183]), .QN(n3530) );
  DFFXL C_reg_17_ ( .D(n2781), .CK(clk), .Q(SHA256_result[177]), .QN(n3539) );
  DFFXL C_reg_18_ ( .D(n2780), .CK(clk), .Q(SHA256_result[178]), .QN(n3536) );
  DFFXL C_reg_12_ ( .D(n2786), .CK(clk), .Q(SHA256_result[172]), .QN(n3828) );
  DFFXL G_reg_27_ ( .D(n2484), .CK(clk), .Q(SHA256_result[59]), .QN(n3856) );
  DFFXL G_reg_26_ ( .D(n2485), .CK(clk), .Q(SHA256_result[58]), .QN(n3771) );
  DFFXL G_reg_25_ ( .D(n2486), .CK(clk), .Q(SHA256_result[57]), .QN(n3783) );
  DFFXL G_reg_24_ ( .D(n2487), .CK(clk), .Q(SHA256_result[56]), .QN(n3782) );
  DFFXL G_reg_23_ ( .D(n2488), .CK(clk), .Q(SHA256_result[55]), .QN(n3793) );
  DFFXL H2_reg_27_ ( .D(n2548), .CK(clk), .Q(H2[27]) );
  DFFXL H2_reg_21_ ( .D(n2554), .CK(clk), .Q(H2[21]) );
  DFFXL B_reg_23_ ( .D(n1572), .CK(clk), .Q(SHA256_result[215]), .QN(n3529) );
  DFFXL D_reg_23_ ( .D(n1587), .CK(clk), .Q(SHA256_result[151]) );
  DFFXL G_reg_15_ ( .D(n2496), .CK(clk), .Q(SHA256_result[47]), .QN(n3811) );
  DFFXL D_reg_9_ ( .D(n1591), .CK(clk), .Q(SHA256_result[137]) );
  DFFXL D_reg_10_ ( .D(n2756), .CK(clk), .Q(SHA256_result[138]), .QN(n3803) );
  DFFXL D_reg_8_ ( .D(n2758), .CK(clk), .Q(SHA256_result[136]), .QN(n3799) );
  DFFXL D_reg_14_ ( .D(n2752), .CK(clk), .Q(SHA256_result[142]), .QN(n3786) );
  DFFXL D_reg_13_ ( .D(n2753), .CK(clk), .Q(SHA256_result[141]), .QN(n3785) );
  DFFXL D_reg_12_ ( .D(n2754), .CK(clk), .Q(SHA256_result[140]), .QN(n3784) );
  DFFXL H4_reg_31_ ( .D(n3704), .CK(clk), .Q(H4[31]) );
  DFFXL H0_reg_22_ ( .D(n3700), .CK(clk), .Q(H0[22]) );
  DFFXL C_reg_20_ ( .D(n1615), .CK(clk), .Q(SHA256_result[180]), .QN(n3535) );
  DFFXL D_reg_26_ ( .D(n2740), .CK(clk), .Q(SHA256_result[154]), .QN(n3846) );
  DFFXL B_reg_12_ ( .D(n1576), .CK(clk), .Q(SHA256_result[204]) );
  DFFHQXL B_reg_19_ ( .D(n1574), .CK(clk), .Q(SHA256_result[211]) );
  DFFHQXL H7_reg_20_ ( .D(n3605), .CK(clk), .Q(H7[20]) );
  DFFHQXL H7_reg_18_ ( .D(n3625), .CK(clk), .Q(H7[18]) );
  DFFHQXL H7_reg_17_ ( .D(n3606), .CK(clk), .Q(H7[17]) );
  DFFHQXL H7_reg_9_ ( .D(n3624), .CK(clk), .Q(H7[9]) );
  DFFHQXL H6_reg_21_ ( .D(n3634), .CK(clk), .Q(H6[21]) );
  DFFHQXL H6_reg_20_ ( .D(n3631), .CK(clk), .Q(H6[20]) );
  DFFHQXL H6_reg_19_ ( .D(n3630), .CK(clk), .Q(H6[19]) );
  DFFHQXL H6_reg_18_ ( .D(n3629), .CK(clk), .Q(H6[18]) );
  DFFHQXL H6_reg_13_ ( .D(n3632), .CK(clk), .Q(H6[13]) );
  DFFHQXL H6_reg_9_ ( .D(n3633), .CK(clk), .Q(H6[9]) );
  DFFHQXL H7_reg_13_ ( .D(n3616), .CK(clk), .Q(H7[13]) );
  DFFHQXL G_reg_19_ ( .D(n1628), .CK(clk), .Q(SHA256_result[51]) );
  DFFHQXL Kt_reg_17_ ( .D(N2963), .CK(clk), .Q(Kt[17]) );
  DFFHQXL H_reg_17_ ( .D(n1601), .CK(clk), .Q(SHA256_result[17]) );
  DFFHQXL D_reg_6_ ( .D(n1593), .CK(clk), .Q(SHA256_result[134]) );
  DFFHQXL D_reg_7_ ( .D(n1592), .CK(clk), .Q(SHA256_result[135]) );
  DFFHQXL B_reg_15_ ( .D(n2816), .CK(clk), .Q(SHA256_result[207]) );
  DFFHQXL H_reg_15_ ( .D(n2464), .CK(clk), .Q(SHA256_result[15]) );
  DFFHQXL C_reg_15_ ( .D(n2783), .CK(clk), .Q(SHA256_result[175]) );
  DFFXL F_reg_26_ ( .D(n1553), .CK(clk), .Q(SHA256_result[90]), .QN(n1142) );
  DFFXL F_reg_23_ ( .D(n1554), .CK(clk), .Q(SHA256_result[87]), .QN(n1145) );
  DFFXL F_reg_27_ ( .D(n2675), .CK(clk), .Q(SHA256_result[91]), .QN(n1141) );
  DFFXL F_reg_24_ ( .D(n2678), .CK(clk), .Q(SHA256_result[88]), .QN(n1144) );
  DFFXL D_reg_15_ ( .D(n2751), .CK(clk), .Q(SHA256_result[143]), .QN(n3780) );
  DFFXL F_reg_20_ ( .D(n1557), .CK(clk), .Q(SHA256_result[84]), .QN(n3794) );
  DFFXL D_reg_11_ ( .D(n1590), .CK(clk), .Q(SHA256_result[139]) );
  DFFXL D_reg_3_ ( .D(n2763), .CK(clk), .Q(SHA256_result[131]), .QN(n3804) );
  DFFXL C_reg_11_ ( .D(n1617), .CK(clk), .Q(SHA256_result[171]), .QN(n3543) );
  DFFXL C_reg_10_ ( .D(n1618), .CK(clk), .Q(SHA256_result[170]) );
  DFFXL G_reg_14_ ( .D(n2497), .CK(clk), .Q(SHA256_result[46]), .QN(n3821) );
  DFFXL D_reg_1_ ( .D(n2765), .CK(clk), .Q(SHA256_result[129]), .QN(n3813) );
  DFFXL B_reg_24_ ( .D(n2807), .CK(clk), .Q(SHA256_result[216]), .QN(n3792) );
  DFFXL B_reg_25_ ( .D(n2806), .CK(clk), .Q(SHA256_result[217]), .QN(n3528) );
  DFFXL H_reg_8_ ( .D(n2471), .CK(clk), .Q(SHA256_result[8]), .QN(n3824) );
  DFFXL F_reg_13_ ( .D(n2689), .CK(clk), .Q(SHA256_result[77]), .QN(n3818) );
  DFFXL H3_reg_17_ ( .D(n2589), .CK(clk), .Q(H3[17]) );
  DFFXL H3_reg_16_ ( .D(n2590), .CK(clk), .Q(H3[16]) );
  DFFXL H3_reg_15_ ( .D(n2591), .CK(clk), .Q(H3[15]) );
  DFFXL H3_reg_14_ ( .D(n2592), .CK(clk), .Q(H3[14]) );
  DFFXL H3_reg_13_ ( .D(n2593), .CK(clk), .Q(H3[13]) );
  DFFXL H3_reg_12_ ( .D(n2594), .CK(clk), .Q(H3[12]) );
  DFFXL H3_reg_10_ ( .D(n2596), .CK(clk), .Q(H3[10]) );
  DFFXL H3_reg_8_ ( .D(n2598), .CK(clk), .Q(H3[8]) );
  DFFXL H1_reg_17_ ( .D(n2846), .CK(clk), .Q(H1[17]) );
  DFFXL H1_reg_16_ ( .D(n2847), .CK(clk), .Q(H1[16]) );
  DFFXL H1_reg_15_ ( .D(n2848), .CK(clk), .Q(H1[15]) );
  DFFXL H1_reg_13_ ( .D(n2850), .CK(clk), .Q(H1[13]) );
  DFFXL H1_reg_11_ ( .D(n2852), .CK(clk), .Q(H1[11]) );
  DFFXL H1_reg_10_ ( .D(n2853), .CK(clk), .Q(H1[10]) );
  DFFXL H1_reg_9_ ( .D(n2854), .CK(clk), .Q(H1[9]) );
  DFFXL H0_reg_30_ ( .D(n2897), .CK(clk), .Q(H0[30]) );
  DFFXL H1_reg_18_ ( .D(n2845), .CK(clk), .Q(H1[18]) );
  DFFXL G_reg_28_ ( .D(n2483), .CK(clk), .Q(SHA256_result[60]), .QN(n3855) );
  DFFXL B_reg_22_ ( .D(n2809), .CK(clk), .Q(SHA256_result[214]), .QN(n3533) );
  DFFXL B_reg_21_ ( .D(n2810), .CK(clk), .Q(SHA256_result[213]), .QN(n3532) );
  DFFXL B_reg_18_ ( .D(n2813), .CK(clk), .Q(SHA256_result[210]), .QN(n3537) );
  DFFXL B_reg_17_ ( .D(n2814), .CK(clk), .Q(SHA256_result[209]), .QN(n3541) );
  DFFXL H_reg_26_ ( .D(n1597), .CK(clk), .Q(SHA256_result[26]) );
  DFFXL C_reg_27_ ( .D(n2771), .CK(clk), .Q(SHA256_result[187]), .QN(n3852) );
  DFFXL B_reg_27_ ( .D(n2804), .CK(clk), .Q(SHA256_result[219]), .QN(n3551) );
  DFFXL H3_reg_31_ ( .D(n2575), .CK(clk), .Q(H3[31]) );
  DFFXL H3_reg_29_ ( .D(n2577), .CK(clk), .Q(H3[29]) );
  DFFXL H3_reg_26_ ( .D(n2580), .CK(clk), .Q(H3[26]) );
  DFFXL H3_reg_24_ ( .D(n2582), .CK(clk), .Q(H3[24]) );
  DFFXL H3_reg_22_ ( .D(n2584), .CK(clk), .Q(H3[22]) );
  DFFXL H3_reg_19_ ( .D(n2587), .CK(clk), .Q(H3[19]) );
  DFFXL H3_reg_18_ ( .D(n2588), .CK(clk), .Q(H3[18]) );
  DFFXL H2_reg_8_ ( .D(n2567), .CK(clk), .Q(H2[8]) );
  DFFXL H2_reg_6_ ( .D(n2569), .CK(clk), .Q(H2[6]) );
  DFFXL A_reg_21_ ( .D(n3576), .CK(clk), .Q(SHA256_result[245]) );
  DFFXL D_reg_27_ ( .D(n1585), .CK(clk), .Q(SHA256_result[155]) );
  DFFXL H0_reg_23_ ( .D(n3678), .CK(clk), .Q(H0[23]) );
  DFFXL F_reg_29_ ( .D(n1552), .CK(clk), .Q(SHA256_result[93]), .QN(n3848) );
  DFFXL H_reg_27_ ( .D(n2452), .CK(clk), .Q(SHA256_result[27]), .QN(n3854) );
  DFFXL C_reg_28_ ( .D(n2770), .CK(clk), .Q(SHA256_result[188]), .QN(n3853) );
  DFFXL G_reg_29_ ( .D(n1624), .CK(clk), .Q(SHA256_result[61]), .QN(n3851) );
  DFFXL H7_reg_15_ ( .D(n2432), .CK(clk), .Q(H7[15]) );
  DFFXL H7_reg_14_ ( .D(n2433), .CK(clk), .Q(H7[14]) );
  DFFXL H7_reg_11_ ( .D(n2436), .CK(clk), .Q(H7[11]) );
  DFFXL H7_reg_10_ ( .D(n2437), .CK(clk), .Q(H7[10]) );
  DFFXL H7_reg_8_ ( .D(n2439), .CK(clk), .Q(H7[8]) );
  DFFXL H6_reg_28_ ( .D(n2514), .CK(clk), .Q(H6[28]) );
  DFFXL H6_reg_27_ ( .D(n2515), .CK(clk), .Q(H6[27]) );
  DFFXL H6_reg_26_ ( .D(n2516), .CK(clk), .Q(H6[26]) );
  DFFXL H6_reg_25_ ( .D(n2517), .CK(clk), .Q(H6[25]) );
  DFFXL H6_reg_24_ ( .D(n2518), .CK(clk), .Q(H6[24]) );
  DFFXL C_reg_14_ ( .D(n2784), .CK(clk), .Q(SHA256_result[174]), .QN(n3814) );
  DFFXL D_reg_4_ ( .D(n2762), .CK(clk), .Q(SHA256_result[132]), .QN(n3801) );
  DFFXL H7_reg_31_ ( .D(n3687), .CK(clk), .Q(H7[31]) );
  DFFXL H4_reg_27_ ( .D(n3679), .CK(clk), .Q(H4[27]) );
  DFFXL H0_reg_28_ ( .D(n3703), .CK(clk), .Q(H0[28]) );
  DFFXL H0_reg_24_ ( .D(n3702), .CK(clk), .Q(H0[24]) );
  DFFXL H0_reg_18_ ( .D(n3677), .CK(clk), .Q(H0[18]) );
  DFFXL H0_reg_11_ ( .D(n3588), .CK(clk), .Q(H0[11]) );
  DFFXL H7_reg_29_ ( .D(n3690), .CK(clk), .Q(H7[29]) );
  DFFXL C_reg_16_ ( .D(n1616), .CK(clk), .Q(SHA256_result[176]) );
  DFFXL D_reg_5_ ( .D(n2761), .CK(clk), .Q(SHA256_result[133]), .QN(n3802) );
  DFFXL H4_reg_10_ ( .D(n3666), .CK(clk), .Q(H4[10]) );
  DFFXL H3_reg_25_ ( .D(n3668), .CK(clk), .Q(H3[25]) );
  DFFXL H3_reg_23_ ( .D(n3669), .CK(clk), .Q(H3[23]) );
  DFFXL H2_reg_23_ ( .D(n3672), .CK(clk), .Q(H2[23]) );
  DFFXL H_reg_16_ ( .D(n1602), .CK(clk), .Q(SHA256_result[16]) );
  DFFXL F_reg_19_ ( .D(n1558), .CK(clk), .Q(SHA256_result[83]), .QN(n3795) );
  DFFXL G_reg_17_ ( .D(n2494), .CK(clk), .Q(SHA256_result[49]), .QN(n3810) );
  DFFXL G_reg_16_ ( .D(n2495), .CK(clk), .Q(SHA256_result[48]), .QN(n3809) );
  DFFXL F_reg_18_ ( .D(n2684), .CK(clk), .Q(SHA256_result[82]), .QN(n3800) );
  DFFXL B_reg_16_ ( .D(n2815), .CK(clk), .Q(SHA256_result[208]), .QN(n3858) );
  DFFXL H5_reg_30_ ( .D(n3697), .CK(clk), .Q(H5[30]) );
  DFFXL H5_reg_29_ ( .D(n3692), .CK(clk), .Q(H5[29]) );
  DFFXL H5_reg_23_ ( .D(n3656), .CK(clk), .Q(H5[23]) );
  DFFXL H5_reg_15_ ( .D(n3646), .CK(clk), .Q(H5[15]) );
  DFFXL H5_reg_12_ ( .D(n3627), .CK(clk), .Q(H5[12]) );
  DFFXL H5_reg_5_ ( .D(n3600), .CK(clk), .Q(H5[5]) );
  DFFXL H5_reg_4_ ( .D(n3604), .CK(clk), .Q(H5[4]) );
  DFFXL H4_reg_29_ ( .D(n3683), .CK(clk), .Q(H4[29]) );
  DFFXL H4_reg_26_ ( .D(n3685), .CK(clk), .Q(H4[26]) );
  DFFXL H4_reg_23_ ( .D(n3684), .CK(clk), .Q(H4[23]) );
  DFFXL H4_reg_22_ ( .D(n3686), .CK(clk), .Q(H4[22]) );
  DFFXL H3_reg_28_ ( .D(n3693), .CK(clk), .Q(H3[28]) );
  DFFXL H3_reg_7_ ( .D(n3595), .CK(clk), .Q(H3[7]) );
  DFFXL H2_reg_11_ ( .D(n3640), .CK(clk), .Q(H2[11]) );
  DFFXL H2_reg_7_ ( .D(n3641), .CK(clk), .Q(H2[7]) );
  DFFXL H1_reg_19_ ( .D(n3652), .CK(clk), .Q(H1[19]) );
  DFFXL H1_reg_6_ ( .D(n3592), .CK(clk), .Q(H1[6]) );
  DFFXL H0_reg_12_ ( .D(n3587), .CK(clk), .Q(H0[12]) );
  DFFXL H0_reg_8_ ( .D(n3586), .CK(clk), .Q(H0[8]) );
  DFFXL H0_reg_4_ ( .D(n3589), .CK(clk), .Q(H0[4]) );
  DFFXL H5_reg_17_ ( .D(n3618), .CK(clk), .Q(H5[17]) );
  DFFXL H5_reg_8_ ( .D(n3619), .CK(clk), .Q(H5[8]) );
  DFFXL H1_reg_12_ ( .D(n3622), .CK(clk), .Q(H1[12]) );
  DFFXL H0_reg_3_ ( .D(n3621), .CK(clk), .Q(H0[3]) );
  DFFXL H3_reg_20_ ( .D(n3628), .CK(clk), .Q(H3[20]) );
  DFFXL H2_reg_25_ ( .D(n3670), .CK(clk), .Q(H2[25]) );
  DFFXL H3_reg_21_ ( .D(n3593), .CK(clk), .Q(H3[21]) );
  DFFXL H5_reg_22_ ( .D(n3607), .CK(clk), .Q(H5[22]) );
  DFFXL H5_reg_20_ ( .D(n3609), .CK(clk), .Q(H5[20]) );
  DFFXL H5_reg_19_ ( .D(n3608), .CK(clk), .Q(H5[19]) );
  DFFXL H5_reg_9_ ( .D(n3611), .CK(clk), .Q(H5[9]) );
  DFFXL H1_reg_30_ ( .D(n3699), .CK(clk), .Q(H1[30]) );
  DFFXL H1_reg_14_ ( .D(n3602), .CK(clk), .Q(H1[14]) );
  DFFXL H1_reg_8_ ( .D(n3603), .CK(clk), .Q(H1[8]) );
  DFFXL H0_reg_26_ ( .D(n3701), .CK(clk), .Q(H0[26]) );
  DFFXL H5_reg_21_ ( .D(n3610), .CK(clk), .Q(H5[21]) );
  DFFXL H5_reg_10_ ( .D(n3612), .CK(clk), .Q(H5[10]) );
  DFFXL H5_reg_6_ ( .D(n3613), .CK(clk), .Q(H5[6]) );
  DFFXL H3_reg_30_ ( .D(n3696), .CK(clk), .Q(H3[30]) );
  DFFXL H3_reg_27_ ( .D(n3694), .CK(clk), .Q(H3[27]) );
  DFFXL H3_reg_9_ ( .D(n3614), .CK(clk), .Q(H3[9]) );
  DFFXL H2_reg_30_ ( .D(n3698), .CK(clk), .Q(H2[30]) );
  DFFXL H7_reg_26_ ( .D(n3674), .CK(clk), .Q(H7[26]) );
  DFFXL F_reg_16_ ( .D(n2686), .CK(clk), .Q(SHA256_result[80]), .QN(n1152) );
  DFFXL F_reg_28_ ( .D(n2674), .CK(clk), .Q(SHA256_result[92]), .QN(n1140) );
  DFFXL F_reg_25_ ( .D(n2677), .CK(clk), .Q(SHA256_result[89]), .QN(n1143) );
  DFFXL F_reg_14_ ( .D(n2688), .CK(clk), .Q(SHA256_result[78]), .QN(n1154) );
  DFFXL F_reg_7_ ( .D(n2695), .CK(clk), .Q(SHA256_result[71]), .QN(n1161) );
  DFFX4 F_reg_3_ ( .D(n2699), .CK(clk), .Q(SHA256_result[67]), .QN(n1165) );
  DFFXL H3_reg_2_ ( .D(n3599), .CK(clk), .Q(H3[2]) );
  DFFX1 F_reg_8_ ( .D(n1564), .CK(clk), .Q(SHA256_result[72]), .QN(n2401) );
  INVX3 U3 ( .A(n2801), .Y(n2384) );
  BUFX8 U4 ( .A(next_E[30]), .Y(n2405) );
  DLY1X1 U5 ( .A(next_A[9]), .Y(n2381) );
  NAND3X2 U6 ( .A(n3298), .B(n3297), .C(n3296), .Y(n2868) );
  NAND2X1 U7 ( .A(N822), .B(n2945), .Y(n3296) );
  AND2X4 U8 ( .A(N950), .B(n2382), .Y(n2727) );
  CLKINVX20 U9 ( .A(n2954), .Y(n2382) );
  DLY1X1 U10 ( .A(next_A[11]), .Y(n2383) );
  CLKBUFX8 U11 ( .A(SHA256_result[96]), .Y(n2934) );
  NAND3BX4 U12 ( .AN(n2799), .B(n2384), .C(n2385), .Y(n3555) );
  CLKINVX20 U13 ( .A(n2805), .Y(n2385) );
  AOI2BB2X1 U14 ( .B0(N986), .B1(n2935), .A0N(n2683), .A1N(n3062), .Y(n830) );
  NOR2BX4 U15 ( .AN(N952), .B(n2386), .Y(n2799) );
  CLKINVX20 U16 ( .A(n2387), .Y(n2386) );
  NAND2X1 U17 ( .A(N951), .B(n2946), .Y(n3359) );
  CLKINVX20 U18 ( .A(n2963), .Y(n2387) );
  BUFX12 U19 ( .A(next_E[28]), .Y(n2826) );
  OAI21X2 U20 ( .A0(SHA256_result[235]), .A1(SHA256_result[171]), .B0(
        SHA256_result[203]), .Y(n3221) );
  OAI21X2 U21 ( .A0(SHA256_result[170]), .A1(SHA256_result[234]), .B0(
        SHA256_result[202]), .Y(n3222) );
  INVX1 U22 ( .A(n3129), .Y(n3121) );
  INVX1 U23 ( .A(n3128), .Y(n3120) );
  INVX1 U24 ( .A(n3130), .Y(n3125) );
  NOR2X1 U25 ( .A(n3714), .B(round[4]), .Y(n1419) );
  NOR2X2 U26 ( .A(n2931), .B(n996), .Y(n1384) );
  NOR2X1 U27 ( .A(n3760), .B(n1320), .Y(n2711) );
  INVX1 U28 ( .A(n2817), .Y(n1250) );
  INVXL U29 ( .A(n2887), .Y(n2406) );
  NOR2BX2 U30 ( .AN(n3013), .B(first_block), .Y(n494) );
  NAND2XL U31 ( .A(n3168), .B(n3170), .Y(n3169) );
  NOR2X1 U32 ( .A(n3779), .B(n2932), .Y(n1408) );
  OR3X2 U33 ( .A(n495), .B(round[6]), .C(n656), .Y(n2825) );
  NOR2X1 U34 ( .A(n3770), .B(round[0]), .Y(n972) );
  AOI222X1 U35 ( .A0(n2718), .A1(n1260), .B0(n2766), .B1(n1419), .C0(n1261), 
        .C1(n2755), .Y(n1418) );
  INVX1 U36 ( .A(n3128), .Y(n3119) );
  CLKBUFX8 U37 ( .A(SHA256_result[245]), .Y(n2891) );
  CLKINVX3 U38 ( .A(n3152), .Y(n3150) );
  BUFX12 U39 ( .A(SHA256_result[32]), .Y(n2827) );
  AOI222X1 U40 ( .A0(n1467), .A1(n2757), .B0(n1475), .B1(n2718), .C0(n3707), 
        .C1(n1354), .Y(n1512) );
  INVX2 U41 ( .A(SHA256_result[43]), .Y(n3831) );
  INVX1 U42 ( .A(n3068), .Y(n3029) );
  OAI2BB1X1 U43 ( .A0N(H7[3]), .A1N(n3140), .B0(n953), .Y(n2444) );
  OAI2BB1X1 U44 ( .A0N(H7[0]), .A1N(n3139), .B0(n952), .Y(n2447) );
  OAI2BB1X1 U45 ( .A0N(H1[2]), .A1N(n3141), .B0(n711), .Y(n2861) );
  OAI2BB1X1 U46 ( .A0N(H1[0]), .A1N(n3141), .B0(n710), .Y(n2863) );
  OAI2BB1X1 U47 ( .A0N(H6[1]), .A1N(n3138), .B0(n900), .Y(n2541) );
  OAI2BB1X1 U48 ( .A0N(H3[1]), .A1N(n3140), .B0(n860), .Y(n2605) );
  OAI2BB1X1 U49 ( .A0N(H2[1]), .A1N(n3139), .B0(n879), .Y(n2574) );
  INVX1 U50 ( .A(SHA256_result[191]), .Y(n2402) );
  INVX1 U51 ( .A(n3157), .Y(n2403) );
  AOI222X1 U52 ( .A0(n3091), .A1(n1286), .B0(n1287), .B1(n2714), .C0(n2755), 
        .C1(n1289), .Y(n1285) );
  NAND2X1 U53 ( .A(SHA256_result[31]), .B(n3157), .Y(n2707) );
  INVX1 U54 ( .A(n558), .Y(n3682) );
  AOI222X1 U55 ( .A0(n3743), .A1(n2755), .B0(n2711), .B1(n1296), .C0(n2712), 
        .C1(n1265), .Y(n1501) );
  AOI222X1 U56 ( .A0(n2755), .A1(n1455), .B0(n1316), .B1(n3165), .C0(n3090), 
        .C1(n1456), .Y(n1451) );
  AOI222X1 U57 ( .A0(n1321), .A1(n3707), .B0(n3711), .B1(n1354), .C0(n1334), 
        .C1(n2755), .Y(n1435) );
  INVXL U58 ( .A(n3706), .Y(n3025) );
  INVXL U59 ( .A(n2719), .Y(n2996) );
  OR2XL U60 ( .A(n2823), .B(n3169), .Y(n495) );
  INVX1 U61 ( .A(n2828), .Y(n3115) );
  INVXL U62 ( .A(n2719), .Y(n2998) );
  INVXL U63 ( .A(n2719), .Y(n2997) );
  CLKINVX3 U64 ( .A(n3163), .Y(n3157) );
  INVXL U65 ( .A(n2764), .Y(n2971) );
  INVX1 U66 ( .A(n660), .Y(n3130) );
  INVX1 U67 ( .A(n660), .Y(n3127) );
  INVX1 U68 ( .A(n660), .Y(n3129) );
  INVXL U69 ( .A(n2764), .Y(n2966) );
  INVXL U70 ( .A(n2764), .Y(n2972) );
  INVXL U71 ( .A(n2764), .Y(n2965) );
  INVXL U72 ( .A(n2719), .Y(n2999) );
  OR2XL U73 ( .A(n1320), .B(round[1]), .Y(n2817) );
  INVXL U74 ( .A(n2764), .Y(n2967) );
  INVXL U75 ( .A(n2764), .Y(n2974) );
  INVXL U76 ( .A(n2764), .Y(n2973) );
  INVX1 U77 ( .A(n3000), .Y(n3015) );
  OR3XL U78 ( .A(N3079), .B(read_counter[2]), .C(n3725), .Y(n2392) );
  NAND3X1 U79 ( .A(read_counter[2]), .B(n3725), .C(n1237), .Y(n2393) );
  NAND3X1 U80 ( .A(n3725), .B(n3723), .C(n1237), .Y(n2394) );
  NAND3X1 U81 ( .A(n1078), .B(n3723), .C(n1081), .Y(n2395) );
  NAND3X1 U82 ( .A(read_counter[1]), .B(n3723), .C(n1237), .Y(n2396) );
  NAND2X1 U83 ( .A(n1080), .B(n1237), .Y(n2397) );
  INVXL U84 ( .A(n3023), .Y(n3064) );
  AND2X2 U85 ( .A(n3352), .B(n3351), .Y(n2399) );
  AND2X4 U86 ( .A(n3374), .B(n3375), .Y(n2400) );
  INVXL U87 ( .A(n1320), .Y(n3090) );
  OAI2BB1X2 U88 ( .A0N(SHA256_result[193]), .A1N(SHA256_result[161]), .B0(
        n3231), .Y(f2_ABC_32[1]) );
  OAI21X1 U89 ( .A0(SHA256_result[193]), .A1(SHA256_result[161]), .B0(n2906), 
        .Y(n3231) );
  AOI2BB2X4 U90 ( .B0(N890), .B1(n2937), .A0N(n2402), .A1N(n2403), .Y(n969) );
  OAI2BB1X4 U91 ( .A0N(n3078), .A1N(SHA256_result[223]), .B0(n969), .Y(n1050)
         );
  DLY1X1 U92 ( .A(next_A[10]), .Y(n2404) );
  CLKINVX2 U93 ( .A(n2954), .Y(n2946) );
  OR3X4 U94 ( .A(n2727), .B(n2736), .C(n2738), .Y(n3556) );
  OAI211X2 U95 ( .A0(n2979), .A1(n3857), .B0(n830), .C0(n3112), .Y(n2671) );
  AOI2BB2X4 U96 ( .B0(N858), .B1(n2939), .A0N(n2406), .A1N(n3064), .Y(n747) );
  INVX2 U97 ( .A(n2959), .Y(n2945) );
  BUFX3 U98 ( .A(T1_32_2_), .Y(n2697) );
  CLKINVX4 U99 ( .A(T1_32_16_), .Y(n2692) );
  CLKBUFX8 U100 ( .A(SHA256_result[103]), .Y(n2830) );
  DLY1X1 U101 ( .A(SHA256_result[121]), .Y(n2883) );
  OR3X4 U102 ( .A(n2739), .B(n2741), .C(n2743), .Y(n3558) );
  AND2X1 U103 ( .A(next_E[29]), .B(n3036), .Y(n2801) );
  OAI211X2 U104 ( .A0(n3842), .A1(n3706), .B0(n2707), .C0(n2705), .Y(n1048) );
  MXI2X4 U105 ( .A(SHA256_result[32]), .B(SHA256_result[64]), .S0(
        SHA256_result[96]), .Y(n2681) );
  INVX8 U106 ( .A(n2681), .Y(f1_EFG_32[0]) );
  INVXL U107 ( .A(n3315), .Y(n2685) );
  NAND2X4 U108 ( .A(N1018), .B(n2937), .Y(n2708) );
  INVX2 U109 ( .A(T1_32_11_), .Y(n2687) );
  CLKINVX4 U110 ( .A(n2687), .Y(n2690) );
  CLKINVX2 U111 ( .A(T1_32_14_), .Y(n2698) );
  XOR3X4 U112 ( .A(n2901), .B(n2892), .C(SHA256_result[237]), .Y(f3_A_32[0])
         );
  BUFX12 U113 ( .A(T1_32_27_), .Y(n2694) );
  INVX3 U114 ( .A(SHA256_result[33]), .Y(n3315) );
  CLKINVX3 U115 ( .A(n2692), .Y(n2693) );
  NAND2X4 U116 ( .A(N825), .B(n2945), .Y(n3293) );
  NAND3X4 U117 ( .A(n3293), .B(n3294), .C(n3295), .Y(n2865) );
  NAND2X2 U118 ( .A(N824), .B(n2944), .Y(n3263) );
  BUFX8 U119 ( .A(N110), .Y(n2696) );
  NAND2XL U120 ( .A(N821), .B(n2946), .Y(n3456) );
  NAND3X2 U121 ( .A(n3263), .B(n3264), .C(n3265), .Y(n2866) );
  NAND2X4 U122 ( .A(N953), .B(n2945), .Y(n3350) );
  NAND2X4 U123 ( .A(n3350), .B(n2399), .Y(n2704) );
  NAND2X1 U124 ( .A(next_A[27]), .B(n3037), .Y(n3297) );
  INVX4 U125 ( .A(n2698), .Y(n2701) );
  NAND2X4 U126 ( .A(n2400), .B(n3376), .Y(n3570) );
  OAI211X2 U127 ( .A0(n2975), .A1(n3843), .B0(n3109), .C0(n747), .Y(n2800) );
  NAND3X2 U128 ( .A(n3359), .B(n3360), .C(n3361), .Y(n2706) );
  OAI21X4 U129 ( .A0(n3064), .A1(n3857), .B0(n970), .Y(n1049) );
  AND2X4 U130 ( .A(n2708), .B(n2709), .Y(n970) );
  NAND2XL U131 ( .A(n2826), .B(n3036), .Y(n3360) );
  OAI2BB1X4 U132 ( .A0N(n2947), .A1N(N954), .B0(n3397), .Y(n3554) );
  NOR2X2 U133 ( .A(n3765), .B(n1320), .Y(n2712) );
  AOI222X1 U134 ( .A0(n1442), .A1(n1250), .B0(n3711), .B1(n2721), .C0(n1281), 
        .C1(n2713), .Y(n1502) );
  AOI222X1 U135 ( .A0(n1395), .A1(n3707), .B0(n1390), .B1(n1250), .C0(n2713), 
        .C1(n1401), .Y(n1531) );
  AOI222X1 U136 ( .A0(n1337), .A1(n1250), .B0(n1281), .B1(n2713), .C0(n1266), 
        .C1(n2714), .Y(n1495) );
  NOR2X2 U137 ( .A(n3762), .B(n1320), .Y(n2713) );
  NAND2X4 U138 ( .A(N922), .B(n2967), .Y(n2702) );
  NAND2X2 U139 ( .A(SHA256_result[191]), .B(n3029), .Y(n2703) );
  AND2X4 U140 ( .A(n2702), .B(n2703), .Y(n785) );
  OAI211X2 U141 ( .A0(n2979), .A1(n3841), .B0(n3111), .C0(n785), .Y(n2735) );
  AOI22X1 U142 ( .A0(SHA256_result[128]), .A1(n3145), .B0(H3[0]), .B1(n3134), 
        .Y(n625) );
  NAND2X4 U143 ( .A(N1050), .B(n2966), .Y(n2705) );
  INVX2 U144 ( .A(n2955), .Y(n2937) );
  CLKINVX4 U145 ( .A(n2968), .Y(n2958) );
  CLKINVX2 U146 ( .A(n2970), .Y(n2954) );
  INVXL U147 ( .A(n2970), .Y(n2952) );
  INVXL U148 ( .A(n2968), .Y(n2959) );
  NAND2X1 U149 ( .A(SHA256_result[63]), .B(n3157), .Y(n2709) );
  INVX1 U150 ( .A(n3152), .Y(n3151) );
  INVX1 U151 ( .A(n3065), .Y(n3037) );
  INVX1 U152 ( .A(n3067), .Y(n3027) );
  INVXL U153 ( .A(n2995), .Y(n2993) );
  INVX1 U154 ( .A(n3074), .Y(n3073) );
  INVX1 U155 ( .A(n3075), .Y(n3071) );
  INVX1 U156 ( .A(n3017), .Y(n3003) );
  INVX1 U157 ( .A(n3026), .Y(n3018) );
  INVX1 U158 ( .A(n3706), .Y(n3026) );
  AOI221XL U159 ( .A0(n1443), .A1(n3165), .B0(n1419), .B1(n1384), .C0(n1507), 
        .Y(n1503) );
  BUFX8 U160 ( .A(SHA256_result[102]), .Y(n2833) );
  NAND3XL U161 ( .A(n3503), .B(n3502), .C(n3128), .Y(n2663) );
  NAND2BX2 U162 ( .AN(n656), .B(n3166), .Y(n3168) );
  AOI21XL U163 ( .A0(n2798), .A1(n2389), .B0(round[6]), .Y(n3166) );
  BUFX3 U164 ( .A(round[3]), .Y(n2931) );
  NAND2XL U165 ( .A(n3171), .B(n3170), .Y(n2719) );
  AOI211X1 U166 ( .A0(n2718), .A1(n1438), .B0(n1356), .C0(n3712), .Y(n1437) );
  AOI2BB1X1 U167 ( .A0N(n1298), .A1N(n2817), .B0(n3715), .Y(n1433) );
  INVX4 U168 ( .A(n656), .Y(n2746) );
  AOI31X1 U169 ( .A0(round[4]), .A1(n3777), .A2(n3707), .B0(n1505), .Y(n1504)
         );
  AOI22XL U170 ( .A0(n2755), .A1(n1496), .B0(n1497), .B1(n3165), .Y(n1494) );
  NAND2X1 U171 ( .A(N984), .B(n2947), .Y(n3268) );
  BUFX16 U172 ( .A(SHA256_result[113]), .Y(n2899) );
  BUFX16 U173 ( .A(SHA256_result[118]), .Y(n2910) );
  INVX1 U174 ( .A(n2991), .Y(n2975) );
  INVX1 U175 ( .A(n2994), .Y(n2982) );
  INVX1 U176 ( .A(n2995), .Y(n2994) );
  INVX1 U177 ( .A(n3075), .Y(n3070) );
  INVX1 U178 ( .A(n3076), .Y(n3069) );
  INVXL U179 ( .A(n2995), .Y(n2992) );
  INVX1 U180 ( .A(n3016), .Y(n3007) );
  NOR2X1 U181 ( .A(n3720), .B(n3778), .Y(n1356) );
  INVX1 U182 ( .A(n3016), .Y(n3006) );
  NOR2X2 U183 ( .A(n2389), .B(n1320), .Y(n2718) );
  NOR2X2 U184 ( .A(n2398), .B(n1320), .Y(n2714) );
  NOR3X1 U185 ( .A(n3719), .B(n3779), .C(n2391), .Y(n1481) );
  AOI22XL U186 ( .A0(n3711), .A1(n2390), .B0(n1420), .B1(n2718), .Y(n1470) );
  AOI31X1 U187 ( .A0(n2757), .A1(n1354), .A2(n1491), .B0(n1537), .Y(n1535) );
  AOI211X1 U188 ( .A0(n1250), .A1(n1417), .B0(n3713), .C0(n3715), .Y(n1416) );
  NAND2X2 U189 ( .A(N818), .B(n2945), .Y(n3400) );
  NAND2X2 U190 ( .A(N820), .B(n2946), .Y(n3299) );
  NAND2X1 U191 ( .A(N981), .B(n2947), .Y(n3238) );
  XOR3X2 U192 ( .A(n2899), .B(n2910), .C(n2837), .Y(f4_E_32[11]) );
  XOR3X2 U193 ( .A(n2875), .B(n2915), .C(n2843), .Y(f4_E_32[10]) );
  NOR2X2 U194 ( .A(n1320), .B(round[4]), .Y(n2757) );
  NAND2BX4 U195 ( .AN(n656), .B(output_enable), .Y(n3170) );
  AOI221X1 U196 ( .A0(n1336), .A1(n3165), .B0(n1250), .B1(n1401), .C0(n1463), 
        .Y(n1462) );
  NOR2X1 U197 ( .A(n3719), .B(n2932), .Y(n1443) );
  MX2X4 U198 ( .A(SHA256_result[35]), .B(SHA256_result[67]), .S0(n2843), .Y(
        f1_EFG_32[3]) );
  OAI21XL U199 ( .A0(n3052), .A1(n3547), .B0(n466), .Y(n1570) );
  OAI211X1 U200 ( .A0(n2976), .A1(n3721), .B0(n3109), .C0(n748), .Y(n2797) );
  OAI211X1 U201 ( .A0(n2982), .A1(n3820), .B0(n3112), .C0(n940), .Y(n2465) );
  OAI211X1 U202 ( .A0(n2982), .A1(n3823), .B0(n3112), .C0(n939), .Y(n2468) );
  OAI211X1 U203 ( .A0(n2975), .A1(n3822), .B0(n3112), .C0(n938), .Y(n2469) );
  OAI211X1 U204 ( .A0(n2976), .A1(n3829), .B0(n3109), .C0(n750), .Y(n2793) );
  OAI211X1 U205 ( .A0(n2975), .A1(n3538), .B0(n3108), .C0(n736), .Y(n2816) );
  OAI211X1 U206 ( .A0(n2975), .A1(n3832), .B0(n3108), .C0(n732), .Y(n2822) );
  INVXL U207 ( .A(n3019), .Y(n3077) );
  INVXL U208 ( .A(n2712), .Y(n3718) );
  INVXL U209 ( .A(n2713), .Y(n3717) );
  INVXL U210 ( .A(n3076), .Y(n3068) );
  AOI2BB1XL U211 ( .A0N(n1263), .A1N(n1386), .B0(n2817), .Y(n1385) );
  INVXL U212 ( .A(n2718), .Y(n3719) );
  OAI22XL U213 ( .A0(n3750), .A1(n3714), .B0(n3089), .B1(n3738), .Y(n1439) );
  AOI22XL U214 ( .A0(n1261), .A1(n2711), .B0(n1263), .B1(n2718), .Y(n1254) );
  INVXL U215 ( .A(n2968), .Y(n2960) );
  AOI2BB1XL U216 ( .A0N(n1351), .A1N(n1454), .B0(n3718), .Y(n1542) );
  AOI21XL U217 ( .A0(n3736), .A1(n3742), .B0(n3720), .Y(n1302) );
  AOI2BB1XL U218 ( .A0N(n1455), .A1N(n1334), .B0(n2817), .Y(n1482) );
  AOI21XL U219 ( .A0(n1317), .A1(n2713), .B0(n1318), .Y(n1313) );
  AOI2BB2XL U220 ( .B0(n2713), .B1(n1261), .A0N(n3089), .A1N(n1483), .Y(n1479)
         );
  AOI22XL U221 ( .A0(n1391), .A1(n2714), .B0(n3711), .B1(n2766), .Y(n1478) );
  NAND4XL U222 ( .A(n1423), .B(n1424), .C(n1425), .D(n1426), .Y(N2962) );
  AOI221XL U223 ( .A0(n1334), .A1(n2718), .B0(n1291), .B1(n2713), .C0(n1427), 
        .Y(n1426) );
  AOI22XL U224 ( .A0(n2714), .A1(n1276), .B0(n1277), .B1(n2718), .Y(n1272) );
  AOI31XL U225 ( .A0(n3753), .A1(n2390), .A2(n3707), .B0(n1274), .Y(n1273) );
  AOI22XL U226 ( .A0(n2713), .A1(n1422), .B0(n1411), .B1(n2391), .Y(n1414) );
  OR4X1 U227 ( .A(n1301), .B(n1357), .C(n1358), .D(n1359), .Y(N2968) );
  AOI31XL U228 ( .A0(n3768), .A1(n3767), .A2(n3728), .B0(n3719), .Y(n1358) );
  OAI33XL U229 ( .A0(n3720), .A1(n3777), .A2(n3737), .B0(n1244), .B1(n3164), 
        .B2(n3716), .Y(n1421) );
  INVXL U230 ( .A(n2757), .Y(n3709) );
  NAND2XL U231 ( .A(n1389), .B(n2757), .Y(n1382) );
  OAI32XL U232 ( .A0(n3709), .A1(n3777), .A2(n3765), .B0(n3716), .B1(n1476), 
        .Y(n1468) );
  AOI21XL U233 ( .A0(n1330), .A1(n3734), .B0(n3716), .Y(n1329) );
  AOI31XL U234 ( .A0(n2757), .A1(n996), .A2(n1248), .B0(n1249), .Y(n1239) );
  NOR2XL U235 ( .A(n1290), .B(n3714), .Y(n1432) );
  AOI22XL U236 ( .A0(n1280), .A1(n2711), .B0(n3090), .B1(n1472), .Y(n1471) );
  AOI2BB1XL U237 ( .A0N(n1296), .A1N(n1317), .B0(n3720), .Y(n1537) );
  INVXL U238 ( .A(n3000), .Y(n3014) );
  AOI22XL U239 ( .A0(n3090), .A1(n1538), .B0(n1321), .B1(n2718), .Y(n1534) );
  AOI221XL U240 ( .A0(n1337), .A1(n2712), .B0(n3707), .B1(n1308), .C0(n1370), 
        .Y(n1369) );
  AOI22XL U241 ( .A0(n1334), .A1(n2718), .B0(n1335), .B1(n2711), .Y(n1326) );
  NOR2XL U242 ( .A(n1290), .B(n1320), .Y(n1336) );
  AOI221XL U243 ( .A0(n3707), .A1(n1263), .B0(n3092), .B1(n1541), .C0(n1542), 
        .Y(n1540) );
  AOI22XL U244 ( .A0(n3090), .A1(n1527), .B0(n1281), .B1(n2714), .Y(n1522) );
  INVXL U245 ( .A(n3706), .Y(n3024) );
  INVXL U246 ( .A(n3706), .Y(n3023) );
  AOI221XL U247 ( .A0(n1395), .A1(n2712), .B0(n2711), .B1(n1351), .C0(n1396), 
        .Y(n1394) );
  AOI22XL U248 ( .A0(n2712), .A1(n1526), .B0(n1386), .B1(n3707), .Y(n1523) );
  AOI22XL U249 ( .A0(n1265), .A1(n3707), .B0(n1266), .B1(n2712), .Y(n1253) );
  NAND3XL U250 ( .A(n2721), .B(n2391), .C(n2711), .Y(n1529) );
  AOI22X1 U251 ( .A0(n1351), .A1(n1412), .B0(n1250), .B1(n1413), .Y(n1406) );
  AOI22XL U252 ( .A0(n3090), .A1(n1488), .B0(n1303), .B1(n2714), .Y(n1487) );
  AND2X1 U253 ( .A(n1260), .B(n2712), .Y(n1342) );
  NOR2X1 U254 ( .A(n2390), .B(n996), .Y(n2721) );
  INVXL U255 ( .A(next_E[0]), .Y(n3525) );
  XOR3X4 U256 ( .A(n2867), .B(n2872), .C(n2860), .Y(f4_E_32[4]) );
  XOR3X4 U257 ( .A(n2873), .B(n2864), .C(SHA256_result[104]), .Y(f4_E_32[2])
         );
  NAND2XL U258 ( .A(n2887), .B(n3159), .Y(n3374) );
  XOR3X4 U259 ( .A(SHA256_result[103]), .B(n2877), .C(n2859), .Y(f4_E_32[1])
         );
  XOR3X4 U260 ( .A(n2875), .B(n2871), .C(n2858), .Y(f4_E_32[5]) );
  AOI21XL U261 ( .A0(n2871), .A1(n2983), .B0(n3113), .Y(n3352) );
  AOI21XL U262 ( .A0(SHA256_result[251]), .A1(n2984), .B0(n3114), .Y(n3298) );
  NAND3X2 U263 ( .A(n2723), .B(n2724), .C(n2726), .Y(n3571) );
  NAND2X2 U264 ( .A(N823), .B(n2947), .Y(n2723) );
  NAND2XL U265 ( .A(next_A[28]), .B(n3037), .Y(n2724) );
  NAND2XL U266 ( .A(n2862), .B(n3160), .Y(n2726) );
  AND2X1 U267 ( .A(next_E[27]), .B(n3036), .Y(n2736) );
  AND2X1 U268 ( .A(n2864), .B(n3159), .Y(n2738) );
  NAND2XL U269 ( .A(n2877), .B(n3159), .Y(n3365) );
  NAND2XL U270 ( .A(next_E[26]), .B(n3036), .Y(n3366) );
  AOI21XL U271 ( .A0(n2874), .A1(n2983), .B0(n3113), .Y(n3361) );
  XOR3X4 U272 ( .A(n2878), .B(n2874), .C(n2869), .Y(f4_E_32[3]) );
  AOI21XL U273 ( .A0(n2857), .A1(n2983), .B0(n3113), .Y(n3301) );
  NAND2X2 U274 ( .A(N945), .B(n2945), .Y(n3447) );
  NAND2XL U275 ( .A(n2910), .B(n3158), .Y(n3445) );
  NAND2XL U276 ( .A(SHA256_result[90]), .B(n3160), .Y(n3236) );
  NAND2XL U277 ( .A(n2877), .B(n3037), .Y(n3237) );
  AND2X2 U278 ( .A(N948), .B(n2945), .Y(n2739) );
  AND2X1 U279 ( .A(next_E[25]), .B(n3036), .Y(n2741) );
  AND2X1 U280 ( .A(n2883), .B(n3159), .Y(n2743) );
  AOI31XL U281 ( .A0(n2714), .A1(n1384), .A2(n2932), .B0(n1385), .Y(n1383) );
  XOR3X4 U282 ( .A(n2923), .B(n2904), .C(SHA256_result[251]), .Y(f3_A_32[5])
         );
  XOR3X4 U283 ( .A(n2920), .B(n2862), .C(SHA256_result[243]), .Y(f3_A_32[6])
         );
  AND3X4 U284 ( .A(n2746), .B(n2389), .C(n2798), .Y(n2745) );
  NAND2XL U285 ( .A(n3157), .B(n2915), .Y(n3448) );
  NAND2XL U286 ( .A(next_E[21]), .B(n3035), .Y(n3449) );
  XOR3X4 U287 ( .A(n2907), .B(SHA256_result[244]), .C(n2849), .Y(f3_A_32[7])
         );
  XOR3X4 U288 ( .A(n2905), .B(n2903), .C(SHA256_result[238]), .Y(f3_A_32[1])
         );
  XOR3X4 U289 ( .A(n2928), .B(n2857), .C(SHA256_result[240]), .Y(f3_A_32[3])
         );
  XOR3X4 U290 ( .A(n2929), .B(n2888), .C(SHA256_result[239]), .Y(f3_A_32[2])
         );
  NAND2XL U291 ( .A(n2903), .B(n3159), .Y(n3398) );
  NAND2XL U292 ( .A(n2901), .B(n3159), .Y(n3393) );
  NOR2X2 U293 ( .A(n1320), .B(round[0]), .Y(n2755) );
  OAI22XL U294 ( .A0(n3720), .A1(n3741), .B0(n3775), .B1(n1382), .Y(n1463) );
  NAND2XL U295 ( .A(N808), .B(n2944), .Y(n3281) );
  OAI22XL U296 ( .A0(n1331), .A1(n1320), .B0(n2931), .B1(n3708), .Y(n1328) );
  XOR3X4 U297 ( .A(SHA256_result[234]), .B(n2891), .C(n2855), .Y(f3_A_32[8])
         );
  OAI211XL U298 ( .A0(n3746), .A1(n3719), .B0(n1338), .C0(n1339), .Y(N2970) );
  AOI211XL U299 ( .A0(n1340), .A1(n2755), .B0(n1341), .C0(n1342), .Y(n1339) );
  AOI21XL U300 ( .A0(n2714), .A1(n1355), .B0(n1464), .Y(n1461) );
  AOI222XL U301 ( .A0(n1386), .A1(n2718), .B0(n1317), .B1(n3707), .C0(n1454), 
        .C1(n2711), .Y(n1452) );
  AOI22XL U302 ( .A0(n1335), .A1(n2714), .B0(n1395), .B1(n2712), .Y(n1450) );
  NAND2XL U303 ( .A(n1356), .B(n2932), .Y(n1344) );
  AOI33XL U304 ( .A0(n1353), .A1(n996), .A2(n2755), .B0(n1354), .B1(n3745), 
        .B2(n1250), .Y(n1346) );
  AOI222XL U305 ( .A0(n1336), .A1(n3165), .B0(n3090), .B1(n1348), .C0(n1294), 
        .C1(n3707), .Y(n1347) );
  AOI22XL U306 ( .A0(n3090), .A1(n1498), .B0(n2711), .B1(n1246), .Y(n1493) );
  NAND2XL U307 ( .A(next_E[18]), .B(n3035), .Y(n3452) );
  NAND2XL U308 ( .A(n2904), .B(n3158), .Y(n3401) );
  NAND2XL U309 ( .A(SHA256_result[244]), .B(n3158), .Y(n3457) );
  NAND2XL U310 ( .A(N814), .B(n2944), .Y(n3287) );
  AOI221XL U311 ( .A0(n2714), .A1(n1408), .B0(n1324), .B1(n2757), .C0(n1409), 
        .Y(n1407) );
  AOI21XL U312 ( .A0(n2713), .A1(n1353), .B0(n1336), .Y(n1410) );
  NAND3XL U313 ( .A(n2766), .B(round[0]), .C(n2757), .Y(n1506) );
  AOI22XL U314 ( .A0(N838), .A1(n2965), .B0(SHA256_result[235]), .B1(n3033), 
        .Y(n734) );
  AOI31XL U315 ( .A0(n2796), .A1(n3770), .A2(n1508), .B0(n3089), .Y(n1507) );
  NAND2XL U316 ( .A(SHA256_result[234]), .B(n2989), .Y(n3439) );
  NAND3BXL U317 ( .AN(n3349), .B(n3108), .C(n3348), .Y(n2725) );
  NAND2XL U318 ( .A(n2869), .B(n2989), .Y(n3348) );
  NAND3BXL U319 ( .AN(n3386), .B(n3108), .C(n3385), .Y(n2893) );
  NAND2XL U320 ( .A(n2892), .B(n2989), .Y(n3385) );
  NAND3BXL U321 ( .AN(n3412), .B(n3108), .C(n3411), .Y(n2894) );
  NAND2XL U322 ( .A(n2985), .B(n2906), .Y(n3411) );
  NAND3BXL U323 ( .AN(n3444), .B(n3108), .C(n3443), .Y(n2886) );
  NAND2XL U324 ( .A(n2907), .B(n2990), .Y(n3443) );
  NAND3BXL U325 ( .AN(n3475), .B(n3108), .C(n3474), .Y(n2889) );
  NAND2XL U326 ( .A(n2924), .B(n2986), .Y(n3474) );
  NAND3BXL U327 ( .AN(n3479), .B(n3108), .C(n3478), .Y(n2890) );
  NAND2XL U328 ( .A(n2928), .B(n2990), .Y(n3478) );
  NAND3BXL U329 ( .AN(n3519), .B(n3108), .C(n3518), .Y(n2895) );
  NAND2XL U330 ( .A(n2933), .B(n2990), .Y(n3518) );
  NAND3XL U331 ( .A(n2759), .B(n3108), .C(n3526), .Y(n2734) );
  OR2X2 U332 ( .A(n2964), .B(n3524), .Y(n2759) );
  NAND2XL U333 ( .A(n2745), .B(n3553), .Y(n3171) );
  AOI22XL U334 ( .A0(N834), .A1(n2972), .B0(n2923), .B1(n3033), .Y(n731) );
  OAI211XL U335 ( .A0(n2979), .A1(n3831), .B0(n3112), .C0(n922), .Y(n2500) );
  OAI211XL U336 ( .A0(n2979), .A1(n3819), .B0(n3112), .C0(n923), .Y(n2499) );
  AOI22XL U337 ( .A0(N968), .A1(n2935), .B0(n2873), .B1(n3028), .Y(n822) );
  INVXL U338 ( .A(n447), .Y(n3162) );
  OAI211XL U339 ( .A0(n2981), .A1(n3810), .B0(n3112), .C0(n927), .Y(n2494) );
  AOI22XL U340 ( .A0(N1004), .A1(n2936), .B0(n3034), .B1(n3807), .Y(n927) );
  OAI211XL U341 ( .A0(n2979), .A1(n3800), .B0(n3111), .C0(n825), .Y(n2684) );
  AOI22XL U342 ( .A0(N973), .A1(n2935), .B0(SHA256_result[114]), .B1(n3028), 
        .Y(n825) );
  NAND3BXL U343 ( .AN(n3189), .B(n3112), .C(n3188), .Y(n2728) );
  NAND3BXL U344 ( .AN(n3192), .B(n3112), .C(n3191), .Y(n2543) );
  NAND3BXL U345 ( .AN(n3196), .B(n3112), .C(n3195), .Y(n2730) );
  NAND2XL U346 ( .A(n2837), .B(n2988), .Y(n3195) );
  INVXL U347 ( .A(next_E[4]), .Y(n3193) );
  NAND3BXL U348 ( .AN(n3200), .B(n3112), .C(n3199), .Y(n2729) );
  NAND2XL U349 ( .A(n2840), .B(n2985), .Y(n3199) );
  NAND3BXL U350 ( .AN(n3246), .B(n3112), .C(n3245), .Y(n2731) );
  INVXL U351 ( .A(next_E[3]), .Y(n3243) );
  NAND3BXL U352 ( .AN(n3250), .B(n3112), .C(n3249), .Y(n2732) );
  NAND2XL U353 ( .A(n2844), .B(n2985), .Y(n3249) );
  INVXL U354 ( .A(next_E[2]), .Y(n3247) );
  NAND3BXL U355 ( .AN(n3275), .B(n3112), .C(n3274), .Y(n2733) );
  NAND2XL U356 ( .A(n2851), .B(n2986), .Y(n3274) );
  INVXL U357 ( .A(next_E[1]), .Y(n3272) );
  NAND2XL U358 ( .A(n2873), .B(n3159), .Y(n3356) );
  AOI33XL U359 ( .A0(n2718), .A1(n3165), .A2(n3748), .B0(n2757), .B1(n996), 
        .B2(n1491), .Y(n1514) );
  AOI221XL U360 ( .A0(n1475), .A1(n2712), .B0(n3707), .B1(n1354), .C0(n1517), 
        .Y(n1516) );
  NAND2BXL U361 ( .AN(n3044), .B(n2851), .Y(n3511) );
  NAND2XL U362 ( .A(n3722), .B(n3159), .Y(n3510) );
  NAND2BXL U363 ( .AN(n3052), .B(n2859), .Y(n3435) );
  NAND2XL U364 ( .A(SHA256_result[76]), .B(n3158), .Y(n3434) );
  NAND2BXL U365 ( .AN(n2953), .B(N960), .Y(n3259) );
  NAND2BXL U366 ( .AN(n3062), .B(n2840), .Y(n3258) );
  NAND2XL U367 ( .A(SHA256_result[69]), .B(n3160), .Y(n3257) );
  NAND2XL U368 ( .A(n3837), .B(n3160), .Y(n3327) );
  NAND2BXL U369 ( .AN(n3061), .B(SHA256_result[104]), .Y(n3331) );
  NAND2XL U370 ( .A(SHA256_result[72]), .B(n3160), .Y(n3330) );
  AOI21XL U371 ( .A0(SHA256_result[240]), .A1(n2984), .B0(n3114), .Y(n3235) );
  NAND3X1 U372 ( .A(n2760), .B(n3501), .C(n3500), .Y(n1559) );
  OR2XL U373 ( .A(n3068), .B(n3499), .Y(n2760) );
  NAND2XL U374 ( .A(next_E[16]), .B(n3036), .Y(n3363) );
  NAND2XL U375 ( .A(SHA256_result[104]), .B(n3159), .Y(n3343) );
  NAND2XL U376 ( .A(SHA256_result[235]), .B(n3161), .Y(n3463) );
  NAND2XL U377 ( .A(n2920), .B(n3160), .Y(n3466) );
  NAND2XL U378 ( .A(n2923), .B(n3157), .Y(n3469) );
  NAND2XL U379 ( .A(n2929), .B(n3158), .Y(n3480) );
  NAND2XL U380 ( .A(n2919), .B(n3158), .Y(n3460) );
  NAND2XL U381 ( .A(n2905), .B(n3158), .Y(n3406) );
  NAND2XL U382 ( .A(n2858), .B(n3160), .Y(n3333) );
  NAND2BXL U383 ( .AN(n2954), .B(N930), .Y(n3185) );
  NAND2XL U384 ( .A(n2830), .B(n3157), .Y(n3183) );
  NAND2BXL U385 ( .AN(n3048), .B(n2872), .Y(n3497) );
  NAND2XL U386 ( .A(n3808), .B(n3157), .Y(n3496) );
  NAND2XL U387 ( .A(n2823), .B(n3170), .Y(n2764) );
  AOI222XL U388 ( .A0(n1491), .A1(n1337), .B0(n3165), .B1(n3757), .C0(n972), 
        .C1(round[1]), .Y(n1465) );
  AOI22XL U389 ( .A0(n3106), .A1(SHA256_result[89]), .B0(n3104), .B1(n2883), 
        .Y(n1118) );
  AOI22XL U390 ( .A0(n3106), .A1(SHA256_result[90]), .B0(n3104), .B1(n2877), 
        .Y(n1114) );
  AOI22XL U391 ( .A0(n3106), .A1(SHA256_result[91]), .B0(n3104), .B1(n2864), 
        .Y(n1110) );
  AOI22XL U392 ( .A0(n3106), .A1(SHA256_result[92]), .B0(n3104), .B1(n2874), 
        .Y(n1106) );
  INVXL U393 ( .A(n2828), .Y(n3114) );
  INVXL U394 ( .A(n2828), .Y(n3113) );
  AND2X1 U395 ( .A(n3105), .B(n2830), .Y(n3276) );
  AOI211XL U396 ( .A0(n996), .A1(n2388), .B0(n1386), .C0(n1261), .Y(n1446) );
  NOR3XL U397 ( .A(n996), .B(round[1]), .C(n3737), .Y(n1391) );
  NOR2X1 U398 ( .A(n3165), .B(n2931), .Y(n2766) );
  AOI22XL U399 ( .A0(N888), .A1(n2941), .B0(SHA256_result[221]), .B1(n3030), 
        .Y(n766) );
  INVXL U400 ( .A(n2855), .Y(n3547) );
  AOI22XL U401 ( .A0(N1048), .A1(n2944), .B0(SHA256_result[29]), .B1(n3156), 
        .Y(n498) );
  NAND2XL U402 ( .A(n3157), .B(SHA256_result[93]), .Y(n3266) );
  NAND2XL U403 ( .A(SHA256_result[94]), .B(n3160), .Y(n3269) );
  BUFX16 U404 ( .A(SHA256_result[99]), .Y(n2843) );
  BUFX16 U405 ( .A(SHA256_result[106]), .Y(n2867) );
  BUFX16 U406 ( .A(SHA256_result[112]), .Y(n2875) );
  MX2X4 U407 ( .A(SHA256_result[36]), .B(SHA256_result[68]), .S0(n2837), .Y(
        n418) );
  BUFX16 U408 ( .A(SHA256_result[227]), .Y(n2905) );
  NAND3X4 U409 ( .A(n1434), .B(n3553), .C(inner_busy), .Y(n1320) );
  AOI22XL U410 ( .A0(n3149), .A1(SHA256_result[176]), .B0(H2[16]), .B1(n3135), 
        .Y(n591) );
  AOI22XL U411 ( .A0(n3149), .A1(SHA256_result[16]), .B0(H7[16]), .B1(n3135), 
        .Y(n590) );
  AOI22XL U412 ( .A0(n3149), .A1(SHA256_result[19]), .B0(H7[19]), .B1(n3134), 
        .Y(n597) );
  AOI22XL U413 ( .A0(n3149), .A1(SHA256_result[54]), .B0(H6[22]), .B1(n3134), 
        .Y(n604) );
  AOI22XL U414 ( .A0(SHA256_result[156]), .A1(n3147), .B0(H3[28]), .B1(n3140), 
        .Y(n547) );
  AOI22XL U415 ( .A0(SHA256_result[153]), .A1(n3150), .B0(H3[25]), .B1(n3136), 
        .Y(n572) );
  AOI22XL U416 ( .A0(SHA256_result[69]), .A1(n3144), .B0(H5[5]), .B1(n3132), 
        .Y(n640) );
  AOI21XL U417 ( .A0(SHA256_result[179]), .A1(n3005), .B0(n3119), .Y(n891) );
  AOI21XL U418 ( .A0(SHA256_result[141]), .A1(n3006), .B0(n3121), .Y(n867) );
  AOI21XL U419 ( .A0(SHA256_result[213]), .A1(n3010), .B0(n3124), .Y(n721) );
  AOI21XL U420 ( .A0(SHA256_result[55]), .A1(n3003), .B0(n3117), .Y(n911) );
  AOI22XL U421 ( .A0(n3150), .A1(SHA256_result[18]), .B0(H7[18]), .B1(n3133), 
        .Y(n615) );
  AOI22XL U422 ( .A0(n3150), .A1(SHA256_result[17]), .B0(H7[17]), .B1(n3132), 
        .Y(n634) );
  AOI22XL U423 ( .A0(n3150), .A1(SHA256_result[50]), .B0(H6[18]), .B1(n3133), 
        .Y(n611) );
  AOI22XL U424 ( .A0(n3150), .A1(SHA256_result[20]), .B0(H7[20]), .B1(n3132), 
        .Y(n635) );
  AOI22XL U425 ( .A0(n3150), .A1(SHA256_result[53]), .B0(H6[21]), .B1(n3133), 
        .Y(n606) );
  AOI22XL U426 ( .A0(n3150), .A1(SHA256_result[52]), .B0(H6[20]), .B1(n3133), 
        .Y(n609) );
  AOI22XL U427 ( .A0(n3150), .A1(SHA256_result[51]), .B0(H6[19]), .B1(n3133), 
        .Y(n610) );
  AOI22XL U428 ( .A0(n3148), .A1(SHA256_result[184]), .B0(H2[24]), .B1(n3137), 
        .Y(n569) );
  AOI22XL U429 ( .A0(n3148), .A1(SHA256_result[26]), .B0(H7[26]), .B1(n3137), 
        .Y(n566) );
  AOI22XL U430 ( .A0(n3148), .A1(SHA256_result[63]), .B0(H6[31]), .B1(n3138), 
        .Y(n552) );
  AOI22XL U431 ( .A0(n3148), .A1(SHA256_result[191]), .B0(H2[31]), .B1(n3136), 
        .Y(n551) );
  AOI22XL U432 ( .A0(n3148), .A1(SHA256_result[61]), .B0(H6[29]), .B1(n3133), 
        .Y(n549) );
  AOI22XL U433 ( .A0(n3148), .A1(SHA256_result[62]), .B0(H6[30]), .B1(n3138), 
        .Y(n545) );
  AOI22XL U434 ( .A0(n3150), .A1(SHA256_result[31]), .B0(H7[31]), .B1(n3138), 
        .Y(n553) );
  AOI22XL U435 ( .A0(n3151), .A1(SHA256_result[29]), .B0(H7[29]), .B1(n3140), 
        .Y(n550) );
  AOI22XL U436 ( .A0(SHA256_result[72]), .A1(n3146), .B0(H5[8]), .B1(n3134), 
        .Y(n621) );
  AOI22XL U437 ( .A0(SHA256_result[76]), .A1(n3146), .B0(H5[12]), .B1(n3133), 
        .Y(n613) );
  AOI22XL U438 ( .A0(SHA256_result[204]), .A1(n3146), .B0(H1[12]), .B1(n3137), 
        .Y(n618) );
  AOI22XL U439 ( .A0(n3807), .A1(n3146), .B0(H5[17]), .B1(n3140), .Y(n622) );
  AOI22XL U440 ( .A0(SHA256_result[148]), .A1(n3146), .B0(H3[20]), .B1(n3133), 
        .Y(n612) );
  AOI22XL U441 ( .A0(SHA256_result[93]), .A1(n3146), .B0(H5[29]), .B1(n3138), 
        .Y(n548) );
  AOI22XL U442 ( .A0(SHA256_result[158]), .A1(n3146), .B0(H3[30]), .B1(n3138), 
        .Y(n544) );
  AOI22XL U443 ( .A0(SHA256_result[94]), .A1(n3146), .B0(H5[30]), .B1(n3138), 
        .Y(n543) );
  AOI22XL U444 ( .A0(SHA256_result[190]), .A1(n3146), .B0(H2[30]), .B1(n3138), 
        .Y(n542) );
  AOI22XL U445 ( .A0(SHA256_result[206]), .A1(n3145), .B0(H1[14]), .B1(n3132), 
        .Y(n638) );
  AOI22XL U446 ( .A0(SHA256_result[84]), .A1(n3145), .B0(H5[20]), .B1(n3132), 
        .Y(n631) );
  AOI22XL U447 ( .A0(SHA256_result[83]), .A1(n3145), .B0(H5[19]), .B1(n3132), 
        .Y(n632) );
  AOI22XL U448 ( .A0(SHA256_result[86]), .A1(n3145), .B0(H5[22]), .B1(n3132), 
        .Y(n633) );
  AOI22XL U449 ( .A0(SHA256_result[222]), .A1(n3145), .B0(H1[30]), .B1(n3138), 
        .Y(n541) );
  AOI22XL U450 ( .A0(SHA256_result[87]), .A1(n3147), .B0(H5[23]), .B1(n3135), 
        .Y(n584) );
  AOI22XL U451 ( .A0(n3808), .A1(n3147), .B0(H5[15]), .B1(n3135), .Y(n594) );
  AOI22XL U452 ( .A0(SHA256_result[180]), .A1(n3150), .B0(H2[20]), .B1(n3135), 
        .Y(n585) );
  AOI22XL U453 ( .A0(SHA256_result[212]), .A1(n3150), .B0(H1[20]), .B1(n3135), 
        .Y(n589) );
  AOI22XL U454 ( .A0(SHA256_result[211]), .A1(n3147), .B0(H1[19]), .B1(n3135), 
        .Y(n588) );
  AOI22XL U455 ( .A0(SHA256_result[185]), .A1(n3147), .B0(H2[25]), .B1(n3137), 
        .Y(n570) );
  AOI22XL U456 ( .A0(SHA256_result[215]), .A1(n3151), .B0(H1[23]), .B1(n3137), 
        .Y(n567) );
  AOI22XL U457 ( .A0(SHA256_result[218]), .A1(n3150), .B0(H1[26]), .B1(n3137), 
        .Y(n565) );
  AOI22XL U458 ( .A0(SHA256_result[155]), .A1(n3147), .B0(H3[27]), .B1(n3138), 
        .Y(n546) );
  AOI22XL U459 ( .A0(SHA256_result[151]), .A1(n3150), .B0(H3[23]), .B1(n3137), 
        .Y(n571) );
  AOI22XL U460 ( .A0(SHA256_result[183]), .A1(n3150), .B0(H2[23]), .B1(n3137), 
        .Y(n568) );
  AOI22XL U461 ( .A0(SHA256_result[137]), .A1(n3145), .B0(H3[9]), .B1(n3137), 
        .Y(n626) );
  AOI22XL U462 ( .A0(SHA256_result[85]), .A1(n3145), .B0(H5[21]), .B1(n3132), 
        .Y(n630) );
  AOI22XL U463 ( .A0(SHA256_result[139]), .A1(n3150), .B0(H3[11]), .B1(n3136), 
        .Y(n583) );
  AOI22XL U464 ( .A0(SHA256_result[90]), .A1(n3150), .B0(H5[26]), .B1(n3136), 
        .Y(n581) );
  AOI22XL U465 ( .A0(SHA256_result[134]), .A1(n3144), .B0(H3[6]), .B1(n3131), 
        .Y(n646) );
  AOI22XL U466 ( .A0(SHA256_result[135]), .A1(n3144), .B0(H3[7]), .B1(n3131), 
        .Y(n645) );
  AOI22XL U467 ( .A0(SHA256_result[149]), .A1(n3144), .B0(H3[21]), .B1(n3131), 
        .Y(n647) );
  BUFX8 U468 ( .A(SHA256_result[119]), .Y(n2909) );
  BUFX8 U469 ( .A(SHA256_result[120]), .Y(n2930) );
  OAI211XL U470 ( .A0(n2980), .A1(n3824), .B0(n3112), .C0(n937), .Y(n2471) );
  INVXL U471 ( .A(SHA256_result[14]), .Y(n3820) );
  AOI22XL U472 ( .A0(N850), .A1(n2942), .B0(SHA256_result[215]), .B1(n3157), 
        .Y(n469) );
  AOI22XL U473 ( .A0(N1009), .A1(n2938), .B0(SHA256_result[54]), .B1(n3161), 
        .Y(n527) );
  OAI211XL U474 ( .A0(n2980), .A1(n3840), .B0(n3112), .C0(n934), .Y(n2479) );
  INVXL U475 ( .A(SHA256_result[205]), .Y(n3545) );
  INVXL U476 ( .A(SHA256_result[207]), .Y(n3538) );
  NAND3BXL U477 ( .AN(n3523), .B(n3108), .C(n3522), .Y(n2831) );
  OAI211XL U478 ( .A0(n2978), .A1(n3830), .B0(n3109), .C0(n752), .Y(n2790) );
  OAI211XL U479 ( .A0(n2980), .A1(n3839), .B0(n3112), .C0(n936), .Y(n2475) );
  OAI211XL U480 ( .A0(n2980), .A1(n3838), .B0(n3112), .C0(n935), .Y(n2476) );
  OAI211XL U481 ( .A0(n2977), .A1(n3813), .B0(n3110), .C0(n767), .Y(n2765) );
  OAI211XL U482 ( .A0(n2977), .A1(n3833), .B0(n3109), .C0(n749), .Y(n2794) );
  AOI22XL U483 ( .A0(N871), .A1(n2940), .B0(SHA256_result[204]), .B1(n3031), 
        .Y(n754) );
  INVXL U484 ( .A(SHA256_result[173]), .Y(n3546) );
  AOI22XL U485 ( .A0(N872), .A1(n2940), .B0(SHA256_result[205]), .B1(n3031), 
        .Y(n755) );
  OAI211XL U486 ( .A0(n2981), .A1(n3812), .B0(n3112), .C0(n941), .Y(n2464) );
  INVXL U487 ( .A(SHA256_result[15]), .Y(n3812) );
  AOI22XL U488 ( .A0(N1034), .A1(n2937), .B0(SHA256_result[47]), .B1(n3027), 
        .Y(n941) );
  OAI211XL U489 ( .A0(n2981), .A1(n3809), .B0(n3112), .C0(n926), .Y(n2495) );
  AOI22XL U490 ( .A0(N1003), .A1(n2936), .B0(n3034), .B1(SHA256_result[80]), 
        .Y(n926) );
  AOI22XL U491 ( .A0(N906), .A1(n2942), .B0(SHA256_result[175]), .B1(n3030), 
        .Y(n776) );
  AOI22XL U492 ( .A0(N908), .A1(n2966), .B0(SHA256_result[177]), .B1(n3029), 
        .Y(n778) );
  AOI22XL U493 ( .A0(N907), .A1(n2973), .B0(SHA256_result[176]), .B1(n3029), 
        .Y(n777) );
  AOI22XL U494 ( .A0(N910), .A1(n2974), .B0(SHA256_result[179]), .B1(n3029), 
        .Y(n780) );
  AOI22XL U495 ( .A0(N909), .A1(n2967), .B0(SHA256_result[178]), .B1(n3029), 
        .Y(n779) );
  OAI211XL U496 ( .A0(n2976), .A1(n3540), .B0(n3110), .C0(n757), .Y(n2783) );
  INVXL U497 ( .A(SHA256_result[175]), .Y(n3540) );
  AOI22XL U498 ( .A0(N874), .A1(n2940), .B0(SHA256_result[207]), .B1(n3031), 
        .Y(n757) );
  AOI22XL U499 ( .A0(N876), .A1(n2940), .B0(SHA256_result[209]), .B1(n3031), 
        .Y(n758) );
  AOI22XL U500 ( .A0(N873), .A1(n2940), .B0(SHA256_result[206]), .B1(n3031), 
        .Y(n756) );
  AOI22XL U501 ( .A0(N877), .A1(n2940), .B0(SHA256_result[210]), .B1(n3031), 
        .Y(n759) );
  AOI22XL U502 ( .A0(N878), .A1(n2940), .B0(SHA256_result[211]), .B1(n3031), 
        .Y(n760) );
  AOI22XL U503 ( .A0(N905), .A1(n2941), .B0(SHA256_result[174]), .B1(n3030), 
        .Y(n775) );
  AOI22XL U504 ( .A0(N904), .A1(n2941), .B0(SHA256_result[173]), .B1(n3030), 
        .Y(n774) );
  AOI22XL U505 ( .A0(N903), .A1(n2941), .B0(SHA256_result[172]), .B1(n3030), 
        .Y(n773) );
  OAI211XL U506 ( .A0(n2979), .A1(n3802), .B0(n3110), .C0(n770), .Y(n2761) );
  OAI211XL U507 ( .A0(n1154), .A1(n2982), .B0(n3111), .C0(n823), .Y(n2688) );
  NAND3BXL U508 ( .AN(n3175), .B(n3112), .C(n3174), .Y(n2829) );
  NAND3BXL U509 ( .AN(n3181), .B(n3112), .C(n3180), .Y(n2510) );
  NAND3BXL U510 ( .AN(n3242), .B(n3112), .C(n3241), .Y(n2506) );
  NAND3BXL U511 ( .AN(n3280), .B(n3112), .C(n3279), .Y(n2508) );
  NAND3BXL U512 ( .AN(n3307), .B(n3112), .C(n3306), .Y(n2503) );
  NAND3BXL U513 ( .AN(n3314), .B(n3112), .C(n3313), .Y(n2700) );
  OAI211XL U514 ( .A0(n1152), .A1(n2982), .B0(n3111), .C0(n824), .Y(n2686) );
  AOI22XL U515 ( .A0(N875), .A1(n2938), .B0(SHA256_result[176]), .B1(n3157), 
        .Y(n518) );
  AOI22XL U516 ( .A0(N1035), .A1(n2942), .B0(SHA256_result[16]), .B1(n3156), 
        .Y(n504) );
  AOI22XL U517 ( .A0(N1036), .A1(n2944), .B0(SHA256_result[17]), .B1(n3156), 
        .Y(n503) );
  AOI22XL U518 ( .A0(N1005), .A1(n2971), .B0(SHA256_result[50]), .B1(n3157), 
        .Y(n531) );
  AOI22XL U519 ( .A0(N897), .A1(n2944), .B0(SHA256_result[134]), .B1(n3156), 
        .Y(n490) );
  AOI22XL U520 ( .A0(N974), .A1(n2942), .B0(SHA256_result[83]), .B1(n3161), 
        .Y(n454) );
  INVXL U521 ( .A(SHA256_result[50]), .Y(n3798) );
  AOI22XL U522 ( .A0(N1037), .A1(n2943), .B0(SHA256_result[18]), .B1(n3156), 
        .Y(n502) );
  AOI22XL U523 ( .A0(N898), .A1(n2943), .B0(SHA256_result[135]), .B1(n3157), 
        .Y(n489) );
  AOI22XL U524 ( .A0(N902), .A1(n2942), .B0(SHA256_result[139]), .B1(n3157), 
        .Y(n487) );
  AOI22XL U525 ( .A0(N911), .A1(n2943), .B0(SHA256_result[148]), .B1(n3159), 
        .Y(n486) );
  AOI22XL U526 ( .A0(N975), .A1(n2942), .B0(SHA256_result[84]), .B1(n3161), 
        .Y(n453) );
  AOI22XL U527 ( .A0(N1039), .A1(n2944), .B0(SHA256_result[20]), .B1(n3156), 
        .Y(n500) );
  INVXL U528 ( .A(SHA256_result[51]), .Y(n3796) );
  AOI22XL U529 ( .A0(N1038), .A1(n2944), .B0(SHA256_result[19]), .B1(n3156), 
        .Y(n501) );
  AOI22XL U530 ( .A0(N1006), .A1(n2965), .B0(SHA256_result[51]), .B1(n3161), 
        .Y(n530) );
  AOI22XL U531 ( .A0(N879), .A1(n2938), .B0(SHA256_result[180]), .B1(n3157), 
        .Y(n517) );
  AOI22XL U532 ( .A0(N1007), .A1(n2972), .B0(SHA256_result[52]), .B1(n3157), 
        .Y(n529) );
  NAND2XL U533 ( .A(n3137), .B(H5[7]), .Y(n3502) );
  AOI22XL U534 ( .A0(n3099), .A1(SHA256_result[140]), .B0(n1092), .B1(
        SHA256_result[172]), .Y(n1186) );
  AOI22XL U535 ( .A0(n3099), .A1(SHA256_result[141]), .B0(n1092), .B1(
        SHA256_result[173]), .Y(n1182) );
  AOI22XL U536 ( .A0(n3099), .A1(SHA256_result[142]), .B0(n1092), .B1(
        SHA256_result[174]), .Y(n1178) );
  AOI22XL U537 ( .A0(n3099), .A1(SHA256_result[143]), .B0(n1092), .B1(
        SHA256_result[175]), .Y(n1174) );
  AOI22XL U538 ( .A0(n3103), .A1(SHA256_result[15]), .B0(n3101), .B1(
        SHA256_result[47]), .Y(n1175) );
  AOI22XL U539 ( .A0(n3103), .A1(SHA256_result[16]), .B0(n3101), .B1(
        SHA256_result[48]), .Y(n1171) );
  AOI22XL U540 ( .A0(n3103), .A1(SHA256_result[17]), .B0(n3101), .B1(
        SHA256_result[49]), .Y(n1164) );
  AOI22XL U541 ( .A0(n3103), .A1(SHA256_result[18]), .B0(n3101), .B1(
        SHA256_result[50]), .Y(n1155) );
  AOI22XL U542 ( .A0(n3103), .A1(SHA256_result[19]), .B0(n3101), .B1(
        SHA256_result[51]), .Y(n1147) );
  OAI21XL U543 ( .A0(SHA256_result[172]), .A1(SHA256_result[204]), .B0(
        SHA256_result[236]), .Y(n3220) );
  OAI2BB1X1 U544 ( .A0N(SHA256_result[173]), .A1N(SHA256_result[205]), .B0(
        n3219), .Y(f2_ABC_32[13]) );
  NAND3X1 U545 ( .A(n2767), .B(n3177), .C(n3176), .Y(n1635) );
  OR2XL U546 ( .A(n3065), .B(n3182), .Y(n2767) );
  NAND3X1 U547 ( .A(n2768), .B(n3492), .C(n3491), .Y(n1595) );
  OR2XL U548 ( .A(n3070), .B(n3490), .Y(n2768) );
  NAND3X1 U549 ( .A(n2773), .B(n3424), .C(n3423), .Y(n1605) );
  OR2XL U550 ( .A(n3067), .B(n3422), .Y(n2773) );
  NAND3X1 U551 ( .A(n2774), .B(n3427), .C(n3426), .Y(n1632) );
  OR2XL U552 ( .A(n3069), .B(n3425), .Y(n2774) );
  NAND3X1 U553 ( .A(n2775), .B(n3256), .C(n3255), .Y(n1633) );
  OR2XL U554 ( .A(n3070), .B(n3254), .Y(n2775) );
  NAND3X1 U555 ( .A(n2778), .B(n3304), .C(n3303), .Y(n1606) );
  OR2XL U556 ( .A(n3067), .B(n3302), .Y(n2778) );
  NAND3X1 U557 ( .A(n2782), .B(n3317), .C(n3316), .Y(n1610) );
  OR2XL U558 ( .A(n3065), .B(n3315), .Y(n2782) );
  NAND3X1 U559 ( .A(n2787), .B(n3320), .C(n3319), .Y(n1608) );
  OR2XL U560 ( .A(n3066), .B(n3318), .Y(n2787) );
  NAND3X1 U561 ( .A(n2788), .B(n3323), .C(n3322), .Y(n1607) );
  OR2XL U562 ( .A(n3068), .B(n3321), .Y(n2788) );
  NAND3X1 U563 ( .A(n2791), .B(n3326), .C(n3325), .Y(n1609) );
  OR2XL U564 ( .A(n3066), .B(n3324), .Y(n2791) );
  NOR2XL U565 ( .A(n3071), .B(n3486), .Y(n3489) );
  NAND2XL U566 ( .A(SHA256_result[206]), .B(n3160), .Y(n3487) );
  NAND3X1 U567 ( .A(n2795), .B(n3506), .C(n3505), .Y(n1574) );
  OR2XL U568 ( .A(n3069), .B(n3504), .Y(n2795) );
  AOI22XL U569 ( .A0(N839), .A1(n2942), .B0(SHA256_result[204]), .B1(n3161), 
        .Y(n473) );
  AOI22XL U570 ( .A0(N847), .A1(n2943), .B0(SHA256_result[212]), .B1(n3156), 
        .Y(n470) );
  AOI22XL U571 ( .A0(N1008), .A1(n2938), .B0(SHA256_result[53]), .B1(n3157), 
        .Y(n528) );
  INVX1 U572 ( .A(n3066), .Y(n3038) );
  INVX1 U573 ( .A(n3071), .Y(n3033) );
  INVX1 U574 ( .A(n3073), .Y(n3034) );
  INVX1 U575 ( .A(n3072), .Y(n3031) );
  INVX1 U576 ( .A(n3070), .Y(n3030) );
  INVX1 U577 ( .A(n3072), .Y(n3032) );
  INVX1 U578 ( .A(n3073), .Y(n3035) );
  INVX1 U579 ( .A(n3069), .Y(n3036) );
  INVX1 U580 ( .A(n3072), .Y(n3028) );
  INVX1 U581 ( .A(n3088), .Y(n3040) );
  INVX1 U582 ( .A(n3024), .Y(n3065) );
  INVX1 U583 ( .A(n3077), .Y(n3067) );
  INVX1 U584 ( .A(n3077), .Y(n3066) );
  INVX1 U585 ( .A(n3084), .Y(n3047) );
  INVX1 U586 ( .A(n3085), .Y(n3046) );
  INVX1 U587 ( .A(n3083), .Y(n3049) );
  INVX1 U588 ( .A(n3087), .Y(n3042) );
  INVX1 U589 ( .A(n3087), .Y(n3041) );
  INVX1 U590 ( .A(n3084), .Y(n3048) );
  INVX1 U591 ( .A(n3086), .Y(n3044) );
  INVX1 U592 ( .A(n3085), .Y(n3045) );
  INVX1 U593 ( .A(n3086), .Y(n3043) );
  INVX1 U594 ( .A(n3083), .Y(n3050) );
  INVX1 U595 ( .A(n3088), .Y(n3039) );
  INVX1 U596 ( .A(n3079), .Y(n3057) );
  INVX1 U597 ( .A(n2992), .Y(n2979) );
  INVX1 U598 ( .A(n2992), .Y(n2977) );
  INVX1 U599 ( .A(n2993), .Y(n2981) );
  INVX1 U600 ( .A(n2991), .Y(n2978) );
  INVX1 U601 ( .A(n2993), .Y(n2980) );
  INVX1 U602 ( .A(n2991), .Y(n2976) );
  INVX1 U603 ( .A(n3080), .Y(n3059) );
  INVX1 U604 ( .A(n3080), .Y(n3058) );
  INVX1 U605 ( .A(n3080), .Y(n3056) );
  INVX1 U606 ( .A(n3079), .Y(n3060) );
  INVX1 U607 ( .A(n3081), .Y(n3055) );
  INVX1 U608 ( .A(n3081), .Y(n3054) );
  INVX1 U609 ( .A(n3082), .Y(n3053) );
  INVX1 U610 ( .A(n3082), .Y(n3052) );
  INVX1 U611 ( .A(n3082), .Y(n3051) );
  INVX1 U612 ( .A(n3078), .Y(n3061) );
  INVX1 U613 ( .A(n3078), .Y(n3063) );
  INVX1 U614 ( .A(n3078), .Y(n3062) );
  INVX1 U615 ( .A(n2711), .Y(n3720) );
  NOR2X1 U616 ( .A(n3746), .B(n3716), .Y(n1249) );
  INVX1 U617 ( .A(n1251), .Y(n3708) );
  INVX1 U618 ( .A(n2954), .Y(n2940) );
  INVX1 U619 ( .A(n2956), .Y(n2941) );
  INVX1 U620 ( .A(n2953), .Y(n2935) );
  INVX1 U621 ( .A(n2956), .Y(n2938) );
  INVX1 U622 ( .A(n2958), .Y(n2943) );
  INVX1 U623 ( .A(n2957), .Y(n2942) );
  INVX1 U624 ( .A(n2952), .Y(n2939) );
  INVX1 U625 ( .A(n2958), .Y(n2944) );
  INVX1 U626 ( .A(n2955), .Y(n2936) );
  INVX1 U627 ( .A(n3074), .Y(n3072) );
  INVX1 U628 ( .A(n3020), .Y(n3079) );
  INVX1 U629 ( .A(n3022), .Y(n3087) );
  INVX1 U630 ( .A(n3021), .Y(n3084) );
  INVX1 U631 ( .A(n3021), .Y(n3085) );
  INVX1 U632 ( .A(n3022), .Y(n3086) );
  INVX1 U633 ( .A(n3021), .Y(n3083) );
  INVX1 U634 ( .A(n3022), .Y(n3088) );
  NOR2X1 U635 ( .A(n3739), .B(n3719), .Y(n1274) );
  INVX1 U636 ( .A(n2397), .Y(n3097) );
  INVX1 U637 ( .A(n2952), .Y(n2947) );
  INVX1 U638 ( .A(n2999), .Y(n2984) );
  INVX1 U639 ( .A(n2999), .Y(n2983) );
  INVX1 U640 ( .A(n2998), .Y(n2985) );
  INVX1 U641 ( .A(n2998), .Y(n2986) );
  INVX1 U642 ( .A(n2998), .Y(n2987) );
  INVX1 U643 ( .A(n2999), .Y(n2988) );
  INVX1 U644 ( .A(n2997), .Y(n2989) );
  INVX1 U645 ( .A(n2997), .Y(n2990) );
  INVX1 U646 ( .A(n3020), .Y(n3080) );
  INVX1 U647 ( .A(n3020), .Y(n3078) );
  INVX1 U648 ( .A(n3020), .Y(n3081) );
  INVX1 U649 ( .A(n3020), .Y(n3082) );
  INVX1 U650 ( .A(n2996), .Y(n2991) );
  INVX1 U651 ( .A(n1401), .Y(n3746) );
  INVX1 U652 ( .A(n1324), .Y(n3759) );
  INVX1 U653 ( .A(n1374), .Y(n3734) );
  INVX1 U654 ( .A(n1467), .Y(n3763) );
  INVX1 U655 ( .A(n1307), .Y(n3758) );
  INVX1 U656 ( .A(n1287), .Y(n3739) );
  INVX1 U657 ( .A(n1352), .Y(n3733) );
  NAND2X1 U658 ( .A(n3746), .B(n3741), .Y(n1413) );
  INVX1 U659 ( .A(n3015), .Y(n3012) );
  INVX1 U660 ( .A(n3016), .Y(n3004) );
  INVX1 U661 ( .A(n2825), .Y(n3013) );
  INVX1 U662 ( .A(n2714), .Y(n3716) );
  INVX1 U663 ( .A(n1382), .Y(n3711) );
  NOR2X1 U664 ( .A(n3764), .B(n3709), .Y(n1251) );
  INVX1 U665 ( .A(n3014), .Y(n3010) );
  INVX1 U666 ( .A(n3014), .Y(n3011) );
  INVX1 U667 ( .A(n3017), .Y(n3005) );
  INVX1 U668 ( .A(n3017), .Y(n3002) );
  INVX1 U669 ( .A(n3015), .Y(n3009) );
  INVX1 U670 ( .A(n3015), .Y(n3008) );
  INVX1 U671 ( .A(n1424), .Y(n3712) );
  INVX1 U672 ( .A(n2970), .Y(n2953) );
  INVX1 U673 ( .A(n2969), .Y(n2955) );
  INVX1 U674 ( .A(n2969), .Y(n2956) );
  INVX1 U675 ( .A(n2969), .Y(n2957) );
  INVX1 U676 ( .A(n3025), .Y(n3019) );
  INVX1 U677 ( .A(n3023), .Y(n3021) );
  INVX1 U678 ( .A(n3023), .Y(n3022) );
  INVX1 U679 ( .A(n3018), .Y(n3074) );
  INVX1 U680 ( .A(n3018), .Y(n3075) );
  INVX1 U681 ( .A(n3018), .Y(n3076) );
  NOR2X1 U682 ( .A(n1366), .B(n3737), .Y(n1316) );
  NOR2X1 U683 ( .A(n3764), .B(n3089), .Y(n1411) );
  OAI21XL U684 ( .A0(n3089), .A1(n3755), .B0(n3718), .Y(n1412) );
  CLKINVX3 U685 ( .A(n3142), .Y(n3140) );
  CLKINVX3 U686 ( .A(n3142), .Y(n3139) );
  INVX1 U687 ( .A(n2397), .Y(n3096) );
  INVX1 U688 ( .A(n3142), .Y(n3133) );
  INVX1 U689 ( .A(n3143), .Y(n3135) );
  INVX1 U690 ( .A(n3143), .Y(n3132) );
  INVX1 U691 ( .A(n3143), .Y(n3131) );
  INVX1 U692 ( .A(n3142), .Y(n3136) );
  INVX1 U693 ( .A(n3143), .Y(n3137) );
  INVX1 U694 ( .A(n3142), .Y(n3138) );
  INVX1 U695 ( .A(n3143), .Y(n3134) );
  INVX1 U696 ( .A(n2395), .Y(n3101) );
  INVX1 U697 ( .A(n3095), .Y(n3094) );
  INVX1 U698 ( .A(n3143), .Y(n3141) );
  INVX1 U699 ( .A(n1366), .Y(n3707) );
  INVX1 U700 ( .A(n1242), .Y(n3710) );
  INVX1 U701 ( .A(n2394), .Y(n3103) );
  INVX1 U702 ( .A(n2973), .Y(n2951) );
  INVX1 U703 ( .A(n2973), .Y(n2950) );
  INVX1 U704 ( .A(n2974), .Y(n2949) );
  INVX1 U705 ( .A(n2974), .Y(n2948) );
  INVX1 U706 ( .A(n2967), .Y(n2961) );
  INVX1 U707 ( .A(n2967), .Y(n2962) );
  INVX1 U708 ( .A(n2965), .Y(n2963) );
  INVX1 U709 ( .A(n2965), .Y(n2964) );
  INVX1 U710 ( .A(n3024), .Y(n3020) );
  INVX1 U711 ( .A(n2719), .Y(n2995) );
  NOR2X1 U712 ( .A(n3760), .B(n3776), .Y(n1324) );
  NOR2X1 U713 ( .A(n3760), .B(n3779), .Y(n1307) );
  NOR2X1 U714 ( .A(n3776), .B(n3750), .Y(n1401) );
  INVX1 U715 ( .A(n1306), .Y(n3738) );
  INVX1 U716 ( .A(n2721), .Y(n3775) );
  INVX1 U717 ( .A(n1278), .Y(n3743) );
  NOR2X1 U718 ( .A(n3775), .B(n3737), .Y(n1277) );
  INVX1 U719 ( .A(n1311), .Y(n3761) );
  INVX1 U720 ( .A(n1295), .Y(n3766) );
  INVX1 U721 ( .A(n1351), .Y(n3745) );
  NOR2X1 U722 ( .A(n3745), .B(n3778), .Y(n1303) );
  NOR2X1 U723 ( .A(n3747), .B(n3760), .Y(n1309) );
  NOR2X1 U724 ( .A(n3737), .B(n3778), .Y(n1374) );
  NOR2X1 U725 ( .A(n3753), .B(n3779), .Y(n1379) );
  NOR2X1 U726 ( .A(n3765), .B(n3778), .Y(n1467) );
  NAND2X1 U727 ( .A(n3762), .B(n3760), .Y(n1484) );
  INVX1 U728 ( .A(n1283), .Y(n3756) );
  INVX1 U729 ( .A(n1310), .Y(n3764) );
  NOR2X1 U730 ( .A(n3753), .B(n3776), .Y(n1291) );
  NOR2X1 U731 ( .A(n3753), .B(n3775), .Y(n1399) );
  INVX1 U732 ( .A(n1474), .Y(n3755) );
  NAND2X1 U733 ( .A(n3753), .B(n3737), .Y(n1246) );
  INVX1 U734 ( .A(n1390), .Y(n3728) );
  OR2X2 U735 ( .A(n3745), .B(n3776), .Y(n2796) );
  INVX1 U736 ( .A(n2796), .Y(n1334) );
  INVX1 U737 ( .A(n1294), .Y(n3741) );
  INVX1 U738 ( .A(n1377), .Y(n3752) );
  NOR2X1 U739 ( .A(n3748), .B(n1309), .Y(n1376) );
  INVX1 U740 ( .A(n1266), .Y(n3747) );
  NOR2X1 U741 ( .A(n3737), .B(n3755), .Y(n1352) );
  OAI21XL U742 ( .A0(n3779), .A1(n3750), .B0(n3734), .Y(n1455) );
  AOI21X1 U743 ( .A0(n1403), .A1(n1484), .B0(n1309), .Y(n1544) );
  OAI21XL U744 ( .A0(n3778), .A1(n3753), .B0(n3729), .Y(n1496) );
  OAI21XL U745 ( .A0(n3745), .A1(n3775), .B0(n3736), .Y(n1315) );
  NOR2X1 U746 ( .A(n3745), .B(n3779), .Y(n1287) );
  INVX1 U747 ( .A(n1365), .Y(n3735) );
  INVX1 U748 ( .A(n1321), .Y(n3729) );
  NAND2X1 U749 ( .A(n3770), .B(n1319), .Y(n1259) );
  NAND2X1 U750 ( .A(n3770), .B(n1278), .Y(n1276) );
  NAND2X1 U751 ( .A(n3736), .B(n3770), .Y(n1438) );
  INVX1 U752 ( .A(n1280), .Y(n3768) );
  INVX1 U753 ( .A(n1372), .Y(n3754) );
  INVX1 U754 ( .A(n3155), .Y(n3144) );
  INVX1 U755 ( .A(n3154), .Y(n3147) );
  INVX1 U756 ( .A(n3154), .Y(n3146) );
  INVX1 U757 ( .A(n3155), .Y(n3145) );
  INVX1 U758 ( .A(n3153), .Y(n3149) );
  INVX1 U759 ( .A(n3153), .Y(n3148) );
  INVX1 U760 ( .A(n3127), .Y(n3116) );
  INVX1 U761 ( .A(n3127), .Y(n3117) );
  INVX1 U762 ( .A(n3129), .Y(n3124) );
  INVX1 U763 ( .A(n3130), .Y(n3122) );
  INVX1 U764 ( .A(n3130), .Y(n3126) );
  INVX1 U765 ( .A(n3127), .Y(n3118) );
  INVX1 U766 ( .A(n3129), .Y(n3123) );
  OAI222XL U767 ( .A0(n3737), .A1(n3714), .B0(n3716), .B1(n1278), .C0(n2389), 
        .C1(n3709), .Y(n1497) );
  OAI221XL U768 ( .A0(n3720), .A1(n3769), .B0(n2817), .B1(n3729), .C0(n1441), 
        .Y(N2960) );
  INVX1 U769 ( .A(n1340), .Y(n3769) );
  AOI222X1 U770 ( .A0(n1442), .A1(n1443), .B0(n3707), .B1(n1444), .C0(n3090), 
        .C1(n1445), .Y(n1441) );
  NAND2X1 U771 ( .A(n3750), .B(n3742), .Y(n1444) );
  OAI221XL U772 ( .A0(n2817), .A1(n3740), .B0(n3716), .B1(n1290), .C0(n1299), 
        .Y(N2973) );
  AOI211X1 U773 ( .A0(n3090), .A1(n1300), .B0(n1301), .C0(n1302), .Y(n1299) );
  NAND4BXL U774 ( .AN(n1303), .B(n3728), .C(n1304), .D(n1305), .Y(n1300) );
  AOI211XL U775 ( .A0(n1399), .A1(n1250), .B0(n1342), .C0(n1249), .Y(n1453) );
  AOI211X1 U776 ( .A0(n1443), .A1(n2721), .B0(n1481), .C0(n1482), .Y(n1480) );
  INVXL U777 ( .A(n2755), .Y(n3714) );
  NAND4X1 U778 ( .A(n1477), .B(n1478), .C(n1479), .D(n1480), .Y(N2956) );
  AOI22XL U779 ( .A0(n2755), .A1(n1401), .B0(n1324), .B1(n2757), .Y(n1477) );
  NAND4X1 U780 ( .A(n1433), .B(n1435), .C(n1436), .D(n1437), .Y(N2961) );
  AOI22X1 U781 ( .A0(n2766), .A1(n1439), .B0(n1411), .B1(n1351), .Y(n1436) );
  NAND4X1 U782 ( .A(n1404), .B(n1405), .C(n1406), .D(n1407), .Y(N2964) );
  OAI21XL U783 ( .A0(n1323), .A1(n1280), .B0(n3707), .Y(n1405) );
  OAI21XL U784 ( .A0(n1379), .A1(n1281), .B0(n2755), .Y(n1404) );
  NAND4BXL U785 ( .AN(n1468), .B(n1469), .C(n1470), .D(n1471), .Y(N2957) );
  AOI22XL U786 ( .A0(n2755), .A1(n1263), .B0(n1475), .B1(n2712), .Y(n1469) );
  NAND2X1 U787 ( .A(n1419), .B(n2721), .Y(n1424) );
  INVX1 U788 ( .A(n3115), .Y(n3108) );
  CLKINVX3 U789 ( .A(n3113), .Y(n3110) );
  CLKINVX3 U790 ( .A(n3115), .Y(n3112) );
  CLKINVX3 U791 ( .A(n3113), .Y(n3111) );
  CLKINVX3 U792 ( .A(n3113), .Y(n3109) );
  INVX1 U793 ( .A(n3162), .Y(n3160) );
  INVX1 U794 ( .A(n3163), .Y(n3159) );
  INVX1 U795 ( .A(n3162), .Y(n3158) );
  INVX1 U796 ( .A(n3163), .Y(n3156) );
  NAND3X1 U797 ( .A(n1325), .B(n1326), .C(n1327), .Y(N2971) );
  AOI22XL U798 ( .A0(n1336), .A1(n996), .B0(n1337), .B1(n2755), .Y(n1325) );
  AOI211X1 U799 ( .A0(n1260), .A1(n2713), .B0(n1328), .C0(n1329), .Y(n1327) );
  NAND3X1 U800 ( .A(n1414), .B(n1415), .C(n1416), .Y(N2963) );
  AOI31X1 U801 ( .A0(n3091), .A1(n996), .A2(n3756), .B0(n1421), .Y(n1415) );
  NAND3X1 U802 ( .A(n1367), .B(n1368), .C(n1369), .Y(N2967) );
  AOI22XL U803 ( .A0(n1250), .A1(n1378), .B0(n1379), .B1(n2718), .Y(n1368) );
  AOI22X1 U804 ( .A0(n1380), .A1(n2713), .B0(n1356), .B1(n2391), .Y(n1367) );
  NAND2X1 U805 ( .A(n1506), .B(n3708), .Y(n1505) );
  NOR3X1 U806 ( .A(n1366), .B(n3777), .C(n2391), .Y(n1357) );
  OAI222XL U807 ( .A0(n1360), .A1(n3089), .B0(n1361), .B1(n3717), .C0(n3720), 
        .C1(n3741), .Y(n1359) );
  AOI21X1 U808 ( .A0(n3775), .A1(n1351), .B0(n1403), .Y(n1476) );
  INVX1 U809 ( .A(n1418), .Y(n3713) );
  INVX1 U810 ( .A(n3162), .Y(n3161) );
  INVX1 U811 ( .A(n2764), .Y(n2970) );
  INVX1 U812 ( .A(n2764), .Y(n2969) );
  INVX1 U813 ( .A(n2764), .Y(n2968) );
  INVX1 U814 ( .A(n3001), .Y(n3017) );
  INVX1 U815 ( .A(n3001), .Y(n3016) );
  OAI221XL U816 ( .A0(n3709), .A1(n1283), .B0(n2817), .B1(n1284), .C0(n1285), 
        .Y(N2974) );
  NAND3BX1 U817 ( .AN(n1277), .B(n3742), .C(n1290), .Y(n1289) );
  NAND4BXL U818 ( .AN(n1291), .B(n3733), .C(n1292), .D(n1293), .Y(n1286) );
  INVX1 U819 ( .A(n1408), .Y(n3770) );
  OAI221XL U820 ( .A0(n3716), .A1(n3730), .B0(n3717), .B1(n3736), .C0(n1540), 
        .Y(N2947) );
  INVX1 U821 ( .A(n1475), .Y(n3730) );
  NAND4BXL U822 ( .AN(n1543), .B(n1278), .C(n3742), .D(n1544), .Y(n1541) );
  AOI31X1 U823 ( .A0(n3758), .A1(n1244), .A2(n1319), .B0(n3089), .Y(n1318) );
  INVX1 U824 ( .A(n1384), .Y(n3779) );
  NAND2X1 U825 ( .A(n1389), .B(n3091), .Y(n1366) );
  OAI211X1 U826 ( .A0(n1238), .A1(n3777), .B0(n1239), .C0(n1240), .Y(N2977) );
  AOI21X1 U827 ( .A0(n3091), .A1(n1241), .B0(n3710), .Y(n1240) );
  AOI21XL U828 ( .A0(n1250), .A1(n1246), .B0(n1251), .Y(n1238) );
  AOI21X1 U829 ( .A0(n1474), .A1(n2757), .B0(n1336), .Y(n1242) );
  AOI31X1 U830 ( .A0(n1371), .A1(n1372), .A2(n1373), .B0(n3089), .Y(n1370) );
  AOI22X1 U831 ( .A0(n1377), .A1(n2766), .B0(n1365), .B1(n996), .Y(n1371) );
  AOI211X1 U832 ( .A0(n1334), .A1(n3762), .B0(n1374), .C0(n1375), .Y(n1373) );
  AOI21X1 U833 ( .A0(n1376), .A1(n3738), .B0(n996), .Y(n1375) );
  AOI31X1 U834 ( .A0(n1397), .A1(n1349), .A2(n1398), .B0(n3089), .Y(n1396) );
  AOI31X1 U835 ( .A0(n3765), .A1(n3778), .A2(n1308), .B0(n1402), .Y(n1397) );
  NOR3X1 U836 ( .A(n3757), .B(n1303), .C(n1399), .Y(n1398) );
  AOI2BB1X1 U837 ( .A0N(n1353), .A1N(n1380), .B0(n3764), .Y(n1402) );
  OAI211X1 U838 ( .A0(n2388), .A1(n1283), .B0(n3733), .C0(n1499), .Y(n1527) );
  AND2X2 U839 ( .A(n972), .B(n2388), .Y(n2798) );
  NAND4X1 U840 ( .A(n1534), .B(n1242), .C(n1535), .D(n1536), .Y(N2948) );
  OAI31XL U841 ( .A0(n1294), .A1(n1374), .A2(n1420), .B0(n2755), .Y(n1536) );
  NAND4X1 U842 ( .A(n1270), .B(n1271), .C(n1272), .D(n1273), .Y(N2975) );
  AOI22XL U843 ( .A0(n3090), .A1(n1279), .B0(n1280), .B1(n1250), .Y(n1271) );
  NAND4X1 U844 ( .A(n1521), .B(n1522), .C(n1523), .D(n1524), .Y(N2950) );
  AOI22XL U845 ( .A0(n3744), .A1(n2755), .B0(n1263), .B1(n2711), .Y(n1521) );
  AOI22XL U846 ( .A0(n1250), .A1(n1525), .B0(n2757), .B1(n1492), .Y(n1524) );
  AOI21X1 U847 ( .A0(n1465), .A1(n1466), .B0(n3089), .Y(n1464) );
  OAI21XL U848 ( .A0(n1467), .A1(n1324), .B0(n1308), .Y(n1466) );
  NAND4X1 U849 ( .A(n1545), .B(n1506), .C(n1546), .D(n1547), .Y(N2946) );
  OAI21XL U850 ( .A0(n1291), .A1(n1303), .B0(n2755), .Y(n1546) );
  NAND3XL U851 ( .A(n2766), .B(n1296), .C(n1250), .Y(n1545) );
  AOI22XL U852 ( .A0(n1295), .A1(n2757), .B0(n3090), .B1(n1548), .Y(n1547) );
  NAND4X1 U853 ( .A(n1252), .B(n1253), .C(n1254), .D(n1255), .Y(N2976) );
  AOI22XL U854 ( .A0(n3757), .A1(n2757), .B0(n2713), .B1(n2766), .Y(n1252) );
  AOI22XL U855 ( .A0(n1250), .A1(n1256), .B0(n3091), .B1(n1257), .Y(n1255) );
  OAI21XL U856 ( .A0(n1379), .A1(n3748), .B0(n1250), .Y(n1423) );
  OAI21XL U857 ( .A0(n1432), .A1(n1316), .B0(n996), .Y(n1425) );
  NAND4X1 U858 ( .A(n1528), .B(n1529), .C(n1530), .D(n1531), .Y(N2949) );
  OAI21XL U859 ( .A0(n1525), .A1(n1386), .B0(n2712), .Y(n1528) );
  AOI22XL U860 ( .A0(n2755), .A1(n1323), .B0(n3091), .B1(n1532), .Y(n1530) );
  AOI21X1 U861 ( .A0(n1281), .A1(n2712), .B0(n1282), .Y(n1270) );
  NAND4BXL U862 ( .AN(n1316), .B(n1392), .C(n1393), .D(n1394), .Y(N2965) );
  OAI21XL U863 ( .A0(n1281), .A1(n1337), .B0(n2718), .Y(n1392) );
  NAND2XL U864 ( .A(n1403), .B(n1250), .Y(n1393) );
  NAND4BXL U865 ( .AN(n1509), .B(n1510), .C(n1511), .D(n1512), .Y(N2952) );
  AOI31X1 U866 ( .A0(n1457), .A1(n3758), .A2(n1513), .B0(n3089), .Y(n1509) );
  OAI21XL U867 ( .A0(n1454), .A1(n1281), .B0(n1250), .Y(n1510) );
  AOI2BB2X1 U868 ( .B0(n1263), .B1(n2711), .A0N(n3716), .A1N(n1361), .Y(n1511)
         );
  NAND4BXL U869 ( .AN(n1282), .B(n1312), .C(n1313), .D(n1314), .Y(N2972) );
  AOI22X1 U870 ( .A0(n1321), .A1(n2714), .B0(n3707), .B1(n2721), .Y(n1312) );
  AOI21XL U871 ( .A0(n2755), .A1(n1315), .B0(n1316), .Y(n1314) );
  INVX1 U872 ( .A(n2393), .Y(n3099) );
  INVX1 U873 ( .A(n2394), .Y(n3102) );
  INVX1 U874 ( .A(n3095), .Y(n3093) );
  INVX1 U875 ( .A(n1094), .Y(n3095) );
  INVX1 U876 ( .A(n2392), .Y(n3105) );
  INVX1 U877 ( .A(n2395), .Y(n3100) );
  NAND3X1 U878 ( .A(n1485), .B(n1486), .C(n1487), .Y(N2955) );
  OAI21XL U880 ( .A0(n1281), .A1(n1335), .B0(n2711), .Y(n1486) );
  AOI31XL U881 ( .A0(n2757), .A1(n2390), .A2(n1364), .B0(n1336), .Y(n1485) );
  INVX1 U882 ( .A(n3092), .Y(n3089) );
  INVX1 U883 ( .A(n2396), .Y(n3107) );
  INVXL U884 ( .A(n495), .Y(n3143) );
  INVXL U885 ( .A(n495), .Y(n3142) );
  NOR2X1 U886 ( .A(n2391), .B(n2388), .Y(n1351) );
  INVX1 U887 ( .A(n1354), .Y(n3776) );
  NOR2X1 U888 ( .A(n3766), .B(n2388), .Y(n1390) );
  INVX1 U889 ( .A(n1491), .Y(n3762) );
  NOR2X1 U890 ( .A(n2389), .B(n2398), .Y(n1389) );
  NOR3X1 U891 ( .A(n2391), .B(n996), .C(n3762), .Y(n1311) );
  INVX1 U892 ( .A(n1457), .Y(n3757) );
  NAND2X1 U893 ( .A(n1400), .B(n2389), .Y(n1278) );
  NOR2X1 U894 ( .A(n3775), .B(n2398), .Y(n1295) );
  NOR2X1 U895 ( .A(n3745), .B(n3777), .Y(n1400) );
  OAI211X1 U896 ( .A0(n2391), .A1(n3764), .B0(n1349), .C0(n1350), .Y(n1348) );
  AOI211X1 U897 ( .A0(n2721), .A1(n1351), .B0(n972), .C0(n1352), .Y(n1350) );
  INVX1 U898 ( .A(n972), .Y(n3767) );
  NOR2X1 U899 ( .A(n3762), .B(n2388), .Y(n1306) );
  INVX1 U900 ( .A(n1442), .Y(n3727) );
  INVX1 U901 ( .A(n1330), .Y(n3731) );
  INVX1 U902 ( .A(n1353), .Y(n3737) );
  AOI221X1 U903 ( .A0(n1294), .A1(n2389), .B0(n1295), .B1(n1296), .C0(n3731), 
        .Y(n1293) );
  AOI222X1 U904 ( .A0(n1306), .A1(n3777), .B0(n1307), .B1(n1308), .C0(n1309), 
        .C1(n3164), .Y(n1305) );
  NOR2X1 U905 ( .A(n3753), .B(n996), .Y(n1263) );
  NOR2X1 U906 ( .A(n3753), .B(n2390), .Y(n1261) );
  NOR2X1 U907 ( .A(n2391), .B(n3776), .Y(n1386) );
  INVX1 U908 ( .A(n1248), .Y(n3760) );
  NOR2X1 U909 ( .A(n3737), .B(n2398), .Y(n1365) );
  NOR2X1 U910 ( .A(n3775), .B(n2391), .Y(n1280) );
  NOR2X1 U911 ( .A(n2388), .B(n3779), .Y(n1321) );
  NOR2X1 U912 ( .A(n3765), .B(n996), .Y(n1310) );
  OAI211X1 U913 ( .A0(n3779), .A1(n3737), .B0(n1499), .C0(n1500), .Y(n1498) );
  AOI211X1 U914 ( .A0(n1475), .A1(n3756), .B0(n972), .C0(n3757), .Y(n1500) );
  INVX1 U915 ( .A(n1265), .Y(n3742) );
  INVX1 U916 ( .A(n1395), .Y(n3736) );
  NOR2X1 U917 ( .A(n3753), .B(n2398), .Y(n1377) );
  NOR2X1 U918 ( .A(n3745), .B(n996), .Y(n1294) );
  NOR2X1 U919 ( .A(n2391), .B(n3778), .Y(n1403) );
  NOR2X1 U920 ( .A(n2389), .B(n3778), .Y(n1474) );
  INVX1 U921 ( .A(n2766), .Y(n3778) );
  INVX1 U922 ( .A(n1364), .Y(n3765) );
  NOR2X1 U923 ( .A(n3750), .B(n2390), .Y(n1266) );
  INVX1 U924 ( .A(n1391), .Y(n3732) );
  NAND4X1 U925 ( .A(n1243), .B(n3732), .C(n2796), .D(n1244), .Y(n1241) );
  NAND2X1 U926 ( .A(n2721), .B(n1246), .Y(n1243) );
  AOI21X1 U927 ( .A0(n1310), .A1(n1308), .B0(n3756), .Y(n1372) );
  OAI21XL U928 ( .A0(n3765), .A1(n3736), .B0(n1298), .Y(n1431) );
  INVX1 U929 ( .A(n1284), .Y(n3748) );
  AOI21X1 U930 ( .A0(n1384), .A1(n1377), .B0(n1442), .Y(n1499) );
  NAND2X1 U931 ( .A(n1340), .B(n1389), .Y(n1283) );
  NOR2XL U932 ( .A(n1265), .B(n1281), .Y(n1361) );
  OAI21XL U933 ( .A0(n2390), .A1(n3737), .B0(n3739), .Y(n1378) );
  INVX1 U934 ( .A(n1420), .Y(n3751) );
  NAND2X1 U935 ( .A(n1284), .B(n1278), .Y(n1258) );
  AOI21X1 U936 ( .A0(n2766), .A1(n3765), .B0(n1390), .Y(n1388) );
  INVX1 U937 ( .A(n1244), .Y(n3744) );
  INVX1 U938 ( .A(n1335), .Y(n3740) );
  NAND2BX1 U939 ( .AN(n1337), .B(n3779), .Y(n1422) );
  AOI22XL U940 ( .A0(n996), .A1(n1297), .B0(n1281), .B1(n2398), .Y(n1292) );
  NAND2X1 U941 ( .A(n1298), .B(n3752), .Y(n1297) );
  AOI221X1 U942 ( .A0(n2398), .A1(n1400), .B0(n3777), .B1(n1391), .C0(n1401), 
        .Y(n1349) );
  INVX1 U943 ( .A(n1308), .Y(n3753) );
  INVX1 U944 ( .A(n1296), .Y(n3750) );
  OR2X2 U945 ( .A(n1259), .B(n1260), .Y(n1256) );
  NOR2X1 U946 ( .A(n3750), .B(n996), .Y(n1323) );
  NOR2X1 U947 ( .A(n2388), .B(n2390), .Y(n1454) );
  NAND2X1 U948 ( .A(n1353), .B(n1354), .Y(n1319) );
  NAND2X1 U949 ( .A(n3747), .B(n2819), .Y(n1355) );
  XOR3X2 U950 ( .A(n2899), .B(n2682), .C(n2859), .Y(f4_E_32[6]) );
  AOI21X1 U951 ( .A0(n2985), .A1(n2855), .B0(n3114), .Y(n3295) );
  NAND2XL U952 ( .A(n2405), .B(n3036), .Y(n3351) );
  AOI21X1 U953 ( .A0(n2849), .A1(n2984), .B0(n3114), .Y(n3265) );
  NAND2XL U954 ( .A(next_A[29]), .B(n3037), .Y(n3264) );
  AND2X2 U955 ( .A(n2860), .B(n3159), .Y(n2805) );
  NAND2XL U956 ( .A(next_A[31]), .B(n3035), .Y(n3375) );
  AOI21XL U957 ( .A0(n3033), .A1(next_E[31]), .B0(n3396), .Y(n3397) );
  NOR2BX1 U958 ( .AN(n3161), .B(n2683), .Y(n3396) );
  XOR3X2 U959 ( .A(n2924), .B(n2919), .C(n2916), .Y(f3_A_32[4]) );
  XOR3X2 U960 ( .A(SHA256_result[235]), .B(n2901), .C(n2887), .Y(f3_A_32[9])
         );
  XOR3X2 U961 ( .A(n2878), .B(n2884), .C(n2851), .Y(f4_E_32[8]) );
  XOR3X2 U962 ( .A(n2872), .B(n2896), .C(n2844), .Y(f4_E_32[9]) );
  NAND3X1 U963 ( .A(n3301), .B(n3300), .C(n3299), .Y(n2870) );
  NAND3X2 U964 ( .A(n3367), .B(n3366), .C(n3365), .Y(n3557) );
  NAND2X2 U965 ( .A(N949), .B(n2946), .Y(n3367) );
  NAND3X1 U966 ( .A(n3456), .B(n3455), .C(n3454), .Y(n3572) );
  NAND2X1 U967 ( .A(n2916), .B(n3158), .Y(n3454) );
  NAND2XL U968 ( .A(next_A[26]), .B(n3035), .Y(n3455) );
  NAND3X1 U969 ( .A(n3379), .B(n3378), .C(n3377), .Y(n3573) );
  NAND2X1 U970 ( .A(n2888), .B(n3159), .Y(n3377) );
  NAND2XL U971 ( .A(next_A[24]), .B(n3035), .Y(n3378) );
  NAND2X2 U972 ( .A(N819), .B(n2947), .Y(n3379) );
  NAND3X1 U973 ( .A(n3485), .B(n3484), .C(n3483), .Y(n2710) );
  AOI21X1 U974 ( .A0(n2930), .A1(n2987), .B0(n3115), .Y(n3485) );
  NAND2XL U975 ( .A(next_E[24]), .B(n3034), .Y(n3484) );
  NAND2X1 U976 ( .A(N947), .B(n2946), .Y(n3483) );
  NAND3X1 U977 ( .A(n3400), .B(n3399), .C(n3398), .Y(n3574) );
  NAND2XL U978 ( .A(n3035), .B(next_A[23]), .Y(n3399) );
  NAND3X1 U979 ( .A(n3395), .B(n3394), .C(n3393), .Y(n3575) );
  NAND2XL U980 ( .A(n3035), .B(next_A[22]), .Y(n3394) );
  NAND2X2 U981 ( .A(N817), .B(n2945), .Y(n3395) );
  XOR3X2 U982 ( .A(n2877), .B(n2915), .C(SHA256_result[104]), .Y(f4_E_32[15])
         );
  XOR3X2 U983 ( .A(n2928), .B(n2919), .C(n2862), .Y(f3_A_32[15]) );
  XOR3X2 U984 ( .A(n2929), .B(SHA256_result[251]), .C(SHA256_result[240]), .Y(
        f3_A_32[14]) );
  XOR3X2 U985 ( .A(n2933), .B(SHA256_result[236]), .C(n2903), .Y(f3_A_32[10])
         );
  XOR3X2 U986 ( .A(n2857), .B(n2892), .C(SHA256_result[238]), .Y(f3_A_32[12])
         );
  XOR3X2 U987 ( .A(n2905), .B(n2916), .C(SHA256_result[239]), .Y(f3_A_32[13])
         );
  XOR3X2 U988 ( .A(n2930), .B(n2884), .C(n2833), .Y(f4_E_32[13]) );
  XOR3X2 U989 ( .A(SHA256_result[114]), .B(n2909), .C(n2840), .Y(f4_E_32[12])
         );
  XOR3X2 U990 ( .A(n2874), .B(n2909), .C(n2867), .Y(f4_E_32[17]) );
  NAND4X1 U991 ( .A(n3108), .B(n3283), .C(n3282), .D(n3281), .Y(n2882) );
  NAND2X1 U992 ( .A(SHA256_result[237]), .B(n2987), .Y(n3283) );
  NAND2XL U993 ( .A(next_A[13]), .B(n3037), .Y(n3282) );
  XOR3X2 U994 ( .A(SHA256_result[121]), .B(n2896), .C(n2830), .Y(f4_E_32[14])
         );
  OAI2BB1X1 U995 ( .A0N(SHA256_result[236]), .A1N(n3161), .B0(n3405), .Y(n3580) );
  AOI2BB2X1 U996 ( .B0(N807), .B1(n2944), .A0N(n3040), .A1N(n3404), .Y(n3405)
         );
  INVXL U997 ( .A(next_A[12]), .Y(n3404) );
  XOR3X2 U998 ( .A(n2869), .B(n2910), .C(n2864), .Y(f4_E_32[16]) );
  XOR3X2 U999 ( .A(n2930), .B(n2860), .C(n2858), .Y(f4_E_32[18]) );
  XOR3X2 U1000 ( .A(n2888), .B(n2906), .C(SHA256_result[237]), .Y(f3_A_32[11])
         );
  NAND3X1 U1001 ( .A(n3447), .B(n3446), .C(n3445), .Y(n3560) );
  NAND3X1 U1002 ( .A(n3389), .B(n3388), .C(n3387), .Y(n3562) );
  NAND2X1 U1003 ( .A(n3157), .B(n2896), .Y(n3387) );
  NAND2X1 U1004 ( .A(N943), .B(n2946), .Y(n3389) );
  NAND3X1 U1005 ( .A(n3238), .B(n3237), .C(n3236), .Y(n1553) );
  NAND3X1 U1006 ( .A(n3453), .B(n3452), .C(n3451), .Y(n2716) );
  AOI21X1 U1007 ( .A0(SHA256_result[114]), .A1(n2983), .B0(n3114), .Y(n3453)
         );
  NAND2X1 U1008 ( .A(N941), .B(n2946), .Y(n3451) );
  OR3XL U1009 ( .A(n2808), .B(n2811), .C(n2812), .Y(n3559) );
  AND2X2 U1010 ( .A(N946), .B(n2945), .Y(n2808) );
  AND2X1 U1011 ( .A(next_E[23]), .B(n3035), .Y(n2811) );
  AND2X2 U1012 ( .A(n3157), .B(n2909), .Y(n2812) );
  NAND3X1 U1013 ( .A(n3382), .B(n3381), .C(n3380), .Y(n3576) );
  NAND2X1 U1014 ( .A(n2891), .B(n3159), .Y(n3380) );
  NAND2XL U1015 ( .A(next_A[21]), .B(n3035), .Y(n3381) );
  NAND2X1 U1016 ( .A(N816), .B(n2945), .Y(n3382) );
  NAND3X1 U1017 ( .A(n3450), .B(n3449), .C(n3448), .Y(n3561) );
  NAND2X2 U1018 ( .A(N944), .B(n2946), .Y(n3450) );
  NAND3X1 U1019 ( .A(n3286), .B(n3285), .C(n3284), .Y(n2880) );
  AOI21X1 U1020 ( .A0(SHA256_result[239]), .A1(n2984), .B0(n3114), .Y(n3286)
         );
  NAND2XL U1021 ( .A(next_A[15]), .B(n3036), .Y(n3285) );
  NAND2X1 U1022 ( .A(N810), .B(n2945), .Y(n3284) );
  NAND3X1 U1023 ( .A(n3403), .B(n3402), .C(n3401), .Y(n3578) );
  NAND2XL U1024 ( .A(next_A[18]), .B(n3035), .Y(n3402) );
  NAND2X1 U1025 ( .A(N813), .B(n2945), .Y(n3403) );
  NAND3X1 U1026 ( .A(n3373), .B(n3372), .C(n3371), .Y(n2715) );
  AOI21X1 U1027 ( .A0(n2985), .A1(n2884), .B0(n3114), .Y(n3373) );
  NAND2X1 U1028 ( .A(next_E[19]), .B(n3036), .Y(n3372) );
  NAND2X1 U1029 ( .A(N942), .B(n2946), .Y(n3371) );
  NAND3X1 U1030 ( .A(n3459), .B(n3458), .C(n3457), .Y(n3577) );
  NAND2XL U1031 ( .A(next_A[20]), .B(n3034), .Y(n3458) );
  NAND2X1 U1032 ( .A(N815), .B(n2946), .Y(n3459) );
  NAND3X1 U1033 ( .A(n3289), .B(n3288), .C(n3287), .Y(n2876) );
  AOI21X1 U1034 ( .A0(SHA256_result[243]), .A1(n2984), .B0(n3114), .Y(n3289)
         );
  NAND2XL U1035 ( .A(next_A[19]), .B(n3036), .Y(n3288) );
  NAND3X1 U1036 ( .A(n3235), .B(n3234), .C(n3233), .Y(n2879) );
  NAND2XL U1037 ( .A(next_A[16]), .B(n3036), .Y(n3234) );
  NAND2X1 U1038 ( .A(N811), .B(n2946), .Y(n3233) );
  NAND3X1 U1039 ( .A(n3292), .B(n3291), .C(n3290), .Y(n2881) );
  AOI21X1 U1040 ( .A0(SHA256_result[238]), .A1(n2984), .B0(n3114), .Y(n3292)
         );
  NAND2XL U1041 ( .A(next_A[14]), .B(n3037), .Y(n3291) );
  NAND2X1 U1042 ( .A(N809), .B(n2944), .Y(n3290) );
  NAND3X1 U1043 ( .A(n3355), .B(n3354), .C(n3353), .Y(n3564) );
  NAND2X1 U1044 ( .A(n2872), .B(n3159), .Y(n3353) );
  NAND2XL U1045 ( .A(next_E[15]), .B(n3036), .Y(n3354) );
  NAND2X1 U1046 ( .A(N938), .B(n2945), .Y(n3355) );
  NAND3X1 U1047 ( .A(n3364), .B(n3363), .C(n3362), .Y(n3563) );
  NAND2X1 U1048 ( .A(n2875), .B(n3159), .Y(n3362) );
  NAND2X1 U1049 ( .A(N939), .B(n2945), .Y(n3364) );
  NAND3X1 U1050 ( .A(n3370), .B(n3369), .C(n3368), .Y(n2720) );
  AOI21X1 U1051 ( .A0(n2878), .A1(n2983), .B0(n3113), .Y(n3370) );
  NAND2XL U1052 ( .A(next_E[14]), .B(n3036), .Y(n3369) );
  NAND2X1 U1053 ( .A(N937), .B(n2947), .Y(n3368) );
  NAND3X1 U1054 ( .A(n3392), .B(n3391), .C(n3390), .Y(n2717) );
  AOI21X1 U1055 ( .A0(n2899), .A1(n2983), .B0(n3114), .Y(n3392) );
  NAND2XL U1056 ( .A(next_E[17]), .B(n3035), .Y(n3391) );
  NAND2X1 U1057 ( .A(N940), .B(n2947), .Y(n3390) );
  NAND3X1 U1058 ( .A(n3462), .B(n3461), .C(n3460), .Y(n3579) );
  NAND2XL U1059 ( .A(next_A[17]), .B(n3035), .Y(n3461) );
  NAND2X1 U1060 ( .A(N812), .B(n2947), .Y(n3462) );
  INVX1 U1061 ( .A(n2825), .Y(n3000) );
  INVX1 U1062 ( .A(n2825), .Y(n3001) );
  INVXL U1063 ( .A(n660), .Y(n3128) );
  INVX1 U1064 ( .A(n494), .Y(n3154) );
  INVX1 U1065 ( .A(n494), .Y(n3153) );
  INVX1 U1066 ( .A(n494), .Y(n3155) );
  INVX1 U1067 ( .A(n494), .Y(n3152) );
  NOR3X1 U1068 ( .A(n3778), .B(n2932), .C(n2817), .Y(n1301) );
  OAI221XL U1069 ( .A0(n1381), .A1(n3089), .B0(n2931), .B1(n1382), .C0(n1383), 
        .Y(N2966) );
  NOR4BXL U1070 ( .AN(n3732), .B(n1281), .C(n1387), .D(n1334), .Y(n1381) );
  OAI221XL U1071 ( .A0(n2932), .A1(n1388), .B0(n1389), .B1(n3742), .C0(n1376), 
        .Y(n1387) );
  AOI22X1 U1072 ( .A0(N999), .A1(n2935), .B0(n3034), .B1(SHA256_result[76]), 
        .Y(n923) );
  OAI211X1 U1073 ( .A0(n2980), .A1(n3771), .B0(n3112), .C0(n931), .Y(n2485) );
  AOI22X1 U1074 ( .A0(N1013), .A1(n2936), .B0(n3034), .B1(SHA256_result[90]), 
        .Y(n931) );
  AOI22X1 U1075 ( .A0(N998), .A1(n2935), .B0(n3034), .B1(SHA256_result[75]), 
        .Y(n922) );
  OAI211X1 U1076 ( .A0(n2976), .A1(n3792), .B0(n3109), .C0(n742), .Y(n2807) );
  AOI22X1 U1077 ( .A0(N851), .A1(n2939), .B0(n2888), .B1(n3032), .Y(n742) );
  OAI211X1 U1078 ( .A0(n2975), .A1(n3528), .B0(n3109), .C0(n743), .Y(n2806) );
  AOI22X1 U1079 ( .A0(N852), .A1(n2939), .B0(n2857), .B1(n3032), .Y(n743) );
  OAI211X1 U1080 ( .A0(n2981), .A1(n3793), .B0(n3112), .C0(n928), .Y(n2488) );
  AOI22X1 U1081 ( .A0(N1010), .A1(n2936), .B0(n3034), .B1(SHA256_result[87]), 
        .Y(n928) );
  OAI211X1 U1082 ( .A0(n2978), .A1(n3827), .B0(n3108), .C0(n734), .Y(n2820) );
  OAI211X1 U1083 ( .A0(n2981), .A1(n3825), .B0(n3111), .C0(n731), .Y(n2824) );
  OAI211X1 U1084 ( .A0(n2980), .A1(n3856), .B0(n3112), .C0(n932), .Y(n2484) );
  AOI22X1 U1085 ( .A0(N1014), .A1(n2936), .B0(n3034), .B1(SHA256_result[91]), 
        .Y(n932) );
  OAI211X1 U1086 ( .A0(n2980), .A1(n3855), .B0(n3112), .C0(n933), .Y(n2483) );
  AOI22X1 U1087 ( .A0(N1015), .A1(n2936), .B0(n3033), .B1(SHA256_result[92]), 
        .Y(n933) );
  OAI211X1 U1088 ( .A0(n2979), .A1(n3811), .B0(n3112), .C0(n925), .Y(n2496) );
  AOI22X1 U1089 ( .A0(N1002), .A1(n2941), .B0(n3034), .B1(n3808), .Y(n925) );
  OAI211X1 U1090 ( .A0(n2980), .A1(n3783), .B0(n3112), .C0(n930), .Y(n2486) );
  AOI22X1 U1091 ( .A0(N1012), .A1(n2936), .B0(n3034), .B1(SHA256_result[89]), 
        .Y(n930) );
  OAI211X1 U1092 ( .A0(n2980), .A1(n3782), .B0(n3112), .C0(n929), .Y(n2487) );
  AOI22X1 U1093 ( .A0(N1011), .A1(n2936), .B0(n3034), .B1(SHA256_result[88]), 
        .Y(n929) );
  OAI211X1 U1094 ( .A0(n3073), .A1(n3358), .B0(n3357), .C0(n3356), .Y(n3565)
         );
  INVX1 U1095 ( .A(next_E[13]), .Y(n3358) );
  NAND2X1 U1096 ( .A(N936), .B(n2946), .Y(n3357) );
  AOI211X1 U1097 ( .A0(n1307), .A1(round[4]), .B0(n1332), .C0(n1333), .Y(n1331) );
  AOI21X1 U1098 ( .A0(n3738), .A1(n3752), .B0(n2931), .Y(n1333) );
  NAND2XL U1099 ( .A(n3170), .B(n3167), .Y(n3706) );
  OAI22X1 U1100 ( .A0(n2960), .A1(n3190), .B0(n3040), .B1(n1168), .Y(n3192) );
  XOR3X2 U1101 ( .A(n2923), .B(n2855), .C(SHA256_result[243]), .Y(f3_A_32[17])
         );
  XOR3X2 U1102 ( .A(n2920), .B(SHA256_result[244]), .C(n2887), .Y(f3_A_32[18])
         );
  OAI211X1 U1103 ( .A0(n2979), .A1(n3818), .B0(n3111), .C0(n822), .Y(n2689) );
  XOR3X2 U1104 ( .A(n2924), .B(n2904), .C(n2849), .Y(f3_A_32[16]) );
  XOR3X2 U1105 ( .A(n2883), .B(n2871), .C(n2859), .Y(f4_E_32[19]) );
  NAND4X1 U1106 ( .A(n1450), .B(n1451), .C(n1452), .D(n1453), .Y(N2959) );
  NAND4X1 U1107 ( .A(n1501), .B(n1502), .C(n1503), .D(n1504), .Y(N2953) );
  NAND4X1 U1108 ( .A(n1459), .B(n1460), .C(n1461), .D(n1462), .Y(N2958) );
  OAI21XL U1109 ( .A0(n3707), .A1(n2712), .B0(n1334), .Y(n1460) );
  AOI31XL U1110 ( .A0(n1391), .A1(n2931), .A2(n2755), .B0(n1274), .Y(n1459) );
  XOR3X2 U1111 ( .A(n2877), .B(n2682), .C(n2873), .Y(f4_E_32[20]) );
  INVX1 U1112 ( .A(n1440), .Y(n3715) );
  AOI31X1 U1113 ( .A0(n2712), .A1(n2931), .A2(n2932), .B0(n1249), .Y(n1440) );
  INVX1 U1114 ( .A(N923), .Y(n3524) );
  OAI21XL U1115 ( .A0(n3060), .A1(n3816), .B0(n450), .Y(n1554) );
  INVX1 U1116 ( .A(n2909), .Y(n3816) );
  AOI22X1 U1117 ( .A0(N978), .A1(n2942), .B0(n3157), .B1(SHA256_result[87]), 
        .Y(n450) );
  NAND3X1 U1118 ( .A(n3329), .B(n3328), .C(n3327), .Y(n1569) );
  NAND2BX1 U1119 ( .AN(n2960), .B(N955), .Y(n3329) );
  NAND3X1 U1120 ( .A(n3465), .B(n3464), .C(n3463), .Y(n3581) );
  NAND2BX1 U1121 ( .AN(n2961), .B(N806), .Y(n3465) );
  NAND2BX1 U1122 ( .AN(n2963), .B(N972), .Y(n3501) );
  NAND2X1 U1123 ( .A(n3807), .B(n3157), .Y(n3500) );
  NAND3X1 U1124 ( .A(n3259), .B(n3258), .C(n3257), .Y(n1566) );
  NAND3X1 U1125 ( .A(n3332), .B(n3331), .C(n3330), .Y(n1564) );
  NAND2BX1 U1126 ( .AN(n2961), .B(N963), .Y(n3332) );
  NAND3X1 U1127 ( .A(n3436), .B(n3435), .C(n3434), .Y(n1561) );
  NAND2BX1 U1128 ( .AN(n2962), .B(N967), .Y(n3436) );
  NAND3X1 U1129 ( .A(n3498), .B(n3497), .C(n3496), .Y(n1560) );
  NAND2BX1 U1130 ( .AN(n2948), .B(N970), .Y(n3498) );
  NAND3X1 U1131 ( .A(n3512), .B(n3511), .C(n3510), .Y(n1568) );
  NAND2BX1 U1132 ( .AN(n2964), .B(N956), .Y(n3512) );
  OAI22X1 U1133 ( .A0(n2949), .A1(n3194), .B0(n3044), .B1(n3193), .Y(n3196) );
  OAI22X1 U1134 ( .A0(n2951), .A1(n3198), .B0(n3044), .B1(n3197), .Y(n3200) );
  INVXL U1135 ( .A(next_E[5]), .Y(n3197) );
  NAND2X1 U1136 ( .A(n2843), .B(n2986), .Y(n3245) );
  OAI22X1 U1137 ( .A0(n2960), .A1(n3244), .B0(n3045), .B1(n3243), .Y(n3246) );
  NAND3BX1 U1138 ( .AN(n3339), .B(n3112), .C(n3338), .Y(n2722) );
  NAND2X1 U1139 ( .A(n2859), .B(n2988), .Y(n3338) );
  OAI22X1 U1140 ( .A0(n2951), .A1(n3337), .B0(n3047), .B1(n3336), .Y(n3339) );
  INVXL U1141 ( .A(next_E[12]), .Y(n3336) );
  OAI22X1 U1142 ( .A0(n2951), .A1(n3347), .B0(n3048), .B1(n3346), .Y(n3349) );
  INVXL U1143 ( .A(next_E[9]), .Y(n3346) );
  OAI22X1 U1144 ( .A0(n2950), .A1(n3248), .B0(n3045), .B1(n3247), .Y(n3250) );
  OAI22X1 U1145 ( .A0(n2951), .A1(n3273), .B0(n3046), .B1(n3272), .Y(n3275) );
  OAI22X1 U1146 ( .A0(n2949), .A1(n3384), .B0(n3041), .B1(n3383), .Y(n3386) );
  INVXL U1147 ( .A(next_A[2]), .Y(n3383) );
  OAI22X1 U1148 ( .A0(n2950), .A1(n3410), .B0(n3041), .B1(n3409), .Y(n3412) );
  INVXL U1149 ( .A(next_A[1]), .Y(n3409) );
  NAND3BX1 U1150 ( .AN(n3440), .B(n3108), .C(n3439), .Y(n2885) );
  OAI22X1 U1151 ( .A0(n2950), .A1(n3438), .B0(n3048), .B1(n3437), .Y(n3440) );
  INVXL U1152 ( .A(n2404), .Y(n3437) );
  OAI22X1 U1153 ( .A0(n2949), .A1(n3442), .B0(n3049), .B1(n3441), .Y(n3444) );
  INVXL U1154 ( .A(n2381), .Y(n3441) );
  OAI22X1 U1155 ( .A0(n2949), .A1(n3473), .B0(n3042), .B1(n3472), .Y(n3475) );
  INVXL U1156 ( .A(next_A[6]), .Y(n3472) );
  OAI22X1 U1157 ( .A0(n2948), .A1(n3477), .B0(n3049), .B1(n3476), .Y(n3479) );
  INVXL U1158 ( .A(next_A[5]), .Y(n3476) );
  OAI22X1 U1159 ( .A0(n2948), .A1(n3517), .B0(n3043), .B1(n3516), .Y(n3519) );
  INVXL U1160 ( .A(next_A[0]), .Y(n3516) );
  NAND2X1 U1161 ( .A(n2833), .B(n2987), .Y(n3188) );
  OAI22X1 U1162 ( .A0(n2948), .A1(n3187), .B0(n3039), .B1(n3186), .Y(n3189) );
  INVXL U1163 ( .A(next_E[6]), .Y(n3186) );
  NAND3X1 U1164 ( .A(n3185), .B(n3184), .C(n3183), .Y(n3569) );
  NAND2BXL U1165 ( .AN(n3059), .B(next_E[7]), .Y(n3184) );
  NAND3X1 U1166 ( .A(n1493), .B(n1494), .C(n1495), .Y(N2954) );
  NAND3X1 U1167 ( .A(n3335), .B(n3334), .C(n3333), .Y(n3566) );
  NAND2BXL U1168 ( .AN(n3053), .B(next_E[11]), .Y(n3334) );
  NAND2BX1 U1169 ( .AN(n2960), .B(N934), .Y(n3335) );
  NAND3X1 U1170 ( .A(n3342), .B(n3341), .C(n3340), .Y(n3567) );
  NAND2BXL U1171 ( .AN(n3061), .B(next_E[10]), .Y(n3341) );
  NAND2BX1 U1172 ( .AN(n2961), .B(N933), .Y(n3342) );
  NAND2X1 U1173 ( .A(n2867), .B(n3159), .Y(n3340) );
  NAND3X1 U1174 ( .A(n3345), .B(n3344), .C(n3343), .Y(n3568) );
  NAND2BX1 U1175 ( .AN(n2962), .B(N931), .Y(n3345) );
  NAND2BXL U1176 ( .AN(n3060), .B(next_E[8]), .Y(n3344) );
  NAND3X1 U1177 ( .A(n3408), .B(n3407), .C(n3406), .Y(n3585) );
  NAND2BX1 U1178 ( .AN(n2962), .B(N798), .Y(n3408) );
  NAND2BXL U1179 ( .AN(n3055), .B(next_A[3]), .Y(n3407) );
  NAND3X1 U1180 ( .A(n3468), .B(n3467), .C(n3466), .Y(n3582) );
  NAND2BX1 U1181 ( .AN(n2964), .B(N803), .Y(n3468) );
  NAND2BXL U1182 ( .AN(n3043), .B(next_A[8]), .Y(n3467) );
  NAND3X1 U1183 ( .A(n3471), .B(n3470), .C(n3469), .Y(n3583) );
  NAND2BX1 U1184 ( .AN(n2963), .B(N802), .Y(n3471) );
  NAND2BXL U1185 ( .AN(n3051), .B(next_A[7]), .Y(n3470) );
  NAND3X1 U1186 ( .A(n3482), .B(n3481), .C(n3480), .Y(n3584) );
  NAND2BX1 U1187 ( .AN(n2949), .B(N799), .Y(n3482) );
  NAND2BXL U1188 ( .AN(n3042), .B(next_A[4]), .Y(n3481) );
  INVX1 U1189 ( .A(N935), .Y(n3337) );
  OAI2BB2X1 U1190 ( .B0(n1410), .B1(n3165), .A0N(n2931), .A1N(n1411), .Y(n1409) );
  INVX1 U1191 ( .A(n1320), .Y(n3092) );
  INVX1 U1192 ( .A(n447), .Y(n3163) );
  OAI22X1 U1193 ( .A0(n2817), .A1(n3751), .B0(n1322), .B1(n3089), .Y(n1282) );
  AOI22X1 U1194 ( .A0(n1323), .A1(n1248), .B0(n1324), .B1(n2932), .Y(n1322) );
  AOI22X1 U1195 ( .A0(n2713), .A1(n1259), .B0(n3711), .B1(n3165), .Y(n1338) );
  AOI31X1 U1196 ( .A0(n3763), .A1(n1284), .A2(n1343), .B0(n3089), .Y(n1341) );
  AOI22X1 U1197 ( .A0(n1380), .A1(n3765), .B0(n1324), .B1(n2932), .Y(n1508) );
  AOI31X1 U1198 ( .A0(n1518), .A1(n1519), .A2(n1520), .B0(n3089), .Y(n1517) );
  AOI22X1 U1199 ( .A0(n1420), .A1(n1484), .B0(n3756), .B1(round[4]), .Y(n1518)
         );
  AOI21XL U1200 ( .A0(n1281), .A1(n1248), .B0(n1332), .Y(n1519) );
  NOR4BX1 U1201 ( .AN(n3746), .B(n3743), .C(n1334), .D(n1309), .Y(n1520) );
  XOR3X2 U1202 ( .A(n2933), .B(n2907), .C(n2891), .Y(f3_A_32[19]) );
  XOR3X2 U1203 ( .A(SHA256_result[234]), .B(n2906), .C(n2901), .Y(f3_A_32[20])
         );
  XOR3X2 U1204 ( .A(SHA256_result[235]), .B(n2903), .C(n2892), .Y(f3_A_32[21])
         );
  AOI22X1 U1205 ( .A0(n3106), .A1(SHA256_result[88]), .B0(n3104), .B1(n2930), 
        .Y(n1122) );
  NOR2BX1 U1206 ( .AN(n1080), .B(N3079), .Y(n1094) );
  XOR3X2 U1207 ( .A(n2875), .B(n2860), .C(n2844), .Y(f4_E_32[23]) );
  XOR3X2 U1208 ( .A(SHA256_result[114]), .B(n2682), .C(n2837), .Y(f4_E_32[25])
         );
  NAND4X1 U1209 ( .A(n1344), .B(n1345), .C(n1346), .D(n1347), .Y(N2969) );
  OAI21XL U1210 ( .A0(n1303), .A1(n1355), .B0(n2713), .Y(n1345) );
  XOR3X2 U1211 ( .A(n2872), .B(n2874), .C(n2851), .Y(f4_E_32[22]) );
  XOR3X2 U1212 ( .A(n2899), .B(n2871), .C(n2843), .Y(f4_E_32[24]) );
  AOI21X1 U1213 ( .A0(n1428), .A1(n1429), .B0(n3089), .Y(n1427) );
  AOI211X1 U1214 ( .A0(n1258), .A1(n3165), .B0(n1390), .C0(n1430), .Y(n1429)
         );
  AOI211X1 U1215 ( .A0(n3757), .A1(n3164), .B0(n1431), .C0(n3731), .Y(n1428)
         );
  AOI21X1 U1216 ( .A0(n3767), .A1(n3761), .B0(n2388), .Y(n1430) );
  INVX1 U1217 ( .A(n2396), .Y(n3106) );
  INVX1 U1218 ( .A(n2393), .Y(n3098) );
  INVX1 U1219 ( .A(n2392), .Y(n3104) );
  NAND3X1 U1220 ( .A(n1514), .B(n1515), .C(n1516), .Y(N2951) );
  OAI21XL U1221 ( .A0(n1390), .A1(n1374), .B0(n1250), .Y(n1515) );
  INVX1 U1222 ( .A(N800), .Y(n3477) );
  INVX1 U1223 ( .A(N929), .Y(n3187) );
  INVX1 U1224 ( .A(N801), .Y(n3473) );
  INVX1 U1225 ( .A(N932), .Y(n3347) );
  INVX1 U1226 ( .A(n1320), .Y(n3091) );
  OAI211X1 U1227 ( .A0(n3723), .A1(n3724), .B0(n1078), .C0(n1079), .Y(N3081)
         );
  AOI31X1 U1228 ( .A0(n3725), .A1(n3723), .A2(n3724), .B0(n1080), .Y(n1079) );
  XOR3X2 U1229 ( .A(n2905), .B(SHA256_result[236]), .C(n2888), .Y(f3_A_32[22])
         );
  XOR3X2 U1230 ( .A(n2929), .B(n2857), .C(SHA256_result[237]), .Y(f3_A_32[23])
         );
  XOR3X2 U1231 ( .A(n2928), .B(n2916), .C(SHA256_result[238]), .Y(f3_A_32[24])
         );
  INVX1 U1232 ( .A(N927), .Y(n3194) );
  INVX1 U1233 ( .A(N928), .Y(n3198) );
  INVX1 U1234 ( .A(N925), .Y(n3248) );
  XOR3X2 U1235 ( .A(n2920), .B(n2919), .C(n2849), .Y(f3_A_32[27]) );
  XOR3X2 U1236 ( .A(n2924), .B(SHA256_result[251]), .C(SHA256_result[239]), 
        .Y(f3_A_32[25]) );
  XOR3X2 U1237 ( .A(n2923), .B(n2862), .C(SHA256_result[240]), .Y(f3_A_32[26])
         );
  XOR3X2 U1238 ( .A(n2851), .B(n2896), .C(n2833), .Y(f4_E_32[27]) );
  XOR3X2 U1239 ( .A(SHA256_result[104]), .B(n2910), .C(n2843), .Y(f4_E_32[29])
         );
  XOR3X2 U1240 ( .A(n2844), .B(n2915), .C(n2830), .Y(f4_E_32[28]) );
  NOR2X1 U1241 ( .A(n2388), .B(n2932), .Y(n1353) );
  NOR3X1 U1242 ( .A(n3776), .B(round[0]), .C(n2388), .Y(n1442) );
  AOI32X1 U1243 ( .A0(n2721), .A1(n2389), .A2(n1296), .B0(round[1]), .B1(n1277), .Y(n1330) );
  NOR2X1 U1244 ( .A(n3777), .B(n3165), .Y(n1354) );
  NOR2X1 U1245 ( .A(n3776), .B(n2932), .Y(n1337) );
  NOR2X1 U1246 ( .A(n2398), .B(round[1]), .Y(n1491) );
  OAI221XL U1247 ( .A0(n3752), .A1(n3775), .B0(n3763), .B1(n2932), .C0(n1465), 
        .Y(n1543) );
  AOI211XL U1248 ( .A0(n2766), .A1(n1362), .B0(n1363), .C0(n3744), .Y(n1360)
         );
  OAI21XL U1249 ( .A0(n1364), .A1(n3753), .B0(n3735), .Y(n1362) );
  AOI21X1 U1250 ( .A0(n3759), .A1(n3727), .B0(n2932), .Y(n1363) );
  NAND3X1 U1251 ( .A(n2931), .B(n2391), .C(n1389), .Y(n1457) );
  OAI211X1 U1252 ( .A0(n1446), .A1(n3765), .B0(n1447), .C0(n1448), .Y(n1445)
         );
  AOI21X1 U1253 ( .A0(n1449), .A1(n3165), .B0(n1391), .Y(n1447) );
  AOI222X1 U1254 ( .A0(n1295), .A1(n3745), .B0(n1294), .B1(n1248), .C0(n3743), 
        .C1(round[0]), .Y(n1448) );
  NAND4X1 U1255 ( .A(n3728), .B(n3727), .C(n1489), .D(n1490), .Y(n1488) );
  AOI22X1 U1256 ( .A0(n1491), .A1(n1261), .B0(n1308), .B1(n1492), .Y(n1489) );
  AOI221X1 U1257 ( .A0(n1391), .A1(round[0]), .B0(n3743), .B1(n3165), .C0(
        n3731), .Y(n1490) );
  XOR3X2 U1258 ( .A(n2869), .B(n2909), .C(n2837), .Y(f4_E_32[30]) );
  XOR3X2 U1259 ( .A(SHA256_result[234]), .B(n2887), .C(SHA256_result[243]), 
        .Y(f3_A_32[29]) );
  XOR3X2 U1260 ( .A(n2907), .B(n2904), .C(n2855), .Y(f3_A_32[28]) );
  XOR3X2 U1261 ( .A(n2933), .B(SHA256_result[235]), .C(SHA256_result[244]), 
        .Y(f3_A_32[30]) );
  INVX1 U1262 ( .A(N795), .Y(n3517) );
  INVX1 U1263 ( .A(n2931), .Y(n3777) );
  NOR2X1 U1264 ( .A(n2391), .B(round[4]), .Y(n1308) );
  NOR2X1 U1265 ( .A(round[4]), .B(n2932), .Y(n1296) );
  NOR2X1 U1266 ( .A(n2389), .B(round[0]), .Y(n1248) );
  NOR2X1 U1267 ( .A(n3750), .B(n2931), .Y(n1525) );
  OAI221XL U1268 ( .A0(n2931), .A1(n3732), .B0(n996), .B1(n3735), .C0(n3763), 
        .Y(n1279) );
  NOR2X1 U1269 ( .A(n3745), .B(n2931), .Y(n1335) );
  NAND2X1 U1270 ( .A(n1525), .B(round[1]), .Y(n1290) );
  NOR2X1 U1271 ( .A(n3753), .B(n2931), .Y(n1420) );
  NOR2X1 U1272 ( .A(n2391), .B(n2931), .Y(n1340) );
  OAI22X1 U1273 ( .A0(round[1]), .A1(n3778), .B0(n3760), .B1(n3775), .Y(n1492)
         );
  NOR2X1 U1274 ( .A(n3745), .B(n3165), .Y(n1265) );
  OAI211X1 U1275 ( .A0(n2932), .A1(n2390), .B0(n3740), .C0(n3776), .Y(n1526)
         );
  NOR2X1 U1276 ( .A(round[0]), .B(round[1]), .Y(n1364) );
  OAI211X1 U1277 ( .A0(n3750), .A1(n3766), .B0(n1473), .C0(n3767), .Y(n1472)
         );
  OAI21XL U1278 ( .A0(n1474), .A1(n3757), .B0(round[4]), .Y(n1473) );
  AOI31X1 U1279 ( .A0(n2931), .A1(n2391), .A2(n1310), .B0(n1311), .Y(n1304) );
  NAND2X1 U1280 ( .A(n1525), .B(round[0]), .Y(n1284) );
  NOR2X1 U1281 ( .A(n3737), .B(n2931), .Y(n1395) );
  OAI211X1 U1282 ( .A0(round[4]), .A1(n3164), .B0(n3751), .C0(n3747), .Y(n1417) );
  NAND2X1 U1283 ( .A(n1365), .B(n2931), .Y(n1298) );
  NOR2X1 U1284 ( .A(n3753), .B(n3165), .Y(n1260) );
  NAND4X1 U1285 ( .A(n3734), .B(n1278), .C(n3761), .D(n1533), .Y(n1532) );
  AOI22X1 U1286 ( .A0(n1340), .A1(n1484), .B0(n1390), .B1(n2932), .Y(n1533) );
  NAND2X1 U1287 ( .A(n1400), .B(round[1]), .Y(n1244) );
  AOI22X1 U1290 ( .A0(n1311), .A1(n2931), .B0(n1353), .B1(n3762), .Y(n1513) );
  OAI21XL U1291 ( .A0(n2932), .A1(n3762), .B0(n1290), .Y(n1449) );
  OAI2BB2X1 U1292 ( .B0(n3755), .B1(n2388), .A0N(n3165), .A1N(n1258), .Y(n1257) );
  OR2X2 U1293 ( .A(n3750), .B(n3165), .Y(n2819) );
  INVX1 U1294 ( .A(n2819), .Y(n1281) );
  NAND4BXL U1295 ( .AN(n1549), .B(n3759), .C(n1284), .D(n1550), .Y(n1548) );
  AOI211X1 U1296 ( .A0(n3749), .A1(n3165), .B0(n1431), .C0(n3754), .Y(n1550)
         );
  OAI21XL U1297 ( .A0(n3738), .A1(n2390), .B0(n1319), .Y(n1549) );
  INVX1 U1298 ( .A(n1290), .Y(n3749) );
  NAND4X1 U1299 ( .A(n1457), .B(n2796), .C(n3761), .D(n1458), .Y(n1456) );
  AOI22X1 U1300 ( .A0(n1307), .A1(n2932), .B0(n1310), .B1(n1296), .Y(n1458) );
  NAND3X1 U1301 ( .A(n3746), .B(n1298), .C(n1539), .Y(n1538) );
  OAI21XL U1302 ( .A0(n3743), .A1(n1365), .B0(n3165), .Y(n1539) );
  AOI21X1 U1303 ( .A0(n3757), .A1(n3165), .B0(n1307), .Y(n1343) );
  INVX1 U1304 ( .A(N992), .Y(n3240) );
  INVX1 U1305 ( .A(N995), .Y(n3305) );
  AOI221X1 U1306 ( .A0(n1484), .A1(n1321), .B0(round[4]), .B1(n1467), .C0(
        n3756), .Y(n1483) );
  INVX1 U1307 ( .A(n3165), .Y(n3164) );
  NOR2X1 U1308 ( .A(n2388), .B(n3165), .Y(n1475) );
  NOR2X1 U1309 ( .A(n2932), .B(n2931), .Y(n1380) );
  NOR2X1 U1310 ( .A(n2391), .B(n3165), .Y(n1317) );
  NOR2X1 U1311 ( .A(n3723), .B(n3725), .Y(n1080) );
  INVX1 U1312 ( .A(N829), .Y(n3173) );
  INVX1 U1313 ( .A(N990), .Y(n3278) );
  INVX1 U1314 ( .A(SHA256_result[238]), .Y(n3486) );
  INVX1 U1315 ( .A(SHA256_result[243]), .Y(n3504) );
  INVX1 U1316 ( .A(n2899), .Y(n3499) );
  MX2X1 U1317 ( .A(SHA256_result[63]), .B(SHA256_result[95]), .S0(n2682), .Y(
        f1_EFG_32[31]) );
  BUFX20 U1318 ( .A(SHA256_result[225]), .Y(n2906) );
  BUFX20 U1319 ( .A(SHA256_result[98]), .Y(n2844) );
  BUFX20 U1320 ( .A(SHA256_result[224]), .Y(n2933) );
  BUFX20 U1321 ( .A(SHA256_result[97]), .Y(n2851) );
  BUFX20 U1322 ( .A(SHA256_result[228]), .Y(n2929) );
  BUFX20 U1323 ( .A(SHA256_result[123]), .Y(n2864) );
  BUFX20 U1324 ( .A(SHA256_result[226]), .Y(n2892) );
  BUFX20 U1325 ( .A(SHA256_result[105]), .Y(n2869) );
  BUFX20 U1326 ( .A(SHA256_result[246]), .Y(n2901) );
  BUFX20 U1327 ( .A(SHA256_result[124]), .Y(n2874) );
  BUFX20 U1328 ( .A(SHA256_result[247]), .Y(n2903) );
  BUFX20 U1329 ( .A(SHA256_result[122]), .Y(n2877) );
  BUFX20 U1330 ( .A(SHA256_result[111]), .Y(n2872) );
  BUFX20 U1331 ( .A(SHA256_result[248]), .Y(n2888) );
  BUFX20 U1332 ( .A(SHA256_result[107]), .Y(n2858) );
  BUFX20 U1333 ( .A(SHA256_result[108]), .Y(n2859) );
  BUFX20 U1334 ( .A(SHA256_result[100]), .Y(n2837) );
  BUFX20 U1335 ( .A(SHA256_result[110]), .Y(n2878) );
  BUFX20 U1336 ( .A(SHA256_result[101]), .Y(n2840) );
  BUFX20 U1337 ( .A(SHA256_result[109]), .Y(n2873) );
  BUFX8 U1338 ( .A(SHA256_result[255]), .Y(n2887) );
  OAI2BB1X1 U1339 ( .A0N(SHA256_result[196]), .A1N(n2929), .B0(n3228), .Y(
        f2_ABC_32[4]) );
  OAI21XL U1340 ( .A0(SHA256_result[196]), .A1(n2929), .B0(SHA256_result[164]), 
        .Y(n3228) );
  OAI21XL U1341 ( .A0(SHA256_result[163]), .A1(SHA256_result[195]), .B0(n2905), 
        .Y(n3229) );
  OAI2BB1X1 U1342 ( .A0N(n2892), .A1N(SHA256_result[162]), .B0(n3230), .Y(
        f2_ABC_32[2]) );
  OAI21XL U1343 ( .A0(SHA256_result[162]), .A1(n2892), .B0(SHA256_result[194]), 
        .Y(n3230) );
  MX2X1 U1344 ( .A(SHA256_result[42]), .B(SHA256_result[74]), .S0(n2867), .Y(
        n330) );
  BUFX20 U1345 ( .A(SHA256_result[242]), .Y(n2904) );
  BUFX20 U1346 ( .A(SHA256_result[241]), .Y(n2919) );
  MX2X1 U1347 ( .A(SHA256_result[40]), .B(SHA256_result[72]), .S0(
        SHA256_result[104]), .Y(f1_EFG_32[8]) );
  BUFX20 U1348 ( .A(SHA256_result[233]), .Y(n2907) );
  BUFX20 U1349 ( .A(SHA256_result[116]), .Y(n2896) );
  BUFX20 U1350 ( .A(SHA256_result[230]), .Y(n2924) );
  BUFX20 U1351 ( .A(SHA256_result[229]), .Y(n2928) );
  BUFX8 U1352 ( .A(SHA256_result[252]), .Y(n2862) );
  BUFX8 U1353 ( .A(SHA256_result[126]), .Y(n2871) );
  BUFX20 U1354 ( .A(SHA256_result[117]), .Y(n2915) );
  BUFX20 U1355 ( .A(SHA256_result[250]), .Y(n2916) );
  BUFX20 U1356 ( .A(SHA256_result[249]), .Y(n2857) );
  BUFX8 U1357 ( .A(SHA256_result[125]), .Y(n2860) );
  BUFX20 U1358 ( .A(SHA256_result[115]), .Y(n2884) );
  BUFX20 U1359 ( .A(SHA256_result[231]), .Y(n2923) );
  BUFX8 U1360 ( .A(SHA256_result[253]), .Y(n2849) );
  BUFX20 U1361 ( .A(SHA256_result[232]), .Y(n2920) );
  MXI2XL U1362 ( .A(n3809), .B(n1152), .S0(n2875), .Y(f1_EFG_32[16]) );
  MXI2XL U1363 ( .A(n3831), .B(n1157), .S0(n2858), .Y(f1_EFG_32[11]) );
  MXI2XL U1364 ( .A(n3821), .B(n1154), .S0(n2878), .Y(f1_EFG_32[14]) );
  MXI2XL U1365 ( .A(n3819), .B(n1156), .S0(n2859), .Y(f1_EFG_32[12]) );
  MXI2XL U1366 ( .A(n3810), .B(n1151), .S0(n2899), .Y(f1_EFG_32[17]) );
  MXI2XL U1367 ( .A(n3811), .B(n1153), .S0(n2872), .Y(f1_EFG_32[15]) );
  OAI2BB1X1 U1368 ( .A0N(SHA256_result[200]), .A1N(n2920), .B0(n3224), .Y(
        f2_ABC_32[8]) );
  OAI21XL U1369 ( .A0(SHA256_result[200]), .A1(n2920), .B0(SHA256_result[168]), 
        .Y(n3224) );
  OAI21X4 U1370 ( .A0(output_enable), .A1(inner_busy), .B0(n1434), .Y(n656) );
  OAI211X1 U1371 ( .A0(n2977), .A1(n3853), .B0(n3110), .C0(n765), .Y(n2770) );
  AOI22X1 U1372 ( .A0(N887), .A1(n2941), .B0(SHA256_result[220]), .B1(n3030), 
        .Y(n765) );
  INVX1 U1373 ( .A(SHA256_result[159]), .Y(n3841) );
  OAI211X1 U1374 ( .A0(n2978), .A1(n3847), .B0(n3108), .C0(n949), .Y(n2449) );
  INVX1 U1375 ( .A(SHA256_result[30]), .Y(n3847) );
  AOI22X1 U1376 ( .A0(N1049), .A1(n2937), .B0(SHA256_result[62]), .B1(n3032), 
        .Y(n949) );
  OAI211X1 U1377 ( .A0(n2979), .A1(n3844), .B0(n3111), .C0(n784), .Y(n2737) );
  INVX1 U1378 ( .A(SHA256_result[157]), .Y(n3844) );
  AOI22X1 U1379 ( .A0(N920), .A1(n2972), .B0(SHA256_result[189]), .B1(n3029), 
        .Y(n784) );
  OAI211X1 U1380 ( .A0(n2981), .A1(n3854), .B0(n3112), .C0(n947), .Y(n2452) );
  AOI22X1 U1381 ( .A0(N1046), .A1(n2937), .B0(SHA256_result[59]), .B1(n3027), 
        .Y(n947) );
  OAI211X1 U1382 ( .A0(n2981), .A1(n3849), .B0(n3112), .C0(n948), .Y(n2451) );
  INVX1 U1383 ( .A(SHA256_result[28]), .Y(n3849) );
  AOI22X1 U1384 ( .A0(N1047), .A1(n2937), .B0(SHA256_result[60]), .B1(n3027), 
        .Y(n948) );
  OAI211X1 U1385 ( .A0(n2975), .A1(n3552), .B0(n3109), .C0(n745), .Y(n2803) );
  INVX1 U1386 ( .A(SHA256_result[220]), .Y(n3552) );
  AOI22XL U1387 ( .A0(N855), .A1(n2939), .B0(n2862), .B1(n3032), .Y(n745) );
  OAI211X1 U1388 ( .A0(n2980), .A1(n3846), .B0(n3111), .C0(n783), .Y(n2740) );
  AOI22X1 U1389 ( .A0(N917), .A1(n2973), .B0(SHA256_result[186]), .B1(n3029), 
        .Y(n783) );
  OAI211X1 U1390 ( .A0(n2977), .A1(n3550), .B0(n3110), .C0(n766), .Y(n2769) );
  INVX1 U1391 ( .A(SHA256_result[189]), .Y(n3550) );
  OAI211X1 U1392 ( .A0(n2975), .A1(n3549), .B0(n3109), .C0(n746), .Y(n2802) );
  INVX1 U1393 ( .A(SHA256_result[221]), .Y(n3549) );
  AOI22XL U1394 ( .A0(N856), .A1(n2939), .B0(n2849), .B1(n3032), .Y(n746) );
  OAI2BB1X1 U1395 ( .A0N(SHA256_result[175]), .A1N(SHA256_result[207]), .B0(
        n3217), .Y(f2_ABC_32[15]) );
  OAI21XL U1396 ( .A0(SHA256_result[207]), .A1(SHA256_result[175]), .B0(
        SHA256_result[239]), .Y(n3217) );
  OAI2BB1X1 U1397 ( .A0N(n2907), .A1N(SHA256_result[169]), .B0(n3223), .Y(
        f2_ABC_32[9]) );
  OAI21XL U1398 ( .A0(n2907), .A1(SHA256_result[169]), .B0(SHA256_result[201]), 
        .Y(n3223) );
  OAI2BB1X2 U1399 ( .A0N(SHA256_result[172]), .A1N(SHA256_result[204]), .B0(
        n3220), .Y(f2_ABC_32[12]) );
  OAI21XL U1400 ( .A0(SHA256_result[205]), .A1(SHA256_result[173]), .B0(
        SHA256_result[237]), .Y(n3219) );
  OAI2BB1X1 U1401 ( .A0N(SHA256_result[174]), .A1N(SHA256_result[206]), .B0(
        n3218), .Y(f2_ABC_32[14]) );
  OAI21XL U1402 ( .A0(SHA256_result[174]), .A1(SHA256_result[206]), .B0(
        SHA256_result[238]), .Y(n3218) );
  OAI211X1 U1403 ( .A0(n1140), .A1(n2982), .B0(n3112), .C0(n829), .Y(n2674) );
  AOI22XL U1404 ( .A0(N983), .A1(n2935), .B0(n2874), .B1(n3028), .Y(n829) );
  OAI211X1 U1405 ( .A0(n1141), .A1(n2982), .B0(n3111), .C0(n828), .Y(n2675) );
  AOI22XL U1406 ( .A0(N982), .A1(n2935), .B0(n2864), .B1(n3028), .Y(n828) );
  OAI211X1 U1407 ( .A0(n1143), .A1(n2982), .B0(n3111), .C0(n827), .Y(n2677) );
  AOI22XL U1408 ( .A0(N980), .A1(n2935), .B0(n2883), .B1(n3028), .Y(n827) );
  MX2X1 U1409 ( .A(SHA256_result[45]), .B(SHA256_result[77]), .S0(n2873), .Y(
        f1_EFG_32[13]) );
  AND2X4 U1410 ( .A(n2745), .B(round[6]), .Y(n2823) );
  OAI21XL U1411 ( .A0(n3053), .A1(n3853), .B0(n481), .Y(n1584) );
  AOI22X1 U1412 ( .A0(N919), .A1(n2942), .B0(SHA256_result[156]), .B1(n3156), 
        .Y(n481) );
  OAI21XL U1413 ( .A0(n3052), .A1(n3852), .B0(n482), .Y(n1585) );
  AOI22X1 U1414 ( .A0(N918), .A1(n2942), .B0(SHA256_result[155]), .B1(n3158), 
        .Y(n482) );
  OAI21XL U1415 ( .A0(n3051), .A1(n3548), .B0(n480), .Y(n1583) );
  INVX1 U1416 ( .A(SHA256_result[190]), .Y(n3548) );
  AOI22X1 U1417 ( .A0(N921), .A1(n2943), .B0(SHA256_result[158]), .B1(n3157), 
        .Y(n480) );
  OAI21XL U1418 ( .A0(n3061), .A1(n3845), .B0(n513), .Y(n1611) );
  INVX1 U1419 ( .A(SHA256_result[222]), .Y(n3845) );
  AOI22X1 U1420 ( .A0(N889), .A1(n2944), .B0(SHA256_result[190]), .B1(n3156), 
        .Y(n513) );
  INVX1 U1421 ( .A(SHA256_result[63]), .Y(n3842) );
  OAI21XL U1422 ( .A0(n3058), .A1(n3851), .B0(n498), .Y(n1596) );
  OAI21XL U1423 ( .A0(n3063), .A1(n3848), .B0(n526), .Y(n1624) );
  AOI22X1 U1424 ( .A0(N1016), .A1(n2938), .B0(SHA256_result[61]), .B1(n3156), 
        .Y(n526) );
  AOI22X1 U1425 ( .A0(N857), .A1(n2943), .B0(SHA256_result[222]), .B1(n3157), 
        .Y(n466) );
  XOR3X2 U1426 ( .A(n2867), .B(n2930), .C(n2840), .Y(f4_E_32[31]) );
  NAND3X1 U1427 ( .A(n3271), .B(n3270), .C(n3269), .Y(n1551) );
  NAND2XL U1428 ( .A(n2871), .B(n3037), .Y(n3270) );
  NAND2X1 U1429 ( .A(N985), .B(n2947), .Y(n3271) );
  NAND3X1 U1430 ( .A(n3268), .B(n3267), .C(n3266), .Y(n1552) );
  NAND2XL U1431 ( .A(n2860), .B(n3037), .Y(n3267) );
  NAND2XL U1432 ( .A(n3013), .B(SHA256_result[71]), .Y(n3503) );
  OAI2BB1X1 U1433 ( .A0N(H6[0]), .A1N(n3138), .B0(n899), .Y(n2542) );
  OAI2BB1X1 U1434 ( .A0N(H4[0]), .A1N(n3140), .B0(n844), .Y(n2638) );
  BUFX8 U1435 ( .A(SHA256_result[254]), .Y(n2855) );
  OAI2BB1X1 U1436 ( .A0N(SHA256_result[94]), .A1N(n3038), .B0(n525), .Y(n1623)
         );
  AOI22X1 U1437 ( .A0(N1017), .A1(n2938), .B0(SHA256_result[62]), .B1(n3157), 
        .Y(n525) );
  AOI21XL U1438 ( .A0(SHA256_result[192]), .A1(n3008), .B0(n3125), .Y(n710) );
  OAI2BB1X1 U1439 ( .A0N(H1[18]), .A1N(n3140), .B0(n720), .Y(n2845) );
  AOI21XL U1440 ( .A0(SHA256_result[210]), .A1(n3008), .B0(n3125), .Y(n720) );
  OAI2BB1X1 U1441 ( .A0N(H1[15]), .A1N(n3141), .B0(n717), .Y(n2848) );
  AOI21XL U1442 ( .A0(SHA256_result[207]), .A1(n3010), .B0(n3125), .Y(n717) );
  OAI2BB1X1 U1443 ( .A0N(H1[17]), .A1N(n3141), .B0(n719), .Y(n2846) );
  AOI21XL U1444 ( .A0(SHA256_result[209]), .A1(n3010), .B0(n3125), .Y(n719) );
  OAI2BB1X1 U1445 ( .A0N(H1[9]), .A1N(n3141), .B0(n713), .Y(n2854) );
  AOI21XL U1446 ( .A0(SHA256_result[201]), .A1(n3010), .B0(n3125), .Y(n713) );
  OAI2BB1X1 U1447 ( .A0N(H2[4]), .A1N(n3139), .B0(n880), .Y(n2571) );
  AOI21XL U1448 ( .A0(SHA256_result[164]), .A1(n3005), .B0(n3120), .Y(n880) );
  OAI2BB1X1 U1449 ( .A0N(H2[19]), .A1N(n3139), .B0(n891), .Y(n2556) );
  OAI2BB1X1 U1450 ( .A0N(H2[15]), .A1N(n3139), .B0(n888), .Y(n2560) );
  AOI21XL U1451 ( .A0(SHA256_result[175]), .A1(n3005), .B0(n3119), .Y(n888) );
  OAI2BB1X1 U1452 ( .A0N(H1[16]), .A1N(n3141), .B0(n718), .Y(n2847) );
  AOI21XL U1453 ( .A0(SHA256_result[208]), .A1(n3009), .B0(n3125), .Y(n718) );
  OAI2BB1X1 U1454 ( .A0N(H6[11]), .A1N(n3133), .B0(n905), .Y(n2531) );
  AOI21XL U1455 ( .A0(SHA256_result[43]), .A1(n3004), .B0(n3118), .Y(n905) );
  OAI2BB1X1 U1456 ( .A0N(H6[3]), .A1N(n3140), .B0(n901), .Y(n2539) );
  AOI21XL U1457 ( .A0(SHA256_result[35]), .A1(n3004), .B0(n3118), .Y(n901) );
  OAI2BB1X1 U1458 ( .A0N(H2[22]), .A1N(n3139), .B0(n893), .Y(n2553) );
  AOI21XL U1459 ( .A0(SHA256_result[182]), .A1(n3005), .B0(n3119), .Y(n893) );
  OAI2BB1X1 U1460 ( .A0N(H3[13]), .A1N(n3140), .B0(n867), .Y(n2593) );
  OAI2BB1X1 U1461 ( .A0N(H6[23]), .A1N(n3138), .B0(n911), .Y(n2519) );
  OAI2BB1X1 U1462 ( .A0N(H1[21]), .A1N(n3140), .B0(n721), .Y(n2842) );
  OAI2BB1X1 U1463 ( .A0N(H2[5]), .A1N(n3139), .B0(n881), .Y(n2570) );
  AOI21XL U1464 ( .A0(SHA256_result[165]), .A1(n3005), .B0(n3120), .Y(n881) );
  OAI2BB1X1 U1465 ( .A0N(H2[12]), .A1N(n3139), .B0(n885), .Y(n2563) );
  AOI21XL U1466 ( .A0(SHA256_result[172]), .A1(n3005), .B0(n3119), .Y(n885) );
  OAI2BB1X1 U1467 ( .A0N(H2[14]), .A1N(n3139), .B0(n887), .Y(n2561) );
  AOI21XL U1468 ( .A0(SHA256_result[174]), .A1(n3005), .B0(n3119), .Y(n887) );
  OAI2BB1X1 U1469 ( .A0N(H2[26]), .A1N(n3139), .B0(n894), .Y(n2549) );
  AOI21XL U1470 ( .A0(SHA256_result[186]), .A1(n3004), .B0(n3119), .Y(n894) );
  OAI2BB1X1 U1471 ( .A0N(H1[13]), .A1N(n3141), .B0(n716), .Y(n2850) );
  AOI21XL U1472 ( .A0(SHA256_result[205]), .A1(n3008), .B0(n3125), .Y(n716) );
  OAI2BB1X1 U1473 ( .A0N(H1[29]), .A1N(n3135), .B0(n727), .Y(n2834) );
  AOI21XL U1474 ( .A0(SHA256_result[221]), .A1(n3009), .B0(n3124), .Y(n727) );
  OAI2BB1X1 U1475 ( .A0N(H2[13]), .A1N(n3139), .B0(n886), .Y(n2562) );
  AOI21XL U1476 ( .A0(SHA256_result[173]), .A1(n3005), .B0(n3119), .Y(n886) );
  OAI2BB1X1 U1477 ( .A0N(H2[17]), .A1N(n3139), .B0(n889), .Y(n2558) );
  AOI21XL U1478 ( .A0(SHA256_result[177]), .A1(n3005), .B0(n3119), .Y(n889) );
  OAI2BB1X1 U1479 ( .A0N(H2[18]), .A1N(n3139), .B0(n890), .Y(n2557) );
  AOI21XL U1480 ( .A0(SHA256_result[178]), .A1(n3005), .B0(n3119), .Y(n890) );
  OAI2BB1X1 U1481 ( .A0N(H2[29]), .A1N(n3135), .B0(n897), .Y(n2546) );
  AOI21XL U1482 ( .A0(SHA256_result[189]), .A1(n3004), .B0(n3118), .Y(n897) );
  AOI21XL U1483 ( .A0(n2685), .A1(n3004), .B0(n3118), .Y(n900) );
  OAI2BB1X1 U1484 ( .A0N(H1[22]), .A1N(n3131), .B0(n722), .Y(n2841) );
  AOI21XL U1485 ( .A0(SHA256_result[214]), .A1(n3008), .B0(n3124), .Y(n722) );
  OAI2BB1X1 U1486 ( .A0N(H1[28]), .A1N(n3139), .B0(n726), .Y(n2835) );
  AOI21XL U1487 ( .A0(SHA256_result[220]), .A1(n3008), .B0(n3124), .Y(n726) );
  OAI2BB1X1 U1488 ( .A0N(H1[27]), .A1N(n3134), .B0(n725), .Y(n2836) );
  AOI21XL U1489 ( .A0(SHA256_result[219]), .A1(n3009), .B0(n3124), .Y(n725) );
  AOI21XL U1490 ( .A0(SHA256_result[161]), .A1(n3005), .B0(n3120), .Y(n879) );
  OAI2BB1X1 U1491 ( .A0N(H3[22]), .A1N(n3139), .B0(n874), .Y(n2584) );
  AOI21XL U1492 ( .A0(SHA256_result[150]), .A1(n3006), .B0(n3120), .Y(n874) );
  OAI2BB1X1 U1493 ( .A0N(H3[16]), .A1N(n3140), .B0(n870), .Y(n2590) );
  AOI21XL U1494 ( .A0(SHA256_result[144]), .A1(n3006), .B0(n3121), .Y(n870) );
  OAI2BB1X1 U1495 ( .A0N(H3[4]), .A1N(n3140), .B0(n862), .Y(n2602) );
  AOI21XL U1496 ( .A0(SHA256_result[132]), .A1(n3007), .B0(n3121), .Y(n862) );
  OAI2BB1X1 U1497 ( .A0N(H3[19]), .A1N(n3139), .B0(n873), .Y(n2587) );
  AOI21XL U1498 ( .A0(SHA256_result[147]), .A1(n3006), .B0(n3120), .Y(n873) );
  OAI2BB1X1 U1499 ( .A0N(H5[13]), .A1N(n3139), .B0(n835), .Y(n2657) );
  AOI21XL U1500 ( .A0(SHA256_result[77]), .A1(n3009), .B0(n3124), .Y(n835) );
  OAI2BB1X1 U1501 ( .A0N(H7[11]), .A1N(n3136), .B0(n957), .Y(n2436) );
  AOI21XL U1502 ( .A0(SHA256_result[11]), .A1(n3002), .B0(n3116), .Y(n957) );
  OAI2BB1X1 U1503 ( .A0N(H7[8]), .A1N(n3133), .B0(n955), .Y(n2439) );
  AOI21XL U1504 ( .A0(SHA256_result[8]), .A1(n3003), .B0(n3117), .Y(n955) );
  OAI2BB1X1 U1505 ( .A0N(H3[17]), .A1N(n3139), .B0(n871), .Y(n2589) );
  AOI21XL U1506 ( .A0(SHA256_result[145]), .A1(n3006), .B0(n3121), .Y(n871) );
  OAI2BB1X1 U1507 ( .A0N(H3[18]), .A1N(n3139), .B0(n872), .Y(n2588) );
  AOI21XL U1508 ( .A0(SHA256_result[146]), .A1(n3006), .B0(n3120), .Y(n872) );
  AOI21XL U1509 ( .A0(SHA256_result[194]), .A1(n3010), .B0(n3125), .Y(n711) );
  OAI2BB1X1 U1510 ( .A0N(H6[8]), .A1N(n3131), .B0(n904), .Y(n2534) );
  AOI21XL U1511 ( .A0(SHA256_result[40]), .A1(n3004), .B0(n3118), .Y(n904) );
  OAI2BB1X1 U1512 ( .A0N(H2[8]), .A1N(n3139), .B0(n883), .Y(n2567) );
  AOI21XL U1513 ( .A0(SHA256_result[168]), .A1(n3005), .B0(n3120), .Y(n883) );
  OAI2BB1X1 U1514 ( .A0N(H3[26]), .A1N(n3139), .B0(n876), .Y(n2580) );
  AOI21XL U1515 ( .A0(SHA256_result[154]), .A1(n3006), .B0(n3120), .Y(n876) );
  OAI2BB1X1 U1516 ( .A0N(H7[30]), .A1N(n3139), .B0(n967), .Y(n2417) );
  AOI21XL U1517 ( .A0(SHA256_result[30]), .A1(n3002), .B0(n3116), .Y(n967) );
  OAI2BB1X1 U1518 ( .A0N(H7[21]), .A1N(n3139), .B0(n960), .Y(n2426) );
  AOI21XL U1519 ( .A0(SHA256_result[21]), .A1(n3002), .B0(n3116), .Y(n960) );
  OAI2BB1X1 U1521 ( .A0N(H7[22]), .A1N(n3139), .B0(n961), .Y(n2425) );
  AOI21XL U1522 ( .A0(SHA256_result[22]), .A1(n3002), .B0(n3116), .Y(n961) );
  OAI2BB1X1 U1523 ( .A0N(H7[23]), .A1N(n3139), .B0(n962), .Y(n2424) );
  AOI21XL U1524 ( .A0(SHA256_result[23]), .A1(n3002), .B0(n3116), .Y(n962) );
  OAI2BB1X1 U1525 ( .A0N(H7[25]), .A1N(n3140), .B0(n964), .Y(n2422) );
  AOI21XL U1526 ( .A0(SHA256_result[25]), .A1(n3002), .B0(n3116), .Y(n964) );
  OAI2BB1X1 U1527 ( .A0N(H7[24]), .A1N(n3139), .B0(n963), .Y(n2423) );
  AOI21XL U1528 ( .A0(SHA256_result[24]), .A1(n3002), .B0(n3116), .Y(n963) );
  OAI2BB1X1 U1529 ( .A0N(H7[28]), .A1N(n3140), .B0(n966), .Y(n2419) );
  AOI21XL U1530 ( .A0(SHA256_result[28]), .A1(n3002), .B0(n3116), .Y(n966) );
  OAI2BB1X1 U1531 ( .A0N(H7[27]), .A1N(n3141), .B0(n965), .Y(n2420) );
  AOI21XL U1532 ( .A0(SHA256_result[27]), .A1(n3002), .B0(n3116), .Y(n965) );
  OAI2BB1X1 U1533 ( .A0N(H1[24]), .A1N(n3136), .B0(n723), .Y(n2839) );
  AOI21XL U1534 ( .A0(SHA256_result[216]), .A1(n3009), .B0(n3124), .Y(n723) );
  OAI2BB1X1 U1535 ( .A0N(H1[25]), .A1N(n3139), .B0(n724), .Y(n2838) );
  AOI21XL U1536 ( .A0(SHA256_result[217]), .A1(n3008), .B0(n3124), .Y(n724) );
  OAI2BB1X1 U1537 ( .A0N(H2[6]), .A1N(n3139), .B0(n882), .Y(n2569) );
  AOI21XL U1538 ( .A0(n3011), .A1(SHA256_result[166]), .B0(n3120), .Y(n882) );
  OAI2BB1X1 U1539 ( .A0N(H3[29]), .A1N(n3139), .B0(n877), .Y(n2577) );
  AOI21XL U1540 ( .A0(SHA256_result[157]), .A1(n3006), .B0(n3120), .Y(n877) );
  OAI2BB1X1 U1541 ( .A0N(H7[14]), .A1N(n3139), .B0(n958), .Y(n2433) );
  AOI21XL U1542 ( .A0(SHA256_result[14]), .A1(n3002), .B0(n3116), .Y(n958) );
  OAI2BB1X1 U1543 ( .A0N(H3[5]), .A1N(n3140), .B0(n863), .Y(n2601) );
  AOI21XL U1544 ( .A0(SHA256_result[133]), .A1(n3007), .B0(n3121), .Y(n863) );
  OAI2BB1X1 U1545 ( .A0N(H3[14]), .A1N(n3140), .B0(n868), .Y(n2592) );
  AOI21XL U1546 ( .A0(SHA256_result[142]), .A1(n3006), .B0(n3121), .Y(n868) );
  OAI2BB1X1 U1547 ( .A0N(H7[10]), .A1N(n3140), .B0(n956), .Y(n2437) );
  AOI21XL U1548 ( .A0(SHA256_result[10]), .A1(n3002), .B0(n3116), .Y(n956) );
  OAI2BB1X1 U1549 ( .A0N(H7[4]), .A1N(n3134), .B0(n954), .Y(n2443) );
  AOI21XL U1550 ( .A0(SHA256_result[4]), .A1(n3003), .B0(n3117), .Y(n954) );
  AOI21XL U1551 ( .A0(SHA256_result[129]), .A1(n3007), .B0(n3121), .Y(n860) );
  OAI2BB1X1 U1552 ( .A0N(H1[31]), .A1N(n3139), .B0(n728), .Y(n2832) );
  AOI21XL U1553 ( .A0(SHA256_result[223]), .A1(n3008), .B0(n3124), .Y(n728) );
  OAI2BB1X1 U1554 ( .A0N(H6[25]), .A1N(n3141), .B0(n913), .Y(n2517) );
  AOI21XL U1555 ( .A0(SHA256_result[57]), .A1(n3003), .B0(n3117), .Y(n913) );
  OAI2BB1X1 U1556 ( .A0N(H6[24]), .A1N(n3135), .B0(n912), .Y(n2518) );
  AOI21XL U1557 ( .A0(SHA256_result[56]), .A1(n3003), .B0(n3117), .Y(n912) );
  OAI2BB1X1 U1558 ( .A0N(H6[28]), .A1N(n3131), .B0(n916), .Y(n2514) );
  AOI21XL U1559 ( .A0(SHA256_result[60]), .A1(n3003), .B0(n3117), .Y(n916) );
  OAI2BB1X1 U1560 ( .A0N(H6[27]), .A1N(n3134), .B0(n915), .Y(n2515) );
  AOI21XL U1561 ( .A0(SHA256_result[59]), .A1(n3003), .B0(n3117), .Y(n915) );
  OAI2BB1X1 U1562 ( .A0N(H6[15]), .A1N(n3140), .B0(n908), .Y(n2527) );
  AOI21XL U1563 ( .A0(SHA256_result[47]), .A1(n3004), .B0(n3118), .Y(n908) );
  OAI2BB1X1 U1564 ( .A0N(H6[14]), .A1N(n3139), .B0(n907), .Y(n2528) );
  AOI21XL U1565 ( .A0(SHA256_result[46]), .A1(n3004), .B0(n3118), .Y(n907) );
  OAI2BB1X1 U1566 ( .A0N(H5[2]), .A1N(n3138), .B0(n831), .Y(n2668) );
  AOI21XL U1567 ( .A0(SHA256_result[66]), .A1(n3009), .B0(n3124), .Y(n831) );
  OAI2BB1X1 U1568 ( .A0N(H6[5]), .A1N(n3138), .B0(n902), .Y(n2537) );
  AOI21XL U1569 ( .A0(SHA256_result[37]), .A1(n3004), .B0(n3118), .Y(n902) );
  OAI2BB1X1 U1570 ( .A0N(H6[7]), .A1N(n3132), .B0(n903), .Y(n2535) );
  AOI21XL U1571 ( .A0(SHA256_result[39]), .A1(n3004), .B0(n3118), .Y(n903) );
  OAI2BB1X1 U1572 ( .A0N(H1[7]), .A1N(n3141), .B0(n712), .Y(n2856) );
  AOI21XL U1573 ( .A0(SHA256_result[199]), .A1(n3009), .B0(n3125), .Y(n712) );
  OAI2BB1X1 U1574 ( .A0N(H1[10]), .A1N(n3141), .B0(n714), .Y(n2853) );
  AOI21XL U1575 ( .A0(SHA256_result[202]), .A1(n3009), .B0(n3125), .Y(n714) );
  OAI2BB1X1 U1576 ( .A0N(H1[11]), .A1N(n3141), .B0(n715), .Y(n2852) );
  AOI21XL U1577 ( .A0(SHA256_result[203]), .A1(n3010), .B0(n3125), .Y(n715) );
  OAI2BB1X1 U1578 ( .A0N(H3[3]), .A1N(n3140), .B0(n861), .Y(n2603) );
  AOI21XL U1579 ( .A0(SHA256_result[131]), .A1(n3007), .B0(n3121), .Y(n861) );
  OAI2BB1X1 U1580 ( .A0N(H2[9]), .A1N(n3139), .B0(n884), .Y(n2566) );
  AOI21XL U1581 ( .A0(n3012), .A1(SHA256_result[169]), .B0(n3119), .Y(n884) );
  OAI2BB1X1 U1582 ( .A0N(H2[21]), .A1N(n3139), .B0(n892), .Y(n2554) );
  AOI21XL U1583 ( .A0(n3011), .A1(SHA256_result[181]), .B0(n3119), .Y(n892) );
  OAI2BB1X1 U1584 ( .A0N(H7[15]), .A1N(n3139), .B0(n959), .Y(n2432) );
  AOI21XL U1585 ( .A0(SHA256_result[15]), .A1(n3002), .B0(n3116), .Y(n959) );
  AOI21XL U1586 ( .A0(SHA256_result[3]), .A1(n3003), .B0(n3117), .Y(n953) );
  OAI2BB1X1 U1587 ( .A0N(H3[8]), .A1N(n3140), .B0(n864), .Y(n2598) );
  AOI21XL U1588 ( .A0(SHA256_result[136]), .A1(n3007), .B0(n3121), .Y(n864) );
  OAI2BB1X1 U1589 ( .A0N(H3[12]), .A1N(n3140), .B0(n866), .Y(n2594) );
  AOI21XL U1590 ( .A0(SHA256_result[140]), .A1(n3007), .B0(n3121), .Y(n866) );
  OAI2BB1X1 U1591 ( .A0N(H3[10]), .A1N(n3140), .B0(n865), .Y(n2596) );
  AOI21XL U1592 ( .A0(SHA256_result[138]), .A1(n3007), .B0(n3121), .Y(n865) );
  OAI2BB1X1 U1593 ( .A0N(H5[31]), .A1N(n3136), .B0(n843), .Y(n2639) );
  AOI21XL U1594 ( .A0(SHA256_result[95]), .A1(n3008), .B0(n3123), .Y(n843) );
  OAI2BB1X1 U1595 ( .A0N(H3[24]), .A1N(n3139), .B0(n875), .Y(n2582) );
  AOI21XL U1596 ( .A0(SHA256_result[152]), .A1(n3006), .B0(n3120), .Y(n875) );
  OAI2BB1X1 U1597 ( .A0N(H5[18]), .A1N(n3140), .B0(n838), .Y(n2652) );
  AOI21XL U1598 ( .A0(SHA256_result[82]), .A1(n3008), .B0(n3123), .Y(n838) );
  OAI2BB1X1 U1599 ( .A0N(H3[31]), .A1N(n3139), .B0(n878), .Y(n2575) );
  AOI21XL U1600 ( .A0(SHA256_result[159]), .A1(n3006), .B0(n3120), .Y(n878) );
  OAI2BB1X1 U1601 ( .A0N(H2[27]), .A1N(n3132), .B0(n895), .Y(n2548) );
  AOI21XL U1602 ( .A0(n3011), .A1(SHA256_result[187]), .B0(n3119), .Y(n895) );
  OAI2BB1X1 U1603 ( .A0N(H2[28]), .A1N(n3137), .B0(n896), .Y(n2547) );
  AOI21XL U1604 ( .A0(n3012), .A1(SHA256_result[188]), .B0(n3118), .Y(n896) );
  OAI2BB1X1 U1605 ( .A0N(H3[15]), .A1N(n3132), .B0(n869), .Y(n2591) );
  AOI21XL U1606 ( .A0(SHA256_result[143]), .A1(n3006), .B0(n3121), .Y(n869) );
  OAI2BB1X1 U1607 ( .A0N(H6[16]), .A1N(n3136), .B0(n909), .Y(n2526) );
  AOI21XL U1608 ( .A0(SHA256_result[48]), .A1(n3003), .B0(n3117), .Y(n909) );
  OAI2BB1X1 U1609 ( .A0N(H6[17]), .A1N(n3134), .B0(n910), .Y(n2525) );
  AOI21XL U1610 ( .A0(SHA256_result[49]), .A1(n3003), .B0(n3117), .Y(n910) );
  OAI2BB1X1 U1611 ( .A0N(H6[26]), .A1N(n3132), .B0(n914), .Y(n2516) );
  AOI21XL U1612 ( .A0(SHA256_result[58]), .A1(n3003), .B0(n3117), .Y(n914) );
  OAI2BB1X1 U1613 ( .A0N(H6[12]), .A1N(n3133), .B0(n906), .Y(n2530) );
  AOI21XL U1614 ( .A0(SHA256_result[44]), .A1(n3004), .B0(n3118), .Y(n906) );
  OAI2BB1X1 U1615 ( .A0N(H4[6]), .A1N(n3140), .B0(n850), .Y(n2632) );
  AOI21XL U1616 ( .A0(n3012), .A1(n2833), .B0(n3122), .Y(n850) );
  AOI21XL U1617 ( .A0(SHA256_result[0]), .A1(n3003), .B0(n3117), .Y(n952) );
  OAI2BB1X1 U1618 ( .A0N(H5[11]), .A1N(n3139), .B0(n834), .Y(n2659) );
  AOI21XL U1619 ( .A0(n3012), .A1(SHA256_result[75]), .B0(n3124), .Y(n834) );
  OAI2BB1X1 U1620 ( .A0N(H5[25]), .A1N(n3140), .B0(n840), .Y(n2645) );
  AOI21XL U1621 ( .A0(n3011), .A1(SHA256_result[89]), .B0(n3123), .Y(n840) );
  OAI2BB1X1 U1622 ( .A0N(H5[16]), .A1N(n3139), .B0(n837), .Y(n2654) );
  AOI21XL U1623 ( .A0(n3011), .A1(SHA256_result[80]), .B0(n3123), .Y(n837) );
  OAI2BB1X1 U1624 ( .A0N(H5[14]), .A1N(n3131), .B0(n836), .Y(n2656) );
  AOI21XL U1625 ( .A0(n3011), .A1(SHA256_result[78]), .B0(n3123), .Y(n836) );
  OAI2BB1X1 U1626 ( .A0N(H5[24]), .A1N(n3140), .B0(n839), .Y(n2646) );
  AOI21XL U1627 ( .A0(n3011), .A1(SHA256_result[88]), .B0(n3123), .Y(n839) );
  OAI2BB1X1 U1628 ( .A0N(H5[27]), .A1N(n3132), .B0(n841), .Y(n2643) );
  AOI21XL U1629 ( .A0(n3011), .A1(SHA256_result[91]), .B0(n3123), .Y(n841) );
  OAI2BB1X1 U1630 ( .A0N(H5[28]), .A1N(n3136), .B0(n842), .Y(n2642) );
  AOI21XL U1631 ( .A0(n3011), .A1(SHA256_result[92]), .B0(n3123), .Y(n842) );
  OAI2BB1X1 U1632 ( .A0N(H5[3]), .A1N(n3137), .B0(n832), .Y(n2667) );
  AOI21XL U1633 ( .A0(n3011), .A1(SHA256_result[67]), .B0(n3124), .Y(n832) );
  OAI2BB1X1 U1634 ( .A0N(H4[9]), .A1N(n3140), .B0(n851), .Y(n2629) );
  AOI21XL U1635 ( .A0(n3010), .A1(n2869), .B0(n3122), .Y(n851) );
  OAI2BB1X1 U1636 ( .A0N(H4[5]), .A1N(n3140), .B0(n849), .Y(n2633) );
  AOI21XL U1637 ( .A0(n3010), .A1(n2840), .B0(n3122), .Y(n849) );
  OAI2BB1X1 U1638 ( .A0N(H4[12]), .A1N(n3140), .B0(n852), .Y(n2626) );
  AOI21XL U1639 ( .A0(n3011), .A1(n2859), .B0(n3122), .Y(n852) );
  OAI2BB1X1 U1640 ( .A0N(H4[4]), .A1N(n3140), .B0(n848), .Y(n2634) );
  AOI21XL U1641 ( .A0(n3011), .A1(n2837), .B0(n3122), .Y(n848) );
  OAI2BB1X1 U1642 ( .A0N(H4[19]), .A1N(n3140), .B0(n856), .Y(n2619) );
  AOI21XL U1643 ( .A0(n3011), .A1(n2884), .B0(n3122), .Y(n856) );
  OAI2BB1X1 U1644 ( .A0N(H4[1]), .A1N(n3139), .B0(n845), .Y(n2637) );
  AOI21XL U1645 ( .A0(n3010), .A1(n2851), .B0(n3123), .Y(n845) );
  OAI2BB1X1 U1646 ( .A0N(H0[14]), .A1N(n3141), .B0(n668), .Y(n2913) );
  AOI21XL U1647 ( .A0(n3012), .A1(SHA256_result[238]), .B0(n3126), .Y(n668) );
  OAI2BB1X1 U1648 ( .A0N(H0[6]), .A1N(n3140), .B0(n664), .Y(n2921) );
  AOI21XL U1649 ( .A0(n3012), .A1(n2924), .B0(n3126), .Y(n664) );
  OAI2BB1X1 U1650 ( .A0N(H0[5]), .A1N(n3139), .B0(n663), .Y(n2922) );
  AOI21XL U1651 ( .A0(n3012), .A1(n2928), .B0(n3126), .Y(n663) );
  OAI2BB1X1 U1652 ( .A0N(H0[19]), .A1N(n3141), .B0(n671), .Y(n2908) );
  AOI21XL U1653 ( .A0(n3012), .A1(SHA256_result[243]), .B0(n3126), .Y(n671) );
  OAI2BB1X1 U1654 ( .A0N(H4[17]), .A1N(n3140), .B0(n854), .Y(n2621) );
  AOI21XL U1655 ( .A0(n3012), .A1(n2899), .B0(n3122), .Y(n854) );
  OAI2BB1X1 U1656 ( .A0N(H4[30]), .A1N(n3140), .B0(n859), .Y(n2608) );
  AOI21XL U1657 ( .A0(n3012), .A1(n2871), .B0(n3122), .Y(n859) );
  OAI2BB1X1 U1658 ( .A0N(H0[30]), .A1N(n3141), .B0(n675), .Y(n2897) );
  AOI21XL U1659 ( .A0(n3012), .A1(n2855), .B0(n3125), .Y(n675) );
  OAI2BB1X1 U1660 ( .A0N(H0[1]), .A1N(n3135), .B0(n661), .Y(n2926) );
  AOI21XL U1661 ( .A0(n3012), .A1(n2906), .B0(n3119), .Y(n661) );
  OAI2BB1X1 U1662 ( .A0N(H0[15]), .A1N(n3141), .B0(n669), .Y(n2912) );
  AOI21XL U1663 ( .A0(SHA256_result[239]), .A1(n3010), .B0(n3126), .Y(n669) );
  OAI2BB1X1 U1664 ( .A0N(H0[13]), .A1N(n3141), .B0(n667), .Y(n2914) );
  AOI21XL U1665 ( .A0(SHA256_result[237]), .A1(n3010), .B0(n3126), .Y(n667) );
  OAI2BB1X1 U1666 ( .A0N(H0[9]), .A1N(n3140), .B0(n665), .Y(n2918) );
  AOI21XL U1667 ( .A0(n2907), .A1(n3010), .B0(n3126), .Y(n665) );
  OAI2BB1X1 U1668 ( .A0N(H0[27]), .A1N(n3141), .B0(n673), .Y(n2900) );
  AOI21XL U1669 ( .A0(SHA256_result[251]), .A1(n3010), .B0(n3126), .Y(n673) );
  OAI2BB1X1 U1670 ( .A0N(H0[10]), .A1N(n3139), .B0(n666), .Y(n2917) );
  AOI21XL U1671 ( .A0(SHA256_result[234]), .A1(n3009), .B0(n3126), .Y(n666) );
  OAI2BB1X1 U1672 ( .A0N(H4[24]), .A1N(n3140), .B0(n857), .Y(n2614) );
  AOI21XL U1673 ( .A0(n2930), .A1(n3007), .B0(n3122), .Y(n857) );
  OAI2BB1X1 U1674 ( .A0N(H4[2]), .A1N(n3133), .B0(n846), .Y(n2636) );
  AOI21XL U1675 ( .A0(n2844), .A1(n3007), .B0(n3123), .Y(n846) );
  OAI2BB1X1 U1676 ( .A0N(H0[16]), .A1N(n3141), .B0(n670), .Y(n2911) );
  AOI21XL U1677 ( .A0(SHA256_result[240]), .A1(n3008), .B0(n3126), .Y(n670) );
  OAI2BB1X1 U1678 ( .A0N(H0[0]), .A1N(n3137), .B0(n659), .Y(n2927) );
  AOI21XL U1679 ( .A0(n2933), .A1(n3009), .B0(n3119), .Y(n659) );
  OAI2BB1X1 U1680 ( .A0N(H4[14]), .A1N(n3140), .B0(n853), .Y(n2624) );
  AOI21XL U1681 ( .A0(n2878), .A1(n3008), .B0(n3122), .Y(n853) );
  OAI2BB1X1 U1682 ( .A0N(H4[18]), .A1N(n3140), .B0(n855), .Y(n2620) );
  AOI21XL U1683 ( .A0(SHA256_result[114]), .A1(n3007), .B0(n3122), .Y(n855) );
  OAI2BB1X1 U1684 ( .A0N(H0[25]), .A1N(n3141), .B0(n672), .Y(n2902) );
  AOI21XL U1685 ( .A0(n2857), .A1(n3007), .B0(n3126), .Y(n672) );
  OAI2BB1X1 U1686 ( .A0N(H4[28]), .A1N(n3140), .B0(n858), .Y(n2610) );
  AOI21XL U1687 ( .A0(n2874), .A1(n3007), .B0(n3122), .Y(n858) );
  OAI2BB1X1 U1688 ( .A0N(H0[29]), .A1N(n3141), .B0(n674), .Y(n2898) );
  AOI21XL U1689 ( .A0(n2849), .A1(n3009), .B0(n3126), .Y(n674) );
  OAI2BB1X1 U1690 ( .A0N(H4[3]), .A1N(n3140), .B0(n847), .Y(n2635) );
  AOI21XL U1691 ( .A0(n2843), .A1(n3008), .B0(n3123), .Y(n847) );
  OAI2BB1X1 U1692 ( .A0N(H0[2]), .A1N(n3140), .B0(n662), .Y(n2925) );
  AOI21XL U1693 ( .A0(n2892), .A1(n3009), .B0(n3119), .Y(n662) );
  INVX1 U1694 ( .A(n598), .Y(n3642) );
  AOI22XL U1695 ( .A0(n3149), .A1(SHA256_result[163]), .B0(H2[3]), .B1(n3134), 
        .Y(n598) );
  INVX1 U1696 ( .A(n606), .Y(n3634) );
  INVX1 U1697 ( .A(n605), .Y(n3635) );
  AOI22XL U1698 ( .A0(n3149), .A1(SHA256_result[42]), .B0(H6[10]), .B1(n3134), 
        .Y(n605) );
  INVX1 U1699 ( .A(n604), .Y(n3636) );
  INVX1 U1700 ( .A(n551), .Y(n3689) );
  INVX1 U1701 ( .A(n595), .Y(n3645) );
  AOI22XL U1702 ( .A0(n3149), .A1(SHA256_result[170]), .B0(H2[10]), .B1(n3134), 
        .Y(n595) );
  INVX1 U1703 ( .A(n591), .Y(n3649) );
  INVX1 U1704 ( .A(n569), .Y(n3671) );
  INVX1 U1705 ( .A(n592), .Y(n3648) );
  AOI22XL U1706 ( .A0(n3149), .A1(SHA256_result[1]), .B0(H7[1]), .B1(n3135), 
        .Y(n592) );
  INVX1 U1707 ( .A(n590), .Y(n3650) );
  INVX1 U1708 ( .A(n634), .Y(n3606) );
  INVX1 U1709 ( .A(n603), .Y(n3637) );
  AOI22XL U1710 ( .A0(n3149), .A1(SHA256_result[36]), .B0(H6[4]), .B1(n3134), 
        .Y(n603) );
  INVX1 U1711 ( .A(n545), .Y(n3695) );
  INVX1 U1712 ( .A(n615), .Y(n3625) );
  INVX1 U1713 ( .A(n635), .Y(n3605) );
  INVX1 U1714 ( .A(n597), .Y(n3643) );
  INVX1 U1715 ( .A(n566), .Y(n3674) );
  INVX1 U1716 ( .A(n550), .Y(n3690) );
  INVX1 U1717 ( .A(n552), .Y(n3688) );
  INVX1 U1718 ( .A(n608), .Y(n3632) );
  AOI22XL U1719 ( .A0(n3150), .A1(SHA256_result[45]), .B0(H6[13]), .B1(n3133), 
        .Y(n608) );
  INVX1 U1720 ( .A(n611), .Y(n3629) );
  INVX1 U1721 ( .A(n609), .Y(n3631) );
  INVX1 U1722 ( .A(n610), .Y(n3630) );
  INVX1 U1723 ( .A(n549), .Y(n3691) );
  INVX1 U1724 ( .A(n624), .Y(n3616) );
  AOI22XL U1725 ( .A0(n3150), .A1(SHA256_result[13]), .B0(H7[13]), .B1(n3135), 
        .Y(n624) );
  INVX1 U1726 ( .A(n644), .Y(n3596) );
  AOI22XL U1727 ( .A0(n3151), .A1(SHA256_result[12]), .B0(H7[12]), .B1(n3131), 
        .Y(n644) );
  INVX1 U1728 ( .A(n623), .Y(n3617) );
  AOI22XL U1729 ( .A0(n3150), .A1(SHA256_result[5]), .B0(H7[5]), .B1(n3132), 
        .Y(n623) );
  INVX1 U1730 ( .A(n601), .Y(n3639) );
  AOI22XL U1731 ( .A0(n3149), .A1(SHA256_result[34]), .B0(H6[2]), .B1(n3134), 
        .Y(n601) );
  INVX1 U1732 ( .A(n602), .Y(n3638) );
  AOI22XL U1733 ( .A0(n3149), .A1(SHA256_result[38]), .B0(H6[6]), .B1(n3134), 
        .Y(n602) );
  INVX1 U1734 ( .A(n607), .Y(n3633) );
  AOI22XL U1735 ( .A0(n3150), .A1(SHA256_result[41]), .B0(H6[9]), .B1(n3133), 
        .Y(n607) );
  INVX1 U1736 ( .A(n620), .Y(n3620) );
  AOI22XL U1737 ( .A0(n3150), .A1(SHA256_result[2]), .B0(H7[2]), .B1(n3131), 
        .Y(n620) );
  INVX1 U1738 ( .A(n616), .Y(n3624) );
  AOI22XL U1739 ( .A0(n3150), .A1(SHA256_result[9]), .B0(H7[9]), .B1(n3133), 
        .Y(n616) );
  INVX1 U1740 ( .A(n643), .Y(n3597) );
  AOI22XL U1741 ( .A0(n3151), .A1(SHA256_result[6]), .B0(H7[6]), .B1(n3131), 
        .Y(n643) );
  INVX1 U1742 ( .A(n596), .Y(n3644) );
  AOI22XL U1743 ( .A0(n3149), .A1(SHA256_result[7]), .B0(H7[7]), .B1(n3134), 
        .Y(n596) );
  INVX1 U1744 ( .A(n553), .Y(n3687) );
  INVX1 U1745 ( .A(n649), .Y(n3591) );
  AOI22XL U1746 ( .A0(SHA256_result[193]), .A1(n3144), .B0(H1[1]), .B1(n3131), 
        .Y(n649) );
  INVX1 U1747 ( .A(n650), .Y(n3590) );
  AOI22XL U1748 ( .A0(SHA256_result[196]), .A1(n3144), .B0(H1[4]), .B1(n3131), 
        .Y(n650) );
  INVX1 U1749 ( .A(n637), .Y(n3603) );
  AOI22XL U1750 ( .A0(SHA256_result[200]), .A1(n3145), .B0(H1[8]), .B1(n3132), 
        .Y(n637) );
  INVX1 U1751 ( .A(n638), .Y(n3602) );
  INVX1 U1752 ( .A(n587), .Y(n3653) );
  AOI22XL U1753 ( .A0(SHA256_result[197]), .A1(n3147), .B0(H1[5]), .B1(n3135), 
        .Y(n587) );
  INVX1 U1754 ( .A(n493), .Y(n3705) );
  AOI22XL U1755 ( .A0(n3148), .A1(n2887), .B0(H0[31]), .B1(n3134), .Y(n493) );
  INVX1 U1756 ( .A(n542), .Y(n3698) );
  INVX1 U1757 ( .A(n617), .Y(n3623) );
  AOI22XL U1758 ( .A0(SHA256_result[160]), .A1(n3146), .B0(H2[0]), .B1(n3133), 
        .Y(n617) );
  INVX1 U1759 ( .A(n646), .Y(n3594) );
  INVX1 U1760 ( .A(n629), .Y(n3611) );
  AOI22XL U1761 ( .A0(SHA256_result[73]), .A1(n3145), .B0(H5[9]), .B1(n3135), 
        .Y(n629) );
  INVX1 U1762 ( .A(n584), .Y(n3656) );
  INVX1 U1763 ( .A(n593), .Y(n3647) );
  AOI22XL U1764 ( .A0(n3722), .A1(n3151), .B0(H5[1]), .B1(n3135), .Y(n593) );
  INVX1 U1765 ( .A(n641), .Y(n3599) );
  AOI22XL U1766 ( .A0(SHA256_result[130]), .A1(n3144), .B0(H3[2]), .B1(n3132), 
        .Y(n641) );
  INVX1 U1767 ( .A(n614), .Y(n3626) );
  AOI22XL U1768 ( .A0(SHA256_result[162]), .A1(n3146), .B0(H2[2]), .B1(n3133), 
        .Y(n614) );
  INVX1 U1769 ( .A(n586), .Y(n3654) );
  AOI22XL U1770 ( .A0(SHA256_result[195]), .A1(n3150), .B0(H1[3]), .B1(n3135), 
        .Y(n586) );
  INVX1 U1771 ( .A(n636), .Y(n3604) );
  AOI22XL U1772 ( .A0(SHA256_result[68]), .A1(n3144), .B0(H5[4]), .B1(n3132), 
        .Y(n636) );
  INVX1 U1773 ( .A(n642), .Y(n3598) );
  AOI22XL U1774 ( .A0(n3837), .A1(n3144), .B0(H5[0]), .B1(n3132), .Y(n642) );
  INVX1 U1775 ( .A(n648), .Y(n3592) );
  AOI22XL U1776 ( .A0(SHA256_result[198]), .A1(n3144), .B0(H1[6]), .B1(n3131), 
        .Y(n648) );
  INVX1 U1777 ( .A(n621), .Y(n3619) );
  INVX1 U1778 ( .A(n627), .Y(n3613) );
  AOI22XL U1779 ( .A0(SHA256_result[70]), .A1(n3145), .B0(H5[6]), .B1(n3131), 
        .Y(n627) );
  INVX1 U1780 ( .A(n640), .Y(n3600) );
  INVX1 U1781 ( .A(n645), .Y(n3595) );
  INVX1 U1782 ( .A(n599), .Y(n3641) );
  AOI22XL U1783 ( .A0(SHA256_result[167]), .A1(n3147), .B0(H2[7]), .B1(n3134), 
        .Y(n599) );
  INVX1 U1784 ( .A(n626), .Y(n3614) );
  INVX1 U1785 ( .A(n613), .Y(n3627) );
  INVX1 U1786 ( .A(n628), .Y(n3612) );
  AOI22XL U1787 ( .A0(SHA256_result[74]), .A1(n3145), .B0(H5[10]), .B1(n3135), 
        .Y(n628) );
  INVX1 U1788 ( .A(n583), .Y(n3657) );
  INVX1 U1789 ( .A(n600), .Y(n3640) );
  AOI22XL U1790 ( .A0(SHA256_result[171]), .A1(n3147), .B0(H2[11]), .B1(n3134), 
        .Y(n600) );
  INVX1 U1791 ( .A(n618), .Y(n3622) );
  INVX1 U1792 ( .A(n594), .Y(n3646) );
  INVX1 U1793 ( .A(n622), .Y(n3618) );
  INVX1 U1794 ( .A(n652), .Y(n3588) );
  AOI22XL U1795 ( .A0(n3150), .A1(SHA256_result[235]), .B0(H0[11]), .B1(n3131), 
        .Y(n652) );
  INVX1 U1796 ( .A(n619), .Y(n3621) );
  AOI22XL U1797 ( .A0(n2905), .A1(n3146), .B0(H0[3]), .B1(n3133), .Y(n619) );
  INVX1 U1798 ( .A(n630), .Y(n3610) );
  INVX1 U1799 ( .A(n631), .Y(n3609) );
  INVX1 U1800 ( .A(n632), .Y(n3608) );
  INVX1 U1801 ( .A(n647), .Y(n3593) );
  INVX1 U1802 ( .A(n612), .Y(n3628) );
  INVX1 U1803 ( .A(n585), .Y(n3655) );
  INVX1 U1804 ( .A(n589), .Y(n3651) );
  INVX1 U1805 ( .A(n588), .Y(n3652) );
  INVX1 U1806 ( .A(n633), .Y(n3607) );
  INVX1 U1807 ( .A(n653), .Y(n3587) );
  AOI22XL U1808 ( .A0(SHA256_result[236]), .A1(n3144), .B0(H0[12]), .B1(n3131), 
        .Y(n653) );
  INVX1 U1809 ( .A(n654), .Y(n3586) );
  AOI22XL U1810 ( .A0(n2920), .A1(n3144), .B0(H0[8]), .B1(n3131), .Y(n654) );
  INVX1 U1811 ( .A(n651), .Y(n3589) );
  AOI22XL U1812 ( .A0(n2929), .A1(n3144), .B0(H0[4]), .B1(n3131), .Y(n651) );
  INVX1 U1813 ( .A(n582), .Y(n3658) );
  AOI22XL U1814 ( .A0(n3149), .A1(n2891), .B0(H0[21]), .B1(n3136), .Y(n582) );
  INVX1 U1815 ( .A(n581), .Y(n3659) );
  INVX1 U1816 ( .A(n580), .Y(n3660) );
  AOI22XL U1817 ( .A0(n3148), .A1(n2919), .B0(H0[17]), .B1(n3136), .Y(n580) );
  INVX1 U1818 ( .A(n579), .Y(n3661) );
  AOI22XL U1819 ( .A0(SHA256_result[104]), .A1(n3151), .B0(H4[8]), .B1(n3136), 
        .Y(n579) );
  INVX1 U1820 ( .A(n578), .Y(n3662) );
  AOI22XL U1821 ( .A0(n3148), .A1(n2830), .B0(H4[7]), .B1(n3136), .Y(n578) );
  INVX1 U1822 ( .A(n577), .Y(n3663) );
  AOI22XL U1823 ( .A0(n3148), .A1(n2858), .B0(H4[11]), .B1(n3136), .Y(n577) );
  INVX1 U1824 ( .A(n576), .Y(n3664) );
  AOI22XL U1825 ( .A0(n2872), .A1(n3150), .B0(H4[15]), .B1(n3136), .Y(n576) );
  INVX1 U1826 ( .A(n575), .Y(n3665) );
  AOI22XL U1827 ( .A0(n3148), .A1(n2873), .B0(H4[13]), .B1(n3136), .Y(n575) );
  INVX1 U1828 ( .A(n574), .Y(n3666) );
  AOI22XL U1829 ( .A0(n2867), .A1(n3150), .B0(H4[10]), .B1(n3136), .Y(n574) );
  INVX1 U1830 ( .A(n573), .Y(n3667) );
  AOI22XL U1831 ( .A0(n3148), .A1(n2875), .B0(H4[16]), .B1(n3136), .Y(n573) );
  INVX1 U1832 ( .A(n572), .Y(n3668) );
  INVX1 U1833 ( .A(n571), .Y(n3669) );
  INVX1 U1834 ( .A(n570), .Y(n3670) );
  INVX1 U1835 ( .A(n568), .Y(n3672) );
  INVX1 U1836 ( .A(n567), .Y(n3673) );
  INVX1 U1837 ( .A(n565), .Y(n3675) );
  INVX1 U1838 ( .A(n564), .Y(n3676) );
  AOI22XL U1839 ( .A0(SHA256_result[244]), .A1(n3150), .B0(H0[20]), .B1(n3137), 
        .Y(n564) );
  INVX1 U1840 ( .A(n563), .Y(n3677) );
  AOI22XL U1841 ( .A0(n3150), .A1(n2904), .B0(H0[18]), .B1(n3137), .Y(n563) );
  INVX1 U1842 ( .A(n562), .Y(n3678) );
  AOI22XL U1843 ( .A0(n2903), .A1(n3147), .B0(H0[23]), .B1(n3137), .Y(n562) );
  INVX1 U1844 ( .A(n561), .Y(n3679) );
  AOI22XL U1845 ( .A0(n3150), .A1(n2864), .B0(H4[27]), .B1(n3137), .Y(n561) );
  INVX1 U1846 ( .A(n560), .Y(n3680) );
  AOI22XL U1847 ( .A0(n2915), .A1(n3150), .B0(H4[21]), .B1(n3137), .Y(n560) );
  INVX1 U1848 ( .A(n559), .Y(n3681) );
  AOI22XL U1849 ( .A0(n2896), .A1(n3150), .B0(H4[20]), .B1(n3136), .Y(n559) );
  AOI22XL U1850 ( .A0(n3148), .A1(n2883), .B0(H4[25]), .B1(n3133), .Y(n558) );
  INVX1 U1851 ( .A(n557), .Y(n3683) );
  AOI22XL U1852 ( .A0(n2860), .A1(n3147), .B0(H4[29]), .B1(n3140), .Y(n557) );
  INVX1 U1853 ( .A(n556), .Y(n3684) );
  AOI22XL U1854 ( .A0(n2909), .A1(n3147), .B0(H4[23]), .B1(n3139), .Y(n556) );
  INVX1 U1855 ( .A(n555), .Y(n3685) );
  AOI22XL U1856 ( .A0(n2877), .A1(n3147), .B0(H4[26]), .B1(n3140), .Y(n555) );
  INVX1 U1857 ( .A(n554), .Y(n3686) );
  AOI22XL U1858 ( .A0(n2910), .A1(n3146), .B0(H4[22]), .B1(n3139), .Y(n554) );
  INVX1 U1859 ( .A(n548), .Y(n3692) );
  INVX1 U1860 ( .A(n547), .Y(n3693) );
  INVX1 U1861 ( .A(n546), .Y(n3694) );
  INVX1 U1862 ( .A(n544), .Y(n3696) );
  INVX1 U1863 ( .A(n543), .Y(n3697) );
  INVX1 U1864 ( .A(n541), .Y(n3699) );
  INVX1 U1865 ( .A(n540), .Y(n3700) );
  AOI22XL U1866 ( .A0(n3151), .A1(n2901), .B0(H0[22]), .B1(n3138), .Y(n540) );
  INVX1 U1867 ( .A(n539), .Y(n3701) );
  AOI22XL U1868 ( .A0(n2916), .A1(n3145), .B0(H0[26]), .B1(n3138), .Y(n539) );
  INVX1 U1869 ( .A(n538), .Y(n3702) );
  AOI22XL U1870 ( .A0(n3150), .A1(n2888), .B0(H0[24]), .B1(n3138), .Y(n538) );
  INVX1 U1871 ( .A(n497), .Y(n3703) );
  AOI22XL U1872 ( .A0(n3150), .A1(n2862), .B0(H0[28]), .B1(n3138), .Y(n497) );
  INVX1 U1873 ( .A(n496), .Y(n3704) );
  AOI22XL U1874 ( .A0(n3150), .A1(n2682), .B0(H4[31]), .B1(n3138), .Y(n496) );
  INVX1 U1875 ( .A(n625), .Y(n3615) );
  INVX1 U1876 ( .A(n639), .Y(n3601) );
  AOI22XL U1877 ( .A0(n3151), .A1(n2923), .B0(H0[7]), .B1(n3132), .Y(n639) );
  OAI21XL U1878 ( .A0(n3171), .A1(first_block), .B0(n3170), .Y(n447) );
  OAI2BB1X1 U1879 ( .A0N(SHA256_result[208]), .A1N(SHA256_result[176]), .B0(
        n3216), .Y(f2_ABC_32[16]) );
  OAI21XL U1880 ( .A0(SHA256_result[208]), .A1(SHA256_result[176]), .B0(
        SHA256_result[240]), .Y(n3216) );
  OAI211XL U1881 ( .A0(n1161), .A1(n2982), .B0(n3111), .C0(n820), .Y(n2695) );
  AOI22XL U1882 ( .A0(N962), .A1(n2971), .B0(n2830), .B1(n3029), .Y(n820) );
  OAI211XL U1883 ( .A0(n1165), .A1(n2982), .B0(n3111), .C0(n819), .Y(n2699) );
  AOI22XL U1884 ( .A0(N958), .A1(n2967), .B0(n2843), .B1(n3029), .Y(n819) );
  OAI211XL U1885 ( .A0(n1157), .A1(n2982), .B0(n3111), .C0(n821), .Y(n2691) );
  AOI22XL U1886 ( .A0(N966), .A1(n2966), .B0(n2858), .B1(n3029), .Y(n821) );
  OAI211X1 U1887 ( .A0(n2976), .A1(n3858), .B0(n3109), .C0(n737), .Y(n2815) );
  AOI22XL U1888 ( .A0(N843), .A1(n2939), .B0(SHA256_result[240]), .B1(n3033), 
        .Y(n737) );
  OAI211X1 U1889 ( .A0(n2976), .A1(n3859), .B0(n3109), .C0(n751), .Y(n2792) );
  AOI22XL U1890 ( .A0(N865), .A1(n2940), .B0(SHA256_result[198]), .B1(n3032), 
        .Y(n751) );
  OAI211X1 U1891 ( .A0(n2976), .A1(n3544), .B0(n3109), .C0(n753), .Y(n2789) );
  AOI22XL U1892 ( .A0(N868), .A1(n2940), .B0(SHA256_result[201]), .B1(n3031), 
        .Y(n753) );
  OAI211X1 U1893 ( .A0(n2977), .A1(n3531), .B0(n3110), .C0(n761), .Y(n2777) );
  AOI22X1 U1894 ( .A0(N880), .A1(n2940), .B0(SHA256_result[213]), .B1(n3031), 
        .Y(n761) );
  OAI211X1 U1895 ( .A0(n2975), .A1(n3826), .B0(n3108), .C0(n733), .Y(n2821) );
  AOI22XL U1896 ( .A0(N837), .A1(n2972), .B0(SHA256_result[234]), .B1(n3033), 
        .Y(n733) );
  OAI211X1 U1897 ( .A0(n2977), .A1(n3852), .B0(n3110), .C0(n764), .Y(n2771) );
  AOI22X1 U1898 ( .A0(N886), .A1(n2941), .B0(SHA256_result[219]), .B1(n3031), 
        .Y(n764) );
  OAI211XL U1899 ( .A0(n2979), .A1(n3821), .B0(n3112), .C0(n924), .Y(n2497) );
  AOI22X1 U1900 ( .A0(N1001), .A1(n2935), .B0(n3034), .B1(SHA256_result[78]), 
        .Y(n924) );
  OAI211X1 U1901 ( .A0(n2977), .A1(n3860), .B0(n3110), .C0(n762), .Y(n2776) );
  AOI22X1 U1902 ( .A0(N881), .A1(n2940), .B0(SHA256_result[214]), .B1(n3031), 
        .Y(n762) );
  OAI211X1 U1903 ( .A0(n2977), .A1(n3850), .B0(n3110), .C0(n763), .Y(n2772) );
  AOI22X1 U1904 ( .A0(N885), .A1(n2965), .B0(SHA256_result[218]), .B1(n3031), 
        .Y(n763) );
  OAI211X1 U1905 ( .A0(n2977), .A1(n3551), .B0(n3109), .C0(n744), .Y(n2804) );
  AOI22XL U1906 ( .A0(N854), .A1(n2939), .B0(SHA256_result[251]), .B1(n3032), 
        .Y(n744) );
  INVXL U1907 ( .A(SHA256_result[0]), .Y(n3840) );
  INVXL U1908 ( .A(SHA256_result[164]), .Y(n3833) );
  AOI22XL U1909 ( .A0(N863), .A1(n2939), .B0(SHA256_result[196]), .B1(n3032), 
        .Y(n749) );
  INVXL U1910 ( .A(SHA256_result[201]), .Y(n3832) );
  AOI22XL U1911 ( .A0(N836), .A1(n2972), .B0(n2907), .B1(n3033), .Y(n732) );
  INVXL U1912 ( .A(SHA256_result[168]), .Y(n3830) );
  AOI22XL U1913 ( .A0(N867), .A1(n2940), .B0(SHA256_result[200]), .B1(n3032), 
        .Y(n752) );
  INVXL U1914 ( .A(SHA256_result[165]), .Y(n3829) );
  AOI22XL U1915 ( .A0(N864), .A1(n2940), .B0(SHA256_result[197]), .B1(n3032), 
        .Y(n750) );
  OAI211X1 U1916 ( .A0(n2976), .A1(n3828), .B0(n3109), .C0(n754), .Y(n2786) );
  OAI211X1 U1917 ( .A0(n2976), .A1(n3546), .B0(n3109), .C0(n755), .Y(n2785) );
  OAI211X1 U1918 ( .A0(n2976), .A1(n3545), .B0(n3108), .C0(n735), .Y(n2818) );
  AOI22XL U1919 ( .A0(N840), .A1(n2965), .B0(SHA256_result[237]), .B1(n3033), 
        .Y(n735) );
  AOI22XL U1920 ( .A0(N1027), .A1(n2936), .B0(SHA256_result[40]), .B1(n3027), 
        .Y(n937) );
  AOI22XL U1921 ( .A0(N1030), .A1(n2937), .B0(SHA256_result[43]), .B1(n3027), 
        .Y(n939) );
  INVXL U1922 ( .A(SHA256_result[10]), .Y(n3822) );
  AOI22XL U1923 ( .A0(N1029), .A1(n2936), .B0(SHA256_result[42]), .B1(n3027), 
        .Y(n938) );
  AOI22XL U1924 ( .A0(N1033), .A1(n2937), .B0(SHA256_result[46]), .B1(n3027), 
        .Y(n940) );
  OAI211X1 U1925 ( .A0(n2975), .A1(n3541), .B0(n3109), .C0(n738), .Y(n2814) );
  AOI22XL U1926 ( .A0(N844), .A1(n2939), .B0(n2919), .B1(n3033), .Y(n738) );
  OAI211X1 U1927 ( .A0(n2976), .A1(n3539), .B0(n3110), .C0(n758), .Y(n2781) );
  OAI211X1 U1928 ( .A0(n2978), .A1(n3814), .B0(n3109), .C0(n756), .Y(n2784) );
  AOI22XL U1929 ( .A0(N842), .A1(n2966), .B0(SHA256_result[239]), .B1(n3033), 
        .Y(n736) );
  AOI22XL U1930 ( .A0(N892), .A1(n2941), .B0(SHA256_result[161]), .B1(n3030), 
        .Y(n767) );
  OAI211X1 U1931 ( .A0(n2975), .A1(n3537), .B0(n3109), .C0(n739), .Y(n2813) );
  AOI22XL U1932 ( .A0(N845), .A1(n2939), .B0(n2904), .B1(n3033), .Y(n739) );
  OAI211X1 U1933 ( .A0(n2976), .A1(n3536), .B0(n3110), .C0(n759), .Y(n2780) );
  OAI211X1 U1934 ( .A0(n2977), .A1(n3806), .B0(n3110), .C0(n760), .Y(n2779) );
  OAI211X1 U1935 ( .A0(n2981), .A1(n3805), .B0(n3112), .C0(n942), .Y(n2458) );
  AOI22X1 U1936 ( .A0(N1040), .A1(n2937), .B0(SHA256_result[53]), .B1(n3027), 
        .Y(n942) );
  OAI211X1 U1937 ( .A0(n2977), .A1(n3804), .B0(n3110), .C0(n768), .Y(n2763) );
  AOI22XL U1938 ( .A0(N894), .A1(n2941), .B0(SHA256_result[163]), .B1(n3030), 
        .Y(n768) );
  OAI211X1 U1939 ( .A0(n2979), .A1(n3803), .B0(n3110), .C0(n772), .Y(n2756) );
  AOI22XL U1940 ( .A0(N901), .A1(n2941), .B0(SHA256_result[170]), .B1(n3030), 
        .Y(n772) );
  AOI22XL U1941 ( .A0(N896), .A1(n2941), .B0(SHA256_result[165]), .B1(n3030), 
        .Y(n770) );
  OAI211X1 U1942 ( .A0(n2977), .A1(n3801), .B0(n3110), .C0(n769), .Y(n2762) );
  AOI22XL U1943 ( .A0(N895), .A1(n2941), .B0(SHA256_result[164]), .B1(n3030), 
        .Y(n769) );
  OAI211X1 U1944 ( .A0(n2979), .A1(n3799), .B0(n3110), .C0(n771), .Y(n2758) );
  AOI22XL U1945 ( .A0(N899), .A1(n2941), .B0(SHA256_result[168]), .B1(n3030), 
        .Y(n771) );
  OAI211X1 U1946 ( .A0(n2975), .A1(n3533), .B0(n3109), .C0(n741), .Y(n2809) );
  AOI22XL U1947 ( .A0(N849), .A1(n2939), .B0(n2901), .B1(n3033), .Y(n741) );
  OAI211X1 U1948 ( .A0(n2975), .A1(n3532), .B0(n3109), .C0(n740), .Y(n2810) );
  AOI22XL U1949 ( .A0(N848), .A1(n2939), .B0(n2891), .B1(n3033), .Y(n740) );
  OAI211X1 U1950 ( .A0(n2981), .A1(n3791), .B0(n3112), .C0(n946), .Y(n2454) );
  AOI22X1 U1951 ( .A0(N1044), .A1(n2937), .B0(SHA256_result[57]), .B1(n3027), 
        .Y(n946) );
  OAI211X1 U1952 ( .A0(n2981), .A1(n3790), .B0(n3112), .C0(n945), .Y(n2455) );
  AOI22X1 U1953 ( .A0(N1043), .A1(n2937), .B0(SHA256_result[56]), .B1(n3027), 
        .Y(n945) );
  OAI211X1 U1954 ( .A0(n2981), .A1(n3789), .B0(n3112), .C0(n944), .Y(n2456) );
  AOI22X1 U1955 ( .A0(N1042), .A1(n2937), .B0(SHA256_result[55]), .B1(n3027), 
        .Y(n944) );
  OAI211X1 U1956 ( .A0(n2981), .A1(n3788), .B0(n3112), .C0(n943), .Y(n2457) );
  AOI22X1 U1957 ( .A0(N1041), .A1(n2937), .B0(SHA256_result[54]), .B1(n3027), 
        .Y(n943) );
  OAI211X1 U1958 ( .A0(n2978), .A1(n3787), .B0(n3111), .C0(n778), .Y(n2749) );
  OAI211X1 U1959 ( .A0(n2978), .A1(n3786), .B0(n3110), .C0(n775), .Y(n2752) );
  OAI211X1 U1960 ( .A0(n2978), .A1(n3785), .B0(n3110), .C0(n774), .Y(n2753) );
  OAI211X1 U1961 ( .A0(n2978), .A1(n3784), .B0(n3110), .C0(n773), .Y(n2754) );
  OAI211X1 U1962 ( .A0(n2978), .A1(n3781), .B0(n3111), .C0(n777), .Y(n2750) );
  OAI211X1 U1963 ( .A0(n2978), .A1(n3780), .B0(n3110), .C0(n776), .Y(n2751) );
  OAI211X1 U1964 ( .A0(n2980), .A1(n3774), .B0(n3111), .C0(n781), .Y(n2744) );
  AOI22X1 U1965 ( .A0(N913), .A1(n2971), .B0(SHA256_result[182]), .B1(n3029), 
        .Y(n781) );
  OAI211X1 U1966 ( .A0(n2978), .A1(n3773), .B0(n3111), .C0(n780), .Y(n2747) );
  OAI211X1 U1967 ( .A0(n2978), .A1(n3772), .B0(n3111), .C0(n779), .Y(n2748) );
  OAI211X1 U1968 ( .A0(n2980), .A1(n3726), .B0(n3111), .C0(n782), .Y(n2742) );
  AOI22X1 U1969 ( .A0(N915), .A1(n2974), .B0(SHA256_result[184]), .B1(n3029), 
        .Y(n782) );
  INVXL U1970 ( .A(SHA256_result[161]), .Y(n3721) );
  AOI22XL U1971 ( .A0(N860), .A1(n2939), .B0(SHA256_result[193]), .B1(n3032), 
        .Y(n748) );
  OAI2BB1X1 U1972 ( .A0N(SHA256_result[178]), .A1N(SHA256_result[210]), .B0(
        n3214), .Y(f2_ABC_32[18]) );
  OAI21XL U1973 ( .A0(SHA256_result[210]), .A1(SHA256_result[178]), .B0(n2904), 
        .Y(n3214) );
  OAI2BB1X1 U1974 ( .A0N(SHA256_result[177]), .A1N(SHA256_result[209]), .B0(
        n3215), .Y(f2_ABC_32[17]) );
  OAI21XL U1975 ( .A0(SHA256_result[209]), .A1(SHA256_result[177]), .B0(n2919), 
        .Y(n3215) );
  MX2X1 U1976 ( .A(SHA256_result[50]), .B(SHA256_result[82]), .S0(
        SHA256_result[114]), .Y(f1_EFG_32[18]) );
  MX2X1 U1977 ( .A(SHA256_result[51]), .B(SHA256_result[83]), .S0(n2884), .Y(
        n259) );
  MX2X1 U1978 ( .A(SHA256_result[52]), .B(SHA256_result[84]), .S0(n2896), .Y(
        f1_EFG_32[20]) );
  AOI22XL U1979 ( .A0(N971), .A1(n2935), .B0(n2875), .B1(n3028), .Y(n824) );
  INVXL U1980 ( .A(SHA256_result[4]), .Y(n3839) );
  AOI22XL U1981 ( .A0(N1023), .A1(n2936), .B0(SHA256_result[36]), .B1(n3028), 
        .Y(n936) );
  INVXL U1982 ( .A(SHA256_result[3]), .Y(n3838) );
  AOI22XL U1983 ( .A0(N1022), .A1(n2936), .B0(SHA256_result[35]), .B1(n3028), 
        .Y(n935) );
  AOI22XL U1984 ( .A0(N969), .A1(n2935), .B0(n2878), .B1(n3028), .Y(n823) );
  OAI211X1 U1985 ( .A0(n1144), .A1(n2982), .B0(n3111), .C0(n826), .Y(n2678) );
  AOI22XL U1986 ( .A0(N979), .A1(n2935), .B0(n2930), .B1(n3028), .Y(n826) );
  NAND4BXL U1987 ( .AN(n3310), .B(n3309), .C(n3112), .D(n3308), .Y(n2504) );
  NAND2XL U1988 ( .A(SHA256_result[39]), .B(n2988), .Y(n3308) );
  NAND2BX1 U1989 ( .AN(n2956), .B(N994), .Y(n3309) );
  NOR2XL U1990 ( .A(n1161), .B(n3071), .Y(n3310) );
  OAI21XL U1991 ( .A0(n3064), .A1(n3819), .B0(n506), .Y(n1604) );
  AOI22XL U1992 ( .A0(N1031), .A1(n2944), .B0(SHA256_result[12]), .B1(n3156), 
        .Y(n506) );
  OAI21XL U1993 ( .A0(n3063), .A1(n3809), .B0(n504), .Y(n1602) );
  OAI21XL U1994 ( .A0(n3062), .A1(n3810), .B0(n503), .Y(n1601) );
  OAI21XL U1995 ( .A0(n3058), .A1(n3771), .B0(n499), .Y(n1597) );
  AOI22X1 U1996 ( .A0(N1045), .A1(n2943), .B0(SHA256_result[26]), .B1(n3156), 
        .Y(n499) );
  OAI21XL U1997 ( .A0(n3061), .A1(n3858), .B0(n518), .Y(n1616) );
  OAI21XL U1998 ( .A0(n3063), .A1(n3818), .B0(n532), .Y(n1630) );
  AOI22XL U1999 ( .A0(N1000), .A1(n2966), .B0(SHA256_result[45]), .B1(n3157), 
        .Y(n532) );
  OAI21XL U2000 ( .A0(n3055), .A1(n3859), .B0(n490), .Y(n1593) );
  OAI21XL U2001 ( .A0(n3061), .A1(n3792), .B0(n515), .Y(n1613) );
  AOI22X1 U2002 ( .A0(N883), .A1(n2938), .B0(SHA256_result[184]), .B1(n3156), 
        .Y(n515) );
  OAI21XL U2003 ( .A0(n3062), .A1(n3528), .B0(n514), .Y(n1612) );
  AOI22X1 U2004 ( .A0(N884), .A1(n2938), .B0(SHA256_result[185]), .B1(n3156), 
        .Y(n514) );
  OAI21XL U2006 ( .A0(n3056), .A1(n3544), .B0(n488), .Y(n1591) );
  AOI22X1 U2007 ( .A0(N900), .A1(n2935), .B0(SHA256_result[137]), .B1(n3160), 
        .Y(n488) );
  OAI21XL U2008 ( .A0(n3052), .A1(n3531), .B0(n485), .Y(n1588) );
  AOI22X1 U2009 ( .A0(N912), .A1(n2943), .B0(SHA256_result[149]), .B1(n3157), 
        .Y(n485) );
  OAI21XL U2010 ( .A0(n3063), .A1(n3826), .B0(n520), .Y(n1618) );
  AOI22XL U2011 ( .A0(N869), .A1(n2938), .B0(SHA256_result[170]), .B1(n3157), 
        .Y(n520) );
  OAI21XL U2012 ( .A0(n3063), .A1(n3827), .B0(n519), .Y(n1617) );
  AOI22XL U2013 ( .A0(N870), .A1(n2938), .B0(SHA256_result[171]), .B1(n3157), 
        .Y(n519) );
  OAI21XL U2014 ( .A0(n3062), .A1(n3825), .B0(n521), .Y(n1619) );
  AOI22XL U2015 ( .A0(N866), .A1(n2938), .B0(SHA256_result[167]), .B1(n3157), 
        .Y(n521) );
  OAI21XL U2016 ( .A0(n3063), .A1(n3800), .B0(n531), .Y(n1629) );
  OAI21XL U2017 ( .A0(n3063), .A1(n3534), .B0(n517), .Y(n1615) );
  OAI21XL U2018 ( .A0(n3057), .A1(n3529), .B0(n516), .Y(n1614) );
  AOI22X1 U2019 ( .A0(N882), .A1(n2938), .B0(SHA256_result[183]), .B1(n3157), 
        .Y(n516) );
  OAI21XL U2020 ( .A0(n3053), .A1(n3527), .B0(n483), .Y(n1586) );
  AOI22X1 U2021 ( .A0(N916), .A1(n2943), .B0(SHA256_result[153]), .B1(n3159), 
        .Y(n483) );
  OAI21XL U2022 ( .A0(n3056), .A1(n3535), .B0(n486), .Y(n1589) );
  OAI21XL U2023 ( .A0(n3054), .A1(n3530), .B0(n484), .Y(n1587) );
  AOI22X1 U2024 ( .A0(N914), .A1(n2942), .B0(SHA256_result[151]), .B1(n3161), 
        .Y(n484) );
  OAI21XL U2025 ( .A0(n3057), .A1(n3542), .B0(n489), .Y(n1592) );
  INVXL U2026 ( .A(SHA256_result[167]), .Y(n3542) );
  OAI21XL U2027 ( .A0(n3054), .A1(n3543), .B0(n487), .Y(n1590) );
  OAI21XL U2028 ( .A0(n3062), .A1(n3817), .B0(n505), .Y(n1603) );
  INVXL U2029 ( .A(SHA256_result[45]), .Y(n3817) );
  AOI22XL U2030 ( .A0(N1032), .A1(n2943), .B0(SHA256_result[13]), .B1(n3161), 
        .Y(n505) );
  OAI21XL U2031 ( .A0(n3060), .A1(n3798), .B0(n502), .Y(n1600) );
  OAI21XL U2032 ( .A0(n3059), .A1(n3797), .B0(n500), .Y(n1598) );
  INVX1 U2033 ( .A(SHA256_result[52]), .Y(n3797) );
  OAI21XL U2034 ( .A0(n3059), .A1(n3796), .B0(n501), .Y(n1599) );
  OAI21XL U2035 ( .A0(n3064), .A1(n3794), .B0(n529), .Y(n1627) );
  OAI21XL U2036 ( .A0(n3060), .A1(n3795), .B0(n530), .Y(n1628) );
  OAI21XL U2037 ( .A0(n3051), .A1(n3834), .B0(n479), .Y(n1582) );
  INVXL U2038 ( .A(n2906), .Y(n3834) );
  AOI22XL U2039 ( .A0(N828), .A1(n2942), .B0(SHA256_result[193]), .B1(n3157), 
        .Y(n479) );
  OAI21XL U2040 ( .A0(n3055), .A1(n3835), .B0(n453), .Y(n1557) );
  INVXL U2041 ( .A(n2896), .Y(n3835) );
  OAI21XL U2042 ( .A0(n3055), .A1(n3815), .B0(n452), .Y(n1556) );
  INVXL U2043 ( .A(n2915), .Y(n3815) );
  AOI22X1 U2044 ( .A0(N976), .A1(n2943), .B0(SHA256_result[85]), .B1(n3157), 
        .Y(n452) );
  OAI21XL U2045 ( .A0(n3050), .A1(n3836), .B0(n454), .Y(n1558) );
  INVXL U2046 ( .A(n2884), .Y(n3836) );
  NAND2XL U2047 ( .A(SHA256_result[192]), .B(n2989), .Y(n3522) );
  OAI22X1 U2048 ( .A0(n2948), .A1(n3521), .B0(n3050), .B1(n3520), .Y(n3523) );
  INVXL U2049 ( .A(n2933), .Y(n3520) );
  NAND3BX1 U2050 ( .AN(n3489), .B(n3488), .C(n3487), .Y(n1575) );
  NAND2BX1 U2051 ( .AN(n2951), .B(N841), .Y(n3488) );
  NAND2XL U2052 ( .A(SHA256_result[35]), .B(n2987), .Y(n3279) );
  OAI22X1 U2053 ( .A0(n2951), .A1(n3278), .B0(n3046), .B1(n1165), .Y(n3280) );
  NAND2BX1 U2054 ( .AN(n2963), .B(N846), .Y(n3506) );
  NAND2X1 U2055 ( .A(SHA256_result[211]), .B(n3160), .Y(n3505) );
  NAND2BX1 U2056 ( .AN(n2964), .B(N891), .Y(n3492) );
  NAND2XL U2057 ( .A(SHA256_result[128]), .B(n3161), .Y(n3491) );
  NAND2BX1 U2058 ( .AN(n2955), .B(N1026), .Y(n3304) );
  NAND2XL U2059 ( .A(SHA256_result[7]), .B(n3160), .Y(n3303) );
  NAND2BX1 U2060 ( .AN(n2962), .B(N989), .Y(n3177) );
  NAND2XL U2061 ( .A(SHA256_result[34]), .B(n3156), .Y(n3176) );
  NAND2XL U2062 ( .A(SHA256_result[37]), .B(n2985), .Y(n3241) );
  OAI22X1 U2063 ( .A0(n2960), .A1(n3240), .B0(n3040), .B1(n3239), .Y(n3242) );
  INVX1 U2064 ( .A(SHA256_result[69]), .Y(n3239) );
  NAND2BX1 U2065 ( .AN(n2960), .B(N993), .Y(n3256) );
  NAND2XL U2066 ( .A(SHA256_result[38]), .B(n3160), .Y(n3255) );
  NAND2XL U2067 ( .A(SHA256_result[66]), .B(n2990), .Y(n3313) );
  OAI22X1 U2068 ( .A0(n2950), .A1(n3312), .B0(n3043), .B1(n3311), .Y(n3314) );
  INVXL U2069 ( .A(n2844), .Y(n3311) );
  NAND2BX1 U2070 ( .AN(n2959), .B(N1025), .Y(n3323) );
  NAND2XL U2071 ( .A(SHA256_result[6]), .B(n3160), .Y(n3322) );
  NAND2BX1 U2072 ( .AN(n2959), .B(N1021), .Y(n3326) );
  NAND2XL U2073 ( .A(SHA256_result[2]), .B(n3160), .Y(n3325) );
  NAND2BX1 U2074 ( .AN(n2961), .B(N1028), .Y(n3424) );
  NAND2XL U2075 ( .A(SHA256_result[9]), .B(n3158), .Y(n3423) );
  NAND2BX1 U2076 ( .AN(n2964), .B(N996), .Y(n3427) );
  NAND2XL U2077 ( .A(SHA256_result[41]), .B(n3158), .Y(n3426) );
  NAND2BX1 U2078 ( .AN(n2961), .B(N1024), .Y(n3320) );
  NAND2XL U2079 ( .A(SHA256_result[5]), .B(n3160), .Y(n3319) );
  NAND2XL U2080 ( .A(SHA256_result[40]), .B(n2988), .Y(n3306) );
  OAI22X1 U2081 ( .A0(n2950), .A1(n3305), .B0(n3047), .B1(n2401), .Y(n3307) );
  NAND2XL U2082 ( .A(SHA256_result[194]), .B(n2988), .Y(n3174) );
  OAI22X1 U2083 ( .A0(n2949), .A1(n3173), .B0(n3042), .B1(n3172), .Y(n3175) );
  INVXL U2084 ( .A(n2892), .Y(n3172) );
  NAND2BX1 U2085 ( .AN(n2957), .B(N1020), .Y(n3317) );
  NAND2XL U2086 ( .A(SHA256_result[1]), .B(n3160), .Y(n3316) );
  NAND2XL U2087 ( .A(n2685), .B(n2988), .Y(n3180) );
  OAI22X1 U2088 ( .A0(n2948), .A1(n3179), .B0(n3039), .B1(n3178), .Y(n3181) );
  INVX1 U2089 ( .A(n3722), .Y(n3178) );
  NAND3X1 U2090 ( .A(n3415), .B(n3414), .C(n3413), .Y(n1579) );
  NAND2BX1 U2091 ( .AN(n2962), .B(N832), .Y(n3415) );
  NAND2BXL U2092 ( .AN(n3050), .B(n2928), .Y(n3414) );
  NAND2XL U2093 ( .A(SHA256_result[197]), .B(n3158), .Y(n3413) );
  NAND3X1 U2094 ( .A(n3515), .B(n3514), .C(n3513), .Y(n1622) );
  NAND2BX1 U2095 ( .AN(n2964), .B(N859), .Y(n3515) );
  NAND2BXL U2096 ( .AN(n3045), .B(SHA256_result[192]), .Y(n3514) );
  NAND2XL U2097 ( .A(SHA256_result[160]), .B(n3158), .Y(n3513) );
  NAND3X1 U2098 ( .A(n3418), .B(n3417), .C(n3416), .Y(n1578) );
  NAND2BX1 U2099 ( .AN(n2962), .B(N833), .Y(n3418) );
  NAND2BXL U2100 ( .AN(n3049), .B(n2924), .Y(n3417) );
  NAND2XL U2101 ( .A(SHA256_result[198]), .B(n3158), .Y(n3416) );
  NAND3X1 U2102 ( .A(n3253), .B(n3252), .C(n3251), .Y(n1567) );
  NAND2BX1 U2103 ( .AN(n2952), .B(N959), .Y(n3253) );
  NAND2BXL U2104 ( .AN(n3058), .B(n2837), .Y(n3252) );
  NAND2XL U2105 ( .A(SHA256_result[68]), .B(n3161), .Y(n3251) );
  NAND3X1 U2106 ( .A(n3262), .B(n3261), .C(n3260), .Y(n1565) );
  NAND2BX1 U2107 ( .AN(n2958), .B(N961), .Y(n3262) );
  NAND2BXL U2108 ( .AN(n3056), .B(n2833), .Y(n3261) );
  NAND2XL U2109 ( .A(SHA256_result[70]), .B(n3160), .Y(n3260) );
  NAND3X1 U2110 ( .A(n3421), .B(n3420), .C(n3419), .Y(n1621) );
  NAND2BX1 U2111 ( .AN(n2962), .B(N861), .Y(n3421) );
  NAND2BXL U2112 ( .AN(n3054), .B(SHA256_result[194]), .Y(n3420) );
  NAND2XL U2113 ( .A(SHA256_result[162]), .B(n3158), .Y(n3419) );
  NAND3X1 U2114 ( .A(n3430), .B(n3429), .C(n3428), .Y(n1562) );
  NAND2BX1 U2115 ( .AN(n2950), .B(N965), .Y(n3430) );
  NAND2BXL U2116 ( .AN(n3047), .B(n2867), .Y(n3429) );
  NAND2XL U2117 ( .A(SHA256_result[74]), .B(n3158), .Y(n3428) );
  NAND3X1 U2118 ( .A(n3433), .B(n3432), .C(n3431), .Y(n1563) );
  NAND2BX1 U2119 ( .AN(n2961), .B(N964), .Y(n3433) );
  NAND2BXL U2120 ( .AN(n3046), .B(n2869), .Y(n3432) );
  NAND2XL U2121 ( .A(SHA256_result[73]), .B(n3158), .Y(n3431) );
  NAND3X1 U2122 ( .A(n3495), .B(n3494), .C(n3493), .Y(n1594) );
  NAND2BX1 U2123 ( .AN(n2961), .B(N893), .Y(n3495) );
  NAND2BXL U2124 ( .AN(n3041), .B(SHA256_result[162]), .Y(n3494) );
  NAND2XL U2125 ( .A(SHA256_result[130]), .B(n3161), .Y(n3493) );
  NAND3X1 U2126 ( .A(n3509), .B(n3508), .C(n3507), .Y(n1555) );
  NAND2BXL U2127 ( .AN(n3054), .B(n2910), .Y(n3508) );
  NAND2BX1 U2128 ( .AN(n2963), .B(N977), .Y(n3509) );
  NAND2X1 U2129 ( .A(SHA256_result[86]), .B(n3158), .Y(n3507) );
  OAI2BB1X1 U2130 ( .A0N(n3038), .A1N(n2920), .B0(n474), .Y(n1577) );
  AOI22XL U2131 ( .A0(N835), .A1(n2944), .B0(SHA256_result[200]), .B1(n3161), 
        .Y(n474) );
  OAI2BB1X1 U2132 ( .A0N(n3038), .A1N(n2929), .B0(n477), .Y(n1580) );
  AOI22XL U2133 ( .A0(N831), .A1(n2943), .B0(SHA256_result[196]), .B1(n3161), 
        .Y(n477) );
  OAI2BB1X1 U2134 ( .A0N(n3037), .A1N(SHA256_result[195]), .B0(n522), .Y(n1620) );
  AOI22XL U2135 ( .A0(N862), .A1(n2938), .B0(SHA256_result[163]), .B1(n3157), 
        .Y(n522) );
  OAI2BB1X1 U2136 ( .A0N(n3037), .A1N(SHA256_result[85]), .B0(n528), .Y(n1626)
         );
  INVX1 U2137 ( .A(N804), .Y(n3442) );
  OAI2BB1X1 U2138 ( .A0N(n3038), .A1N(SHA256_result[74]), .B0(n533), .Y(n1631)
         );
  AOI22XL U2139 ( .A0(N997), .A1(n2971), .B0(SHA256_result[42]), .B1(n3157), 
        .Y(n533) );
  INVX1 U2140 ( .A(N805), .Y(n3438) );
  OAI2BB1X1 U2141 ( .A0N(n3037), .A1N(SHA256_result[86]), .B0(n527), .Y(n1625)
         );
  OAI2BB1X1 U2142 ( .A0N(n3037), .A1N(SHA256_result[236]), .B0(n473), .Y(n1576) );
  OAI2BB1X1 U2143 ( .A0N(n3038), .A1N(SHA256_result[244]), .B0(n470), .Y(n1573) );
  OAI2BB1X1 U2144 ( .A0N(n3037), .A1N(n2903), .B0(n469), .Y(n1572) );
  OAI2BB1X1 U2145 ( .A0N(n3037), .A1N(n2905), .B0(n478), .Y(n1581) );
  AOI22XL U2146 ( .A0(N830), .A1(n2942), .B0(SHA256_result[195]), .B1(n3161), 
        .Y(n478) );
  OAI2BB1X1 U2147 ( .A0N(n3037), .A1N(n2916), .B0(n468), .Y(n1571) );
  AOI22X1 U2148 ( .A0(N853), .A1(n2943), .B0(SHA256_result[218]), .B1(n3157), 
        .Y(n468) );
  OAI2BB1X1 U2149 ( .A0N(n3038), .A1N(SHA256_result[68]), .B0(n536), .Y(n1634)
         );
  AOI22XL U2150 ( .A0(N991), .A1(n2966), .B0(SHA256_result[36]), .B1(n3157), 
        .Y(n536) );
  BUFX3 U2151 ( .A(n677), .Y(n2828) );
  NAND3BXL U2152 ( .AN(n3171), .B(first_block), .C(n3170), .Y(n677) );
  MX2X1 U2153 ( .A(SHA256_result[53]), .B(SHA256_result[85]), .S0(n2915), .Y(
        n287) );
  MX2X1 U2154 ( .A(SHA256_result[54]), .B(SHA256_result[86]), .S0(n2910), .Y(
        n265) );
  MXI2XL U2155 ( .A(n3793), .B(n1145), .S0(n2909), .Y(f1_EFG_32[23]) );
  OAI2BB1X1 U2156 ( .A0N(SHA256_result[179]), .A1N(SHA256_result[211]), .B0(
        n3213), .Y(f2_ABC_32[19]) );
  OAI21XL U2157 ( .A0(SHA256_result[179]), .A1(SHA256_result[211]), .B0(
        SHA256_result[243]), .Y(n3213) );
  OAI2BB1X1 U2158 ( .A0N(SHA256_result[212]), .A1N(SHA256_result[180]), .B0(
        n3212), .Y(f2_ABC_32[20]) );
  OAI21XL U2159 ( .A0(SHA256_result[180]), .A1(SHA256_result[212]), .B0(
        SHA256_result[244]), .Y(n3212) );
  NAND2X1 U2160 ( .A(n1078), .B(read_counter[0]), .Y(N3079) );
  AOI22XL U2161 ( .A0(n3096), .A1(SHA256_result[193]), .B0(n3093), .B1(n2906), 
        .Y(n1229) );
  AOI22XL U2162 ( .A0(n3096), .A1(SHA256_result[196]), .B0(n3093), .B1(n2929), 
        .Y(n1217) );
  AOI22XL U2163 ( .A0(n3096), .A1(SHA256_result[200]), .B0(n3093), .B1(n2920), 
        .Y(n1201) );
  AOI22XL U2164 ( .A0(n3097), .A1(SHA256_result[206]), .B0(n3094), .B1(
        SHA256_result[238]), .Y(n1177) );
  AOI22XL U2165 ( .A0(n3097), .A1(SHA256_result[210]), .B0(n3094), .B1(n2904), 
        .Y(n1149) );
  AOI22XL U2166 ( .A0(n3096), .A1(SHA256_result[197]), .B0(n3093), .B1(n2928), 
        .Y(n1213) );
  AOI22XL U2167 ( .A0(n3097), .A1(SHA256_result[207]), .B0(n3094), .B1(
        SHA256_result[239]), .Y(n1173) );
  AOI22XL U2168 ( .A0(n3097), .A1(SHA256_result[209]), .B0(n3094), .B1(n2919), 
        .Y(n1159) );
  AOI22XL U2169 ( .A0(n3096), .A1(SHA256_result[201]), .B0(n3093), .B1(n2907), 
        .Y(n1197) );
  AOI22XL U2170 ( .A0(n3097), .A1(SHA256_result[208]), .B0(n3094), .B1(
        SHA256_result[240]), .Y(n1169) );
  AOI22XL U2171 ( .A0(n3096), .A1(SHA256_result[198]), .B0(n3093), .B1(n2924), 
        .Y(n1209) );
  AOI22XL U2172 ( .A0(n3097), .A1(SHA256_result[204]), .B0(n3094), .B1(
        SHA256_result[236]), .Y(n1185) );
  AOI22XL U2173 ( .A0(n3097), .A1(SHA256_result[211]), .B0(n3094), .B1(
        SHA256_result[243]), .Y(n1139) );
  AOI22XL U2174 ( .A0(n3097), .A1(SHA256_result[213]), .B0(n3094), .B1(n2891), 
        .Y(n1131) );
  AOI22XL U2175 ( .A0(n3097), .A1(SHA256_result[212]), .B0(n3094), .B1(
        SHA256_result[244]), .Y(n1135) );
  AOI22XL U2176 ( .A0(n3097), .A1(SHA256_result[215]), .B0(n3094), .B1(n2903), 
        .Y(n1123) );
  AOI22XL U2177 ( .A0(n3097), .A1(SHA256_result[205]), .B0(n3094), .B1(
        SHA256_result[237]), .Y(n1181) );
  AOI22XL U2178 ( .A0(n3106), .A1(SHA256_result[93]), .B0(n3104), .B1(n2860), 
        .Y(n1102) );
  AOI22XL U2179 ( .A0(n3106), .A1(SHA256_result[94]), .B0(n3104), .B1(n2871), 
        .Y(n1098) );
  AOI22XL U2180 ( .A0(n3097), .A1(SHA256_result[214]), .B0(n3094), .B1(n2901), 
        .Y(n1127) );
  AOI22XL U2181 ( .A0(n3096), .A1(SHA256_result[195]), .B0(n3093), .B1(n2905), 
        .Y(n1221) );
  AOI22XL U2182 ( .A0(n3096), .A1(SHA256_result[194]), .B0(n3093), .B1(n2892), 
        .Y(n1225) );
  AOI22XL U2183 ( .A0(n3106), .A1(SHA256_result[95]), .B0(n3104), .B1(n2682), 
        .Y(n1086) );
  AOI22XL U2184 ( .A0(n3096), .A1(SHA256_result[199]), .B0(n3093), .B1(n2923), 
        .Y(n1205) );
  AOI22XL U2185 ( .A0(n3096), .A1(SHA256_result[202]), .B0(n3093), .B1(
        SHA256_result[234]), .Y(n1193) );
  AOI22XL U2186 ( .A0(n3096), .A1(SHA256_result[203]), .B0(n3093), .B1(
        SHA256_result[235]), .Y(n1189) );
  NAND4X1 U2187 ( .A(n1233), .B(n1234), .C(n1235), .D(n1236), .Y(N3047) );
  AOI22XL U2188 ( .A0(n3099), .A1(SHA256_result[128]), .B0(n1092), .B1(
        SHA256_result[160]), .Y(n1234) );
  AOI22XL U2189 ( .A0(n3096), .A1(SHA256_result[192]), .B0(n3093), .B1(n2933), 
        .Y(n1233) );
  NAND4X1 U2190 ( .A(n1209), .B(n1210), .C(n1211), .D(n1212), .Y(N3053) );
  AOI22XL U2191 ( .A0(n3099), .A1(SHA256_result[134]), .B0(n1092), .B1(
        SHA256_result[166]), .Y(n1210) );
  AOI22XL U2192 ( .A0(n3103), .A1(SHA256_result[6]), .B0(n3101), .B1(
        SHA256_result[38]), .Y(n1211) );
  AOI22XL U2193 ( .A0(n3107), .A1(SHA256_result[70]), .B0(n3105), .B1(n2833), 
        .Y(n1212) );
  NAND4X1 U2194 ( .A(n1181), .B(n1182), .C(n1183), .D(n1184), .Y(N3060) );
  AOI22XL U2195 ( .A0(n3103), .A1(SHA256_result[13]), .B0(n3101), .B1(
        SHA256_result[45]), .Y(n1183) );
  AOI22XL U2196 ( .A0(n3107), .A1(SHA256_result[77]), .B0(n3105), .B1(n2873), 
        .Y(n1184) );
  NAND4X1 U2197 ( .A(n1139), .B(n1146), .C(n1147), .D(n1148), .Y(N3066) );
  AOI22X1 U2198 ( .A0(n3099), .A1(SHA256_result[147]), .B0(n1092), .B1(
        SHA256_result[179]), .Y(n1146) );
  AOI22XL U2199 ( .A0(n3106), .A1(SHA256_result[83]), .B0(n3105), .B1(n2884), 
        .Y(n1148) );
  NAND4X1 U2200 ( .A(n1135), .B(n1136), .C(n1137), .D(n1138), .Y(N3067) );
  AOI22X1 U2201 ( .A0(n3098), .A1(SHA256_result[148]), .B0(n1092), .B1(
        SHA256_result[180]), .Y(n1136) );
  AOI22X1 U2202 ( .A0(n3102), .A1(SHA256_result[20]), .B0(n3100), .B1(
        SHA256_result[52]), .Y(n1137) );
  AOI22XL U2203 ( .A0(n3106), .A1(SHA256_result[84]), .B0(n3104), .B1(n2896), 
        .Y(n1138) );
  NAND4X1 U2204 ( .A(n1131), .B(n1132), .C(n1133), .D(n1134), .Y(N3068) );
  AOI22X1 U2205 ( .A0(n3098), .A1(SHA256_result[149]), .B0(n1092), .B1(
        SHA256_result[181]), .Y(n1132) );
  AOI22X1 U2206 ( .A0(n3102), .A1(SHA256_result[21]), .B0(n3100), .B1(
        SHA256_result[53]), .Y(n1133) );
  AOI22XL U2207 ( .A0(n3106), .A1(SHA256_result[85]), .B0(n3104), .B1(n2915), 
        .Y(n1134) );
  NAND4X1 U2208 ( .A(n1099), .B(n1100), .C(n1101), .D(n1102), .Y(N3076) );
  AOI22X1 U2209 ( .A0(n3098), .A1(SHA256_result[157]), .B0(n1092), .B1(
        SHA256_result[189]), .Y(n1100) );
  AOI22XL U2210 ( .A0(n3096), .A1(SHA256_result[221]), .B0(n3093), .B1(n2849), 
        .Y(n1099) );
  AOI22X1 U2211 ( .A0(n3102), .A1(SHA256_result[29]), .B0(n3100), .B1(
        SHA256_result[61]), .Y(n1101) );
  NAND4X1 U2212 ( .A(n1095), .B(n1096), .C(n1097), .D(n1098), .Y(N3077) );
  AOI22X1 U2213 ( .A0(n3098), .A1(SHA256_result[158]), .B0(n1092), .B1(
        SHA256_result[190]), .Y(n1096) );
  AOI22XL U2214 ( .A0(n3097), .A1(SHA256_result[222]), .B0(n1094), .B1(n2855), 
        .Y(n1095) );
  AOI22X1 U2215 ( .A0(n3102), .A1(SHA256_result[30]), .B0(n3100), .B1(
        SHA256_result[62]), .Y(n1097) );
  NAND4X1 U2216 ( .A(n1217), .B(n1218), .C(n1219), .D(n1220), .Y(N3051) );
  AOI22XL U2217 ( .A0(n3099), .A1(SHA256_result[132]), .B0(n1092), .B1(
        SHA256_result[164]), .Y(n1218) );
  AOI22XL U2218 ( .A0(n3103), .A1(SHA256_result[4]), .B0(n3100), .B1(
        SHA256_result[36]), .Y(n1219) );
  AOI22XL U2219 ( .A0(n3107), .A1(SHA256_result[68]), .B0(n3104), .B1(n2837), 
        .Y(n1220) );
  NAND4X1 U2220 ( .A(n1193), .B(n1194), .C(n1195), .D(n1196), .Y(N3057) );
  AOI22XL U2221 ( .A0(n3099), .A1(SHA256_result[138]), .B0(n1092), .B1(
        SHA256_result[170]), .Y(n1194) );
  AOI22XL U2222 ( .A0(n3103), .A1(SHA256_result[10]), .B0(n3101), .B1(
        SHA256_result[42]), .Y(n1195) );
  AOI22XL U2223 ( .A0(n3107), .A1(SHA256_result[74]), .B0(n3105), .B1(n2867), 
        .Y(n1196) );
  NAND4X1 U2224 ( .A(n1127), .B(n1128), .C(n1129), .D(n1130), .Y(N3069) );
  AOI22X1 U2225 ( .A0(n3098), .A1(SHA256_result[150]), .B0(n1092), .B1(
        SHA256_result[182]), .Y(n1128) );
  AOI22X1 U2226 ( .A0(n3102), .A1(SHA256_result[22]), .B0(n3100), .B1(
        SHA256_result[54]), .Y(n1129) );
  AOI22XL U2227 ( .A0(n3106), .A1(SHA256_result[86]), .B0(n3104), .B1(n2910), 
        .Y(n1130) );
  NAND4X1 U2228 ( .A(n1197), .B(n1198), .C(n1199), .D(n1200), .Y(N3056) );
  AOI22XL U2229 ( .A0(n3099), .A1(SHA256_result[137]), .B0(n1092), .B1(
        SHA256_result[169]), .Y(n1198) );
  AOI22XL U2230 ( .A0(n3103), .A1(SHA256_result[9]), .B0(n3101), .B1(
        SHA256_result[41]), .Y(n1199) );
  AOI22XL U2231 ( .A0(n3106), .A1(SHA256_result[73]), .B0(n3105), .B1(n2869), 
        .Y(n1200) );
  NAND4X1 U2232 ( .A(n1225), .B(n1226), .C(n1227), .D(n1228), .Y(N3049) );
  AOI22XL U2233 ( .A0(n3098), .A1(SHA256_result[130]), .B0(n1092), .B1(
        SHA256_result[162]), .Y(n1226) );
  AOI22XL U2234 ( .A0(n3103), .A1(SHA256_result[2]), .B0(n3101), .B1(
        SHA256_result[34]), .Y(n1227) );
  AOI22XL U2235 ( .A0(n3107), .A1(SHA256_result[66]), .B0(n3105), .B1(n2844), 
        .Y(n1228) );
  NAND4X1 U2236 ( .A(n1206), .B(n1207), .C(n1205), .D(n3277), .Y(N3054) );
  AOI22XL U2237 ( .A0(n3098), .A1(SHA256_result[135]), .B0(n1092), .B1(
        SHA256_result[167]), .Y(n1206) );
  AOI22XL U2238 ( .A0(n3103), .A1(SHA256_result[7]), .B0(n3101), .B1(
        SHA256_result[39]), .Y(n1207) );
  AOI21X1 U2239 ( .A0(n3107), .A1(SHA256_result[71]), .B0(n3276), .Y(n3277) );
  NAND4X1 U2240 ( .A(n1083), .B(n1084), .C(n1085), .D(n1086), .Y(N3078) );
  AOI22X1 U2241 ( .A0(n3098), .A1(SHA256_result[159]), .B0(n1092), .B1(
        SHA256_result[191]), .Y(n1084) );
  AOI22XL U2242 ( .A0(n3097), .A1(SHA256_result[223]), .B0(n3094), .B1(n2887), 
        .Y(n1083) );
  AOI22X1 U2243 ( .A0(n3102), .A1(SHA256_result[31]), .B0(n3100), .B1(
        SHA256_result[63]), .Y(n1085) );
  NAND4X1 U2244 ( .A(n1149), .B(n1150), .C(n1155), .D(n1158), .Y(N3065) );
  AOI22X1 U2245 ( .A0(n3099), .A1(SHA256_result[146]), .B0(n1092), .B1(
        SHA256_result[178]), .Y(n1150) );
  AOI22XL U2246 ( .A0(n3107), .A1(SHA256_result[82]), .B0(n3105), .B1(
        SHA256_result[114]), .Y(n1158) );
  NAND4X1 U2247 ( .A(n1221), .B(n1222), .C(n1223), .D(n1224), .Y(N3050) );
  AOI22XL U2248 ( .A0(n3099), .A1(SHA256_result[131]), .B0(n1092), .B1(
        SHA256_result[163]), .Y(n1222) );
  AOI22XL U2249 ( .A0(n3103), .A1(SHA256_result[3]), .B0(n3100), .B1(
        SHA256_result[35]), .Y(n1223) );
  AOI22XL U2250 ( .A0(n3107), .A1(SHA256_result[67]), .B0(n3104), .B1(n2843), 
        .Y(n1224) );
  NAND4X1 U2251 ( .A(n1213), .B(n1214), .C(n1215), .D(n1216), .Y(N3052) );
  AOI22XL U2252 ( .A0(n3098), .A1(SHA256_result[133]), .B0(n1092), .B1(
        SHA256_result[165]), .Y(n1214) );
  AOI22XL U2253 ( .A0(n3103), .A1(SHA256_result[5]), .B0(n3101), .B1(
        SHA256_result[37]), .Y(n1215) );
  AOI22XL U2254 ( .A0(n3107), .A1(SHA256_result[69]), .B0(n3104), .B1(n2840), 
        .Y(n1216) );
  NAND4X1 U2255 ( .A(n1229), .B(n1230), .C(n1231), .D(n1232), .Y(N3048) );
  AOI22XL U2256 ( .A0(n3098), .A1(SHA256_result[129]), .B0(n1092), .B1(
        SHA256_result[161]), .Y(n1230) );
  AOI22XL U2257 ( .A0(n3103), .A1(SHA256_result[1]), .B0(n3100), .B1(n2685), 
        .Y(n1231) );
  AOI22XL U2258 ( .A0(n3107), .A1(n3722), .B0(n3105), .B1(n2851), .Y(n1232) );
  NAND4X1 U2259 ( .A(n1201), .B(n1202), .C(n1203), .D(n1204), .Y(N3055) );
  AOI22XL U2260 ( .A0(n3099), .A1(SHA256_result[136]), .B0(n1092), .B1(
        SHA256_result[168]), .Y(n1202) );
  AOI22XL U2261 ( .A0(n3102), .A1(SHA256_result[8]), .B0(n3101), .B1(
        SHA256_result[40]), .Y(n1203) );
  AOI22XL U2262 ( .A0(n3106), .A1(SHA256_result[72]), .B0(n3105), .B1(
        SHA256_result[104]), .Y(n1204) );
  NAND4X1 U2263 ( .A(n1189), .B(n1190), .C(n1191), .D(n1192), .Y(N3058) );
  AOI22XL U2264 ( .A0(n3099), .A1(SHA256_result[139]), .B0(n1092), .B1(
        SHA256_result[171]), .Y(n1190) );
  AOI22XL U2265 ( .A0(n3103), .A1(SHA256_result[11]), .B0(n3101), .B1(
        SHA256_result[43]), .Y(n1191) );
  AOI22XL U2266 ( .A0(n3107), .A1(SHA256_result[75]), .B0(n3105), .B1(n2858), 
        .Y(n1192) );
  NAND4X1 U2267 ( .A(n1185), .B(n1186), .C(n1187), .D(n1188), .Y(N3059) );
  AOI22XL U2268 ( .A0(n3102), .A1(SHA256_result[12]), .B0(n3101), .B1(
        SHA256_result[44]), .Y(n1187) );
  AOI22XL U2269 ( .A0(n3106), .A1(SHA256_result[76]), .B0(n3105), .B1(n2859), 
        .Y(n1188) );
  NAND4X1 U2270 ( .A(n1177), .B(n1178), .C(n1179), .D(n1180), .Y(N3061) );
  AOI22XL U2271 ( .A0(n3102), .A1(SHA256_result[14]), .B0(n3101), .B1(
        SHA256_result[46]), .Y(n1179) );
  AOI22XL U2272 ( .A0(n3107), .A1(SHA256_result[78]), .B0(n3105), .B1(n2878), 
        .Y(n1180) );
  NAND4X1 U2273 ( .A(n1173), .B(n1174), .C(n1175), .D(n1176), .Y(N3062) );
  AOI22XL U2274 ( .A0(n3107), .A1(n3808), .B0(n3105), .B1(n2872), .Y(n1176) );
  NAND4X1 U2275 ( .A(n1169), .B(n1170), .C(n1171), .D(n1172), .Y(N3063) );
  AOI22X1 U2276 ( .A0(n3099), .A1(SHA256_result[144]), .B0(n1092), .B1(
        SHA256_result[176]), .Y(n1170) );
  AOI22XL U2277 ( .A0(n3107), .A1(SHA256_result[80]), .B0(n3105), .B1(n2875), 
        .Y(n1172) );
  NAND4X1 U2278 ( .A(n1159), .B(n1162), .C(n1164), .D(n1166), .Y(N3064) );
  AOI22X1 U2279 ( .A0(n3099), .A1(SHA256_result[145]), .B0(n1092), .B1(
        SHA256_result[177]), .Y(n1162) );
  AOI22XL U2280 ( .A0(n3107), .A1(n3807), .B0(n3105), .B1(n2899), .Y(n1166) );
  NAND4X1 U2281 ( .A(n1119), .B(n1120), .C(n1121), .D(n1122), .Y(N3071) );
  AOI22X1 U2282 ( .A0(n3098), .A1(SHA256_result[152]), .B0(n1092), .B1(
        SHA256_result[184]), .Y(n1120) );
  AOI22XL U2283 ( .A0(n3097), .A1(SHA256_result[216]), .B0(n1094), .B1(n2888), 
        .Y(n1119) );
  AOI22X1 U2284 ( .A0(n3102), .A1(SHA256_result[24]), .B0(n3100), .B1(
        SHA256_result[56]), .Y(n1121) );
  NAND4X1 U2285 ( .A(n1115), .B(n1116), .C(n1117), .D(n1118), .Y(N3072) );
  AOI22X1 U2286 ( .A0(n3098), .A1(SHA256_result[153]), .B0(n1092), .B1(
        SHA256_result[185]), .Y(n1116) );
  AOI22XL U2287 ( .A0(n3096), .A1(SHA256_result[217]), .B0(n1094), .B1(n2857), 
        .Y(n1115) );
  AOI22X1 U2288 ( .A0(n3102), .A1(SHA256_result[25]), .B0(n3100), .B1(
        SHA256_result[57]), .Y(n1117) );
  NAND4X1 U2289 ( .A(n1111), .B(n1112), .C(n1113), .D(n1114), .Y(N3073) );
  AOI22X1 U2290 ( .A0(n3098), .A1(SHA256_result[154]), .B0(n1092), .B1(
        SHA256_result[186]), .Y(n1112) );
  AOI22XL U2291 ( .A0(n3096), .A1(SHA256_result[218]), .B0(n1094), .B1(n2916), 
        .Y(n1111) );
  AOI22X1 U2292 ( .A0(n3102), .A1(SHA256_result[26]), .B0(n3100), .B1(
        SHA256_result[58]), .Y(n1113) );
  NAND4X1 U2293 ( .A(n1107), .B(n1108), .C(n1109), .D(n1110), .Y(N3074) );
  AOI22X1 U2294 ( .A0(n3098), .A1(SHA256_result[155]), .B0(n1092), .B1(
        SHA256_result[187]), .Y(n1108) );
  AOI22XL U2295 ( .A0(n3096), .A1(SHA256_result[219]), .B0(n1094), .B1(
        SHA256_result[251]), .Y(n1107) );
  AOI22X1 U2296 ( .A0(n3102), .A1(SHA256_result[27]), .B0(n3100), .B1(
        SHA256_result[59]), .Y(n1109) );
  NAND4X1 U2297 ( .A(n1103), .B(n1104), .C(n1105), .D(n1106), .Y(N3075) );
  AOI22X1 U2298 ( .A0(n3098), .A1(SHA256_result[156]), .B0(n1092), .B1(
        SHA256_result[188]), .Y(n1104) );
  AOI22XL U2299 ( .A0(n3097), .A1(SHA256_result[220]), .B0(n3094), .B1(n2862), 
        .Y(n1103) );
  AOI22X1 U2300 ( .A0(n3102), .A1(SHA256_result[28]), .B0(n3100), .B1(
        SHA256_result[60]), .Y(n1105) );
  NAND4X1 U2301 ( .A(n1123), .B(n1124), .C(n1125), .D(n1126), .Y(N3070) );
  AOI22X1 U2302 ( .A0(n3098), .A1(SHA256_result[151]), .B0(n1092), .B1(
        SHA256_result[183]), .Y(n1124) );
  AOI22X1 U2303 ( .A0(n3102), .A1(SHA256_result[23]), .B0(n3100), .B1(
        SHA256_result[55]), .Y(n1125) );
  AOI22XL U2304 ( .A0(n3106), .A1(SHA256_result[87]), .B0(n3104), .B1(n2909), 
        .Y(n1126) );
  AND3X2 U2305 ( .A(n1078), .B(read_counter[2]), .C(n1081), .Y(n1092) );
  NOR3XL U2306 ( .A(n656), .B(round[6]), .C(output_enable), .Y(n40) );
  MXI2XL U2307 ( .A(n3782), .B(n1144), .S0(n2930), .Y(f1_EFG_32[24]) );
  MXI2XL U2308 ( .A(n3783), .B(n1143), .S0(n2883), .Y(f1_EFG_32[25]) );
  MXI2XL U2309 ( .A(n3771), .B(n1142), .S0(n2877), .Y(f1_EFG_32[26]) );
  OAI2BB1X1 U2310 ( .A0N(n2901), .A1N(SHA256_result[214]), .B0(n3210), .Y(
        f2_ABC_32[22]) );
  OAI21XL U2311 ( .A0(n2901), .A1(SHA256_result[214]), .B0(SHA256_result[182]), 
        .Y(n3210) );
  OAI2BB1X1 U2312 ( .A0N(SHA256_result[215]), .A1N(SHA256_result[183]), .B0(
        n3209), .Y(f2_ABC_32[23]) );
  OAI21XL U2313 ( .A0(SHA256_result[183]), .A1(SHA256_result[215]), .B0(n2903), 
        .Y(n3209) );
  OAI2BB1X1 U2314 ( .A0N(SHA256_result[213]), .A1N(SHA256_result[181]), .B0(
        n3211), .Y(f2_ABC_32[21]) );
  OAI21XL U2315 ( .A0(SHA256_result[213]), .A1(SHA256_result[181]), .B0(n2891), 
        .Y(n3211) );
  BUFX3 U2316 ( .A(n995), .Y(n2932) );
  OAI21XL U2317 ( .A0(n1081), .A1(n1082), .B0(n1078), .Y(N3080) );
  NOR2X1 U2318 ( .A(read_counter[0]), .B(n3725), .Y(n1082) );
  INVX1 U2319 ( .A(N926), .Y(n3244) );
  MXI2XL U2320 ( .A(n3856), .B(n1141), .S0(n2864), .Y(f1_EFG_32[27]) );
  MXI2XL U2321 ( .A(n3855), .B(n1140), .S0(n2874), .Y(f1_EFG_32[28]) );
  OAI2BB1X1 U2322 ( .A0N(SHA256_result[186]), .A1N(n2916), .B0(n3206), .Y(
        f2_ABC_32[26]) );
  OAI21XL U2323 ( .A0(SHA256_result[186]), .A1(n2916), .B0(SHA256_result[218]), 
        .Y(n3206) );
  OAI2BB1X1 U2324 ( .A0N(SHA256_result[216]), .A1N(SHA256_result[184]), .B0(
        n3208), .Y(f2_ABC_32[24]) );
  OAI21XL U2325 ( .A0(SHA256_result[216]), .A1(SHA256_result[184]), .B0(n2888), 
        .Y(n3208) );
  OAI2BB1X1 U2326 ( .A0N(SHA256_result[217]), .A1N(SHA256_result[185]), .B0(
        n3207), .Y(f2_ABC_32[25]) );
  OAI21XL U2327 ( .A0(SHA256_result[185]), .A1(SHA256_result[217]), .B0(n2857), 
        .Y(n3207) );
  MX2X1 U2328 ( .A(SHA256_result[61]), .B(SHA256_result[93]), .S0(n2860), .Y(
        f1_EFG_32[29]) );
  INVX1 U2329 ( .A(N924), .Y(n3273) );
  INVX1 U2330 ( .A(N796), .Y(n3410) );
  INVX1 U2331 ( .A(N797), .Y(n3384) );
  MX2X1 U2332 ( .A(SHA256_result[62]), .B(SHA256_result[94]), .S0(n2871), .Y(
        n365) );
  OAI2BB1X1 U2333 ( .A0N(SHA256_result[190]), .A1N(n2855), .B0(n3202), .Y(
        f2_ABC_32[30]) );
  OAI21XL U2334 ( .A0(n2855), .A1(SHA256_result[190]), .B0(SHA256_result[222]), 
        .Y(n3202) );
  OAI2BB1X1 U2335 ( .A0N(SHA256_result[189]), .A1N(SHA256_result[221]), .B0(
        n3203), .Y(f2_ABC_32[29]) );
  OAI21XL U2336 ( .A0(SHA256_result[221]), .A1(SHA256_result[189]), .B0(n2849), 
        .Y(n3203) );
  OAI2BB1X1 U2337 ( .A0N(SHA256_result[251]), .A1N(SHA256_result[219]), .B0(
        n3205), .Y(f2_ABC_32[27]) );
  OAI21XL U2338 ( .A0(SHA256_result[251]), .A1(SHA256_result[219]), .B0(
        SHA256_result[187]), .Y(n3205) );
  OAI2BB1X1 U2339 ( .A0N(n2862), .A1N(SHA256_result[220]), .B0(n3204), .Y(
        f2_ABC_32[28]) );
  OAI21XL U2340 ( .A0(n2862), .A1(SHA256_result[220]), .B0(SHA256_result[188]), 
        .Y(n3204) );
  INVX1 U2341 ( .A(read_counter[0]), .Y(n3724) );
  XOR3X2 U2342 ( .A(SHA256_result[236]), .B(n2906), .C(n2891), .Y(f3_A_32[31])
         );
  OAI2BB1X1 U2343 ( .A0N(SHA256_result[191]), .A1N(n2887), .B0(n3201), .Y(
        f2_ABC_32[31]) );
  OAI21XL U2344 ( .A0(SHA256_result[191]), .A1(n2887), .B0(SHA256_result[223]), 
        .Y(n3201) );
  INVX1 U2345 ( .A(read_counter[1]), .Y(n3725) );
  NOR2X1 U2346 ( .A(n3724), .B(read_counter[1]), .Y(n1081) );
  INVXL U2347 ( .A(n1168), .Y(n3837) );
  INVX1 U2348 ( .A(N957), .Y(n3312) );
  INVX1 U2349 ( .A(N988), .Y(n3179) );
  INVXL U2350 ( .A(n1167), .Y(n3722) );
  INVXL U2351 ( .A(SHA256_result[166]), .Y(n3859) );
  INVXL U2352 ( .A(SHA256_result[169]), .Y(n3544) );
  INVX1 U2353 ( .A(SHA256_result[223]), .Y(n3843) );
  INVXL U2354 ( .A(SHA256_result[199]), .Y(n3825) );
  INVX1 U2355 ( .A(SHA256_result[95]), .Y(n3857) );
  INVXL U2356 ( .A(SHA256_result[160]), .Y(n3490) );
  INVX1 U2357 ( .A(N987), .Y(n3190) );
  INVX1 U2358 ( .A(N827), .Y(n3521) );
  NAND2BXL U2359 ( .AN(n3057), .B(n2934), .Y(n3328) );
  AOI21XL U2360 ( .A0(n3012), .A1(n2934), .B0(n3123), .Y(n844) );
  AOI2BB2XL U2361 ( .B0(n2934), .B1(n2988), .A0N(n3039), .A1N(n3525), .Y(n3526) );
  AOI22XL U2362 ( .A0(n3107), .A1(n3837), .B0(n3104), .B1(n2934), .Y(n1236) );
  XOR3X2 U2363 ( .A(n2934), .B(SHA256_result[114]), .C(n2873), .Y(f4_E_32[7])
         );
  XOR3X2 U2364 ( .A(n2934), .B(n2878), .C(n2864), .Y(f4_E_32[21]) );
  XOR3X2 U2365 ( .A(n2934), .B(n2884), .C(n2840), .Y(f4_E_32[26]) );
  NAND2XL U2366 ( .A(next_A[30]), .B(n3036), .Y(n3294) );
  NAND2XL U2367 ( .A(n3037), .B(next_A[25]), .Y(n3300) );
  NAND2XL U2368 ( .A(next_E[20]), .B(n3035), .Y(n3388) );
  NAND2BXL U2369 ( .AN(n3057), .B(n2383), .Y(n3464) );
  AOI21XL U2370 ( .A0(n2827), .A1(n3004), .B0(n3118), .Y(n899) );
  NAND2XL U2371 ( .A(n2827), .B(n2986), .Y(n3191) );
  AOI22XL U2372 ( .A0(N1019), .A1(n2936), .B0(n2827), .B1(n3028), .Y(n934) );
  AOI22XL U2373 ( .A0(n3103), .A1(SHA256_result[0]), .B0(n3100), .B1(n2827), 
        .Y(n1235) );
  NAND2XL U2374 ( .A(next_E[22]), .B(n3035), .Y(n3446) );
  CLKINVX3 U2375 ( .A(n3168), .Y(n3167) );
  CLKINVX4 U2376 ( .A(SHA256_result[44]), .Y(n3819) );
  CLKINVX4 U2377 ( .A(SHA256_result[66]), .Y(n3182) );
  CLKINVX4 U2378 ( .A(SHA256_result[41]), .Y(n3422) );
  CLKINVX4 U2379 ( .A(SHA256_result[73]), .Y(n3425) );
  MXI2X4 U2380 ( .A(n3422), .B(n3425), .S0(n2869), .Y(n321) );
  CLKINVX4 U2381 ( .A(SHA256_result[39]), .Y(n3302) );
  MXI2X4 U2382 ( .A(n3302), .B(n1161), .S0(n2830), .Y(f1_EFG_32[7]) );
  CLKINVX4 U2383 ( .A(SHA256_result[38]), .Y(n3321) );
  CLKINVX4 U2384 ( .A(SHA256_result[70]), .Y(n3254) );
  MXI2X4 U2385 ( .A(n3321), .B(n3254), .S0(n2833), .Y(n353) );
  CLKINVX4 U2386 ( .A(SHA256_result[37]), .Y(n3318) );
  MXI2X4 U2387 ( .A(n3318), .B(n1163), .S0(n2840), .Y(f1_EFG_32[5]) );
  CLKINVX4 U2388 ( .A(SHA256_result[34]), .Y(n3324) );
  MXI2X4 U2389 ( .A(n3324), .B(n3182), .S0(n2844), .Y(f1_EFG_32[2]) );
  MXI2X4 U2390 ( .A(n3315), .B(n1167), .S0(n2851), .Y(f1_EFG_32[1]) );
  XOR3X4 U2391 ( .A(SHA256_result[102]), .B(SHA256_result[121]), .C(n2858), 
        .Y(f4_E_32[0]) );
  OAI2BB1X4 U2392 ( .A0N(SHA256_result[235]), .A1N(SHA256_result[171]), .B0(
        n3221), .Y(f2_ABC_32[11]) );
  OAI2BB1X4 U2393 ( .A0N(SHA256_result[170]), .A1N(SHA256_result[234]), .B0(
        n3222), .Y(f2_ABC_32[10]) );
  OAI21X4 U2394 ( .A0(n2923), .A1(SHA256_result[167]), .B0(SHA256_result[199]), 
        .Y(n3225) );
  OAI2BB1X4 U2395 ( .A0N(n2923), .A1N(SHA256_result[167]), .B0(n3225), .Y(
        f2_ABC_32[7]) );
  OAI21X4 U2396 ( .A0(SHA256_result[198]), .A1(n2924), .B0(SHA256_result[166]), 
        .Y(n3226) );
  OAI2BB1X4 U2397 ( .A0N(SHA256_result[198]), .A1N(n2924), .B0(n3226), .Y(
        f2_ABC_32[6]) );
  OAI21X4 U2398 ( .A0(SHA256_result[165]), .A1(n2928), .B0(SHA256_result[197]), 
        .Y(n3227) );
  OAI2BB1X4 U2399 ( .A0N(SHA256_result[165]), .A1N(n2928), .B0(n3227), .Y(
        f2_ABC_32[5]) );
  OAI2BB1X4 U2400 ( .A0N(SHA256_result[163]), .A1N(SHA256_result[195]), .B0(
        n3229), .Y(f2_ABC_32[3]) );
  OAI21X4 U2401 ( .A0(n2933), .A1(SHA256_result[192]), .B0(SHA256_result[160]), 
        .Y(n3232) );
  OAI2BB1X4 U2402 ( .A0N(n2933), .A1N(SHA256_result[192]), .B0(n3232), .Y(
        f2_ABC_32[0]) );
  NAND2X4 U2403 ( .A(N826), .B(n2946), .Y(n3376) );
endmodule


module controller_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module controller ( clk, reset, first_block, last_block, output_enable, busy, 
        inner_busy );
  input clk, reset, first_block, last_block;
  output output_enable, busy, inner_busy;
  wire   N11, N24, N25, N26, N27, N28, N29, N30, N47, N48, N49, n12, n19, n5,
         n6, n7, n18, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n40,
         n41, n42, n43;
  wire   [1:0] state;
  wire   [6:0] counter1;
  wire   [2:0] counter2;

  CLKINVX8 U24 ( .A(reset), .Y(n12) );
  CLKINVX4 U26 ( .A(reset), .Y(n18) );
  controller_DW01_inc_0 add_82 ( .A(counter1), .SUM({N30, N29, N28, N27, N26, 
        N25, N24}) );
  DFFHQX1 counter2_reg_2_ ( .D(N49), .CK(clk), .Q(counter2[2]) );
  DFFHQX1 counter2_reg_0_ ( .D(N47), .CK(clk), .Q(counter2[0]) );
  DFFHQX1 counter2_reg_1_ ( .D(N48), .CK(clk), .Q(counter2[1]) );
  DFFTRX1 counter1_reg_1_ ( .D(N25), .RN(n19), .CK(clk), .Q(counter1[1]) );
  DFFTRX1 counter1_reg_3_ ( .D(N27), .RN(n19), .CK(clk), .Q(counter1[3]) );
  DFFTRX1 counter1_reg_2_ ( .D(N26), .RN(n19), .CK(clk), .Q(counter1[2]) );
  DFFTRX1 counter1_reg_6_ ( .D(N30), .RN(n19), .CK(clk), .Q(counter1[6]) );
  DFFTRX1 state_reg_0_ ( .D(n12), .RN(n41), .CK(clk), .Q(state[0]) );
  DFFHQX1 state_reg_1_ ( .D(N11), .CK(clk), .Q(state[1]) );
  DFFTRXL counter1_reg_5_ ( .D(N29), .RN(n19), .CK(clk), .Q(counter1[5]), .QN(
        n6) );
  DFFTRXL counter1_reg_4_ ( .D(N28), .RN(n19), .CK(clk), .Q(counter1[4]), .QN(
        n5) );
  DFFTRXL counter1_reg_0_ ( .D(N24), .RN(n19), .CK(clk), .Q(counter1[0]), .QN(
        n7) );
  AOI22XL U3 ( .A0(n22), .A1(inner_busy), .B0(first_block), .B1(n23), .Y(n21)
         );
  INVX1 U4 ( .A(n23), .Y(busy) );
  INVX1 U5 ( .A(n22), .Y(n40) );
  NOR2BX2 U6 ( .AN(state[1]), .B(state[0]), .Y(output_enable) );
  NOR2X1 U7 ( .A(state[1]), .B(state[0]), .Y(n23) );
  AOI211X1 U8 ( .A0(n24), .A1(n43), .B0(reset), .C0(n40), .Y(n19) );
  INVX1 U9 ( .A(last_block), .Y(n43) );
  INVX1 U10 ( .A(n21), .Y(n41) );
  NOR2BX1 U11 ( .AN(state[0]), .B(state[1]), .Y(inner_busy) );
  NAND2X1 U12 ( .A(output_enable), .B(n18), .Y(n27) );
  OAI211X1 U13 ( .A0(counter2[2]), .A1(n27), .B0(n29), .C0(n25), .Y(N11) );
  NAND3X1 U14 ( .A(inner_busy), .B(n18), .C(n40), .Y(n29) );
  AOI2BB1X1 U15 ( .A0N(counter2[1]), .A1N(n27), .B0(N47), .Y(n25) );
  NOR2X1 U16 ( .A(n27), .B(counter2[0]), .Y(N47) );
  OAI21XL U17 ( .A0(n25), .A1(n42), .B0(n26), .Y(N49) );
  NAND4BXL U18 ( .AN(n27), .B(counter2[1]), .C(counter2[0]), .D(n42), .Y(n26)
         );
  INVX1 U19 ( .A(counter2[2]), .Y(n42) );
  NOR2X1 U20 ( .A(n28), .B(n27), .Y(N48) );
  XNOR2X1 U21 ( .A(counter2[0]), .B(counter2[1]), .Y(n28) );
  NAND2X1 U22 ( .A(n24), .B(counter1[6]), .Y(n22) );
  AND4X2 U23 ( .A(n6), .B(n5), .C(n7), .D(n30), .Y(n24) );
  NOR3X1 U25 ( .A(counter1[2]), .B(counter1[3]), .C(counter1[1]), .Y(n30) );
endmodule


module top ( clk, reset, data, write_enable, last_block, first_block, busy, 
        digest, output_enable );
  input [31:0] data;
  output [31:0] digest;
  input clk, reset, write_enable, last_block, first_block;
  output busy, output_enable;
  wire   inner_busy;
  wire   [31:0] Wt;

  message_schedule our_message_schedule ( .clk(clk), .reset(reset), .data(data), .write_enable(write_enable), .inner_busy(inner_busy), .Wt(Wt) );
  hash_core our_hash_core ( .clk(clk), .reset(reset), .Wt(Wt), .inner_busy(
        inner_busy), .first_block(first_block), .output_enable(output_enable), 
        .digest(digest) );
  controller our_controller ( .clk(clk), .reset(reset), .first_block(
        first_block), .last_block(last_block), .output_enable(output_enable), 
        .busy(busy), .inner_busy(inner_busy) );
endmodule


module sha256_chip ( clk, reset, data, write_enable, last_block, first_block, 
        busy, digest, output_enable );
  input [31:0] data;
  output [31:0] digest;
  input clk, reset, write_enable, last_block, first_block;
  output busy, output_enable;
  wire   net_clk, net_reset, net_write_enable, net_last_block, net_first_block,
         net_busy, net_output_enable;
  wire   [31:0] net_data;
  wire   [31:0] net_digest;

  PIW PIW_clk ( .PAD(clk), .C(net_clk) );
  PIW PIW_reset ( .PAD(reset), .C(net_reset) );
  PIW PIW_data0 ( .PAD(data[0]), .C(net_data[0]) );
  PIW PIW_data1 ( .PAD(data[1]), .C(net_data[1]) );
  PIW PIW_data2 ( .PAD(data[2]), .C(net_data[2]) );
  PIW PIW_data3 ( .PAD(data[3]), .C(net_data[3]) );
  PIW PIW_data4 ( .PAD(data[4]), .C(net_data[4]) );
  PIW PIW_data5 ( .PAD(data[5]), .C(net_data[5]) );
  PIW PIW_data6 ( .PAD(data[6]), .C(net_data[6]) );
  PIW PIW_data7 ( .PAD(data[7]), .C(net_data[7]) );
  PIW PIW_data8 ( .PAD(data[8]), .C(net_data[8]) );
  PIW PIW_data9 ( .PAD(data[9]), .C(net_data[9]) );
  PIW PIW_data10 ( .PAD(data[10]), .C(net_data[10]) );
  PIW PIW_data11 ( .PAD(data[11]), .C(net_data[11]) );
  PIW PIW_data12 ( .PAD(data[12]), .C(net_data[12]) );
  PIW PIW_data13 ( .PAD(data[13]), .C(net_data[13]) );
  PIW PIW_data14 ( .PAD(data[14]), .C(net_data[14]) );
  PIW PIW_data15 ( .PAD(data[15]), .C(net_data[15]) );
  PIW PIW_data16 ( .PAD(data[16]), .C(net_data[16]) );
  PIW PIW_data17 ( .PAD(data[17]), .C(net_data[17]) );
  PIW PIW_data18 ( .PAD(data[18]), .C(net_data[18]) );
  PIW PIW_data19 ( .PAD(data[19]), .C(net_data[19]) );
  PIW PIW_data20 ( .PAD(data[20]), .C(net_data[20]) );
  PIW PIW_data21 ( .PAD(data[21]), .C(net_data[21]) );
  PIW PIW_data22 ( .PAD(data[22]), .C(net_data[22]) );
  PIW PIW_data23 ( .PAD(data[23]), .C(net_data[23]) );
  PIW PIW_data24 ( .PAD(data[24]), .C(net_data[24]) );
  PIW PIW_data25 ( .PAD(data[25]), .C(net_data[25]) );
  PIW PIW_data26 ( .PAD(data[26]), .C(net_data[26]) );
  PIW PIW_data27 ( .PAD(data[27]), .C(net_data[27]) );
  PIW PIW_data28 ( .PAD(data[28]), .C(net_data[28]) );
  PIW PIW_data29 ( .PAD(data[29]), .C(net_data[29]) );
  PIW PIW_data30 ( .PAD(data[30]), .C(net_data[30]) );
  PIW PIW_data31 ( .PAD(data[31]), .C(net_data[31]) );
  PIW PIW_write_enable ( .PAD(write_enable), .C(net_write_enable) );
  PIW PIW_last_block ( .PAD(last_block), .C(net_last_block) );
  PIW PIW_first_block ( .PAD(first_block), .C(net_first_block) );
  PO8W PO8W_busy ( .I(net_busy), .PAD(busy) );
  PO8W PO8W_digest0 ( .I(net_digest[0]), .PAD(digest[0]) );
  PO8W PO8W_digest1 ( .I(net_digest[1]), .PAD(digest[1]) );
  PO8W PO8W_digest2 ( .I(net_digest[2]), .PAD(digest[2]) );
  PO8W PO8W_digest3 ( .I(net_digest[3]), .PAD(digest[3]) );
  PO8W PO8W_digest4 ( .I(net_digest[4]), .PAD(digest[4]) );
  PO8W PO8W_digest5 ( .I(net_digest[5]), .PAD(digest[5]) );
  PO8W PO8W_digest6 ( .I(net_digest[6]), .PAD(digest[6]) );
  PO8W PO8W_digest7 ( .I(net_digest[7]), .PAD(digest[7]) );
  PO8W PO8W_digest8 ( .I(net_digest[8]), .PAD(digest[8]) );
  PO8W PO8W_digest9 ( .I(net_digest[9]), .PAD(digest[9]) );
  PO8W PO8W_digest10 ( .I(net_digest[10]), .PAD(digest[10]) );
  PO8W PO8W_digest11 ( .I(net_digest[11]), .PAD(digest[11]) );
  PO8W PO8W_digest12 ( .I(net_digest[12]), .PAD(digest[12]) );
  PO8W PO8W_digest13 ( .I(net_digest[13]), .PAD(digest[13]) );
  PO8W PO8W_digest14 ( .I(net_digest[14]), .PAD(digest[14]) );
  PO8W PO8W_digest15 ( .I(net_digest[15]), .PAD(digest[15]) );
  PO8W PO8W_digest16 ( .I(net_digest[16]), .PAD(digest[16]) );
  PO8W PO8W_digest17 ( .I(net_digest[17]), .PAD(digest[17]) );
  PO8W PO8W_digest18 ( .I(net_digest[18]), .PAD(digest[18]) );
  PO8W PO8W_digest19 ( .I(net_digest[19]), .PAD(digest[19]) );
  PO8W PO8W_digest20 ( .I(net_digest[20]), .PAD(digest[20]) );
  PO8W PO8W_digest21 ( .I(net_digest[21]), .PAD(digest[21]) );
  PO8W PO8W_digest22 ( .I(net_digest[22]), .PAD(digest[22]) );
  PO8W PO8W_digest23 ( .I(net_digest[23]), .PAD(digest[23]) );
  PO8W PO8W_digest24 ( .I(net_digest[24]), .PAD(digest[24]) );
  PO8W PO8W_digest25 ( .I(net_digest[25]), .PAD(digest[25]) );
  PO8W PO8W_digest26 ( .I(net_digest[26]), .PAD(digest[26]) );
  PO8W PO8W_digest27 ( .I(net_digest[27]), .PAD(digest[27]) );
  PO8W PO8W_digest28 ( .I(net_digest[28]), .PAD(digest[28]) );
  PO8W PO8W_digest29 ( .I(net_digest[29]), .PAD(digest[29]) );
  PO8W PO8W_digest30 ( .I(net_digest[30]), .PAD(digest[30]) );
  PO8W PO8W_digest31 ( .I(net_digest[31]), .PAD(digest[31]) );
  PO8W PO8W_output_enable ( .I(net_output_enable), .PAD(output_enable) );
  top inst_top ( .clk(net_clk), .reset(net_reset), .data(net_data), 
        .write_enable(net_write_enable), .last_block(net_last_block), 
        .first_block(net_first_block), .busy(net_busy), .digest(net_digest), 
        .output_enable(net_output_enable) );
endmodule



module message_schedule_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module message_schedule_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module message_schedule_DW01_add_17 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1;
  wire   [31:1] carry;

  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX4 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX4 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX4 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX4 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX4 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX4 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX4 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX4 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX4 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX4 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX4 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX4 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  INVX2 U1 ( .A(n1), .Y(carry[1]) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X4 U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module message_schedule_DW01_add_20 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215;

  OR2X4 U2 ( .A(A[3]), .B(B[3]), .Y(n212) );
  OR2X2 U3 ( .A(n11), .B(n181), .Y(n1) );
  NAND2X1 U4 ( .A(n1), .B(n157), .Y(n179) );
  CLKINVX3 U5 ( .A(n182), .Y(n181) );
  OAI21X4 U6 ( .A0(n184), .A1(n161), .B0(n162), .Y(n182) );
  NOR2X1 U7 ( .A(A[9]), .B(B[9]), .Y(n8) );
  NAND2X1 U8 ( .A(n94), .B(n95), .Y(n74) );
  OAI21X2 U9 ( .A0(n160), .A1(n7), .B0(n149), .Y(n145) );
  INVX1 U10 ( .A(n150), .Y(n149) );
  NAND2X1 U11 ( .A(n115), .B(n110), .Y(n113) );
  OR2X2 U12 ( .A(A[5]), .B(B[5]), .Y(n36) );
  NAND2X1 U13 ( .A(B[4]), .B(A[4]), .Y(n39) );
  INVX1 U14 ( .A(n159), .Y(n202) );
  INVX1 U15 ( .A(n189), .Y(n194) );
  INVX1 U16 ( .A(n18), .Y(n201) );
  OAI21XL U17 ( .A0(n178), .A1(n12), .B0(n158), .Y(n176) );
  INVX1 U18 ( .A(n179), .Y(n178) );
  NOR2X2 U19 ( .A(n49), .B(n51), .Y(n210) );
  NAND2X4 U20 ( .A(n145), .B(n146), .Y(n122) );
  OAI21X4 U21 ( .A0(n9), .A1(n184), .B0(n23), .Y(n18) );
  INVX4 U22 ( .A(n21), .Y(n184) );
  NOR2XL U23 ( .A(n40), .B(n45), .Y(n214) );
  NAND2XL U24 ( .A(B[9]), .B(A[9]), .Y(n20) );
  OR2X1 U25 ( .A(A[4]), .B(B[4]), .Y(n37) );
  NAND2X1 U26 ( .A(B[6]), .B(A[6]), .Y(n30) );
  OR2X1 U27 ( .A(A[1]), .B(B[1]), .Y(n64) );
  OR2X2 U28 ( .A(A[6]), .B(B[6]), .Y(n206) );
  OAI21X2 U29 ( .A0(n204), .A1(n205), .B0(n26), .Y(n165) );
  NOR2BXL U30 ( .AN(n48), .B(n49), .Y(n47) );
  XNOR2X1 U31 ( .A(n113), .B(n4), .Y(SUM[22]) );
  NAND2X1 U32 ( .A(n106), .B(n101), .Y(n4) );
  XNOR2X1 U33 ( .A(n56), .B(n2), .Y(SUM[30]) );
  NAND2X1 U34 ( .A(B[1]), .B(A[1]), .Y(n65) );
  NAND2XL U35 ( .A(B[2]), .B(A[2]), .Y(n52) );
  OAI21XL U36 ( .A0(n139), .A1(n128), .B0(n127), .Y(n137) );
  OAI21XL U37 ( .A0(n50), .A1(n51), .B0(n52), .Y(n46) );
  NOR2XL U38 ( .A(n39), .B(n40), .Y(n33) );
  OAI21XL U39 ( .A0(n12), .A1(n157), .B0(n158), .Y(n154) );
  OAI21XL U40 ( .A0(n151), .A1(n13), .B0(n152), .Y(n150) );
  INVX1 U41 ( .A(n156), .Y(n155) );
  NAND2X1 U42 ( .A(n142), .B(n132), .Y(n140) );
  NOR2X1 U43 ( .A(A[13]), .B(B[13]), .Y(n12) );
  NAND2XL U44 ( .A(B[5]), .B(A[5]), .Y(n34) );
  NAND2X1 U45 ( .A(B[8]), .B(A[8]), .Y(n23) );
  OAI2BB1X2 U46 ( .A0N(n202), .A1N(n38), .B0(n203), .Y(n21) );
  OAI21X2 U47 ( .A0(n8), .A1(n201), .B0(n20), .Y(n199) );
  NAND2XL U48 ( .A(n206), .B(n207), .Y(n205) );
  NAND3BX2 U49 ( .AN(n170), .B(n48), .C(n168), .Y(n38) );
  NOR2BXL U50 ( .AN(n156), .B(n173), .Y(n177) );
  XOR2X2 U51 ( .A(n174), .B(n175), .Y(SUM[15]) );
  NOR2BXL U52 ( .AN(n152), .B(n13), .Y(n175) );
  INVXL U53 ( .A(n212), .Y(n49) );
  NAND2X1 U54 ( .A(n54), .B(n57), .Y(n2) );
  OAI21X1 U55 ( .A0(n58), .A1(n59), .B0(n60), .Y(n56) );
  NOR2BX1 U56 ( .AN(n133), .B(n125), .Y(n124) );
  XNOR2X1 U57 ( .A(n89), .B(n3), .Y(SUM[26]) );
  NAND2X1 U58 ( .A(n82), .B(n77), .Y(n3) );
  NOR2BXL U59 ( .AN(n39), .B(n45), .Y(n44) );
  NOR2BXL U60 ( .AN(n30), .B(n29), .Y(n32) );
  NOR2BXL U61 ( .AN(n132), .B(n130), .Y(n144) );
  NOR2BXL U62 ( .AN(n23), .B(n9), .Y(n22) );
  INVXL U63 ( .A(n161), .Y(n166) );
  AOI21XL U64 ( .A0(n167), .A1(n168), .B0(n159), .Y(n164) );
  NOR2XL U65 ( .A(n169), .B(n170), .Y(n167) );
  NAND3XL U66 ( .A(n36), .B(n37), .C(n38), .Y(n35) );
  NAND2X2 U67 ( .A(n118), .B(n119), .Y(n98) );
  XNOR2X1 U68 ( .A(n94), .B(n5), .Y(SUM[24]) );
  NAND2X1 U69 ( .A(n85), .B(n95), .Y(n5) );
  XOR2XL U70 ( .A(n67), .B(n59), .Y(SUM[29]) );
  XNOR2X1 U71 ( .A(n68), .B(n6), .Y(SUM[28]) );
  NAND2X1 U72 ( .A(n71), .B(n69), .Y(n6) );
  NAND2XL U73 ( .A(n52), .B(n66), .Y(n62) );
  NAND2XL U74 ( .A(n56), .B(n57), .Y(n55) );
  NAND2XL U75 ( .A(B[3]), .B(A[3]), .Y(n48) );
  NAND2XL U76 ( .A(B[7]), .B(A[7]), .Y(n26) );
  NAND2XL U77 ( .A(B[10]), .B(A[10]), .Y(n191) );
  NAND2XL U78 ( .A(B[11]), .B(A[11]), .Y(n188) );
  NOR2XL U79 ( .A(A[0]), .B(B[0]), .Y(n15) );
  AND2X1 U80 ( .A(B[0]), .B(A[0]), .Y(n16) );
  NOR2XL U81 ( .A(A[12]), .B(B[12]), .Y(n11) );
  NAND2XL U82 ( .A(B[0]), .B(A[0]), .Y(n17) );
  NAND2XL U83 ( .A(B[17]), .B(A[17]), .Y(n132) );
  NAND2XL U84 ( .A(B[13]), .B(A[13]), .Y(n158) );
  NAND2XL U85 ( .A(B[15]), .B(A[15]), .Y(n152) );
  NAND3XL U86 ( .A(A[0]), .B(B[0]), .C(n64), .Y(n63) );
  AND2X1 U87 ( .A(n65), .B(n63), .Y(n50) );
  INVX1 U88 ( .A(n165), .Y(n203) );
  NAND2X1 U89 ( .A(n214), .B(n215), .Y(n159) );
  NOR2X1 U90 ( .A(n27), .B(n29), .Y(n215) );
  AND2X2 U91 ( .A(n162), .B(n163), .Y(n7) );
  INVX1 U92 ( .A(n36), .Y(n40) );
  INVX1 U93 ( .A(n206), .Y(n29) );
  AOI21X1 U94 ( .A0(n185), .A1(n186), .B0(n187), .Y(n162) );
  INVX1 U95 ( .A(n188), .Y(n187) );
  OAI2BB1X1 U96 ( .A0N(n189), .A1N(n190), .B0(n191), .Y(n186) );
  OAI21XL U97 ( .A0(n8), .A1(n23), .B0(n20), .Y(n190) );
  NOR2X1 U98 ( .A(n208), .B(n209), .Y(n204) );
  NAND2X1 U99 ( .A(n30), .B(n34), .Y(n209) );
  INVX1 U100 ( .A(n37), .Y(n45) );
  INVX1 U101 ( .A(n66), .Y(n51) );
  INVX1 U102 ( .A(n207), .Y(n27) );
  XOR2X1 U103 ( .A(n199), .B(n200), .Y(SUM[10]) );
  NOR2BX1 U104 ( .AN(n191), .B(n194), .Y(n200) );
  XOR2X1 U105 ( .A(n179), .B(n180), .Y(SUM[13]) );
  NOR2BX1 U106 ( .AN(n158), .B(n12), .Y(n180) );
  XOR2X1 U107 ( .A(n18), .B(n19), .Y(SUM[9]) );
  NOR2BX1 U108 ( .AN(n20), .B(n8), .Y(n19) );
  XOR2X1 U109 ( .A(n176), .B(n177), .Y(SUM[14]) );
  XOR2X1 U110 ( .A(n24), .B(n25), .Y(SUM[7]) );
  NOR2BX1 U111 ( .AN(n26), .B(n27), .Y(n25) );
  OAI21XL U112 ( .A0(n28), .A1(n29), .B0(n30), .Y(n24) );
  INVX1 U113 ( .A(n31), .Y(n28) );
  XOR2X1 U114 ( .A(n196), .B(n197), .Y(SUM[11]) );
  NOR2BX1 U115 ( .AN(n188), .B(n195), .Y(n197) );
  OAI21XL U116 ( .A0(n198), .A1(n194), .B0(n191), .Y(n196) );
  INVX1 U117 ( .A(n199), .Y(n198) );
  OAI2BB1X1 U118 ( .A0N(n153), .A1N(n176), .B0(n156), .Y(n174) );
  NAND3BX1 U119 ( .AN(n33), .B(n34), .C(n35), .Y(n31) );
  NOR2X1 U120 ( .A(n40), .B(n39), .Y(n208) );
  INVX1 U121 ( .A(n213), .Y(n170) );
  NAND2BX1 U122 ( .AN(n52), .B(n212), .Y(n213) );
  AOI21X1 U123 ( .A0(n68), .A1(n69), .B0(n70), .Y(n59) );
  INVX1 U124 ( .A(n71), .Y(n70) );
  OAI21XL U125 ( .A0(n122), .A1(n123), .B0(n124), .Y(n118) );
  NAND3BX1 U126 ( .AN(n10), .B(n134), .C(n135), .Y(n123) );
  INVX1 U127 ( .A(n61), .Y(n58) );
  INVX1 U128 ( .A(n134), .Y(n128) );
  XOR2X1 U129 ( .A(n92), .B(n93), .Y(SUM[25]) );
  NOR2BX1 U130 ( .AN(n86), .B(n84), .Y(n93) );
  NAND2X1 U131 ( .A(n60), .B(n61), .Y(n67) );
  XOR2X1 U132 ( .A(n41), .B(n42), .Y(SUM[5]) );
  NAND2X1 U133 ( .A(n36), .B(n34), .Y(n41) );
  AOI21X1 U134 ( .A0(n38), .A1(n37), .B0(n43), .Y(n42) );
  INVX1 U135 ( .A(n39), .Y(n43) );
  INVX1 U136 ( .A(n135), .Y(n130) );
  INVX1 U137 ( .A(n153), .Y(n173) );
  INVX1 U138 ( .A(n185), .Y(n195) );
  XOR2X1 U139 ( .A(n46), .B(n47), .Y(SUM[3]) );
  XOR2X1 U140 ( .A(n38), .B(n44), .Y(SUM[4]) );
  AOI21X1 U141 ( .A0(n126), .A1(n127), .B0(n10), .Y(n125) );
  NAND2BX1 U142 ( .AN(n128), .B(n129), .Y(n126) );
  OAI21XL U143 ( .A0(n130), .A1(n131), .B0(n132), .Y(n129) );
  XOR2X1 U144 ( .A(n118), .B(n120), .Y(SUM[20]) );
  NOR2BX1 U145 ( .AN(n109), .B(n121), .Y(n120) );
  INVX1 U146 ( .A(n119), .Y(n121) );
  XOR2X1 U147 ( .A(n182), .B(n183), .Y(SUM[12]) );
  NOR2BX1 U148 ( .AN(n157), .B(n11), .Y(n183) );
  XOR2X1 U149 ( .A(n31), .B(n32), .Y(SUM[6]) );
  XOR2X1 U150 ( .A(n137), .B(n138), .Y(SUM[19]) );
  NOR2BX1 U151 ( .AN(n133), .B(n10), .Y(n138) );
  INVX1 U152 ( .A(n140), .Y(n139) );
  XOR2X1 U153 ( .A(n143), .B(n144), .Y(SUM[17]) );
  XOR2X1 U154 ( .A(n116), .B(n117), .Y(SUM[21]) );
  NOR2BX1 U155 ( .AN(n110), .B(n108), .Y(n117) );
  XOR2X1 U156 ( .A(n62), .B(n50), .Y(SUM[2]) );
  XOR2X1 U157 ( .A(n111), .B(n112), .Y(SUM[23]) );
  NAND2X1 U158 ( .A(n104), .B(n100), .Y(n111) );
  AOI21X1 U159 ( .A0(n101), .A1(n113), .B0(n114), .Y(n112) );
  INVX1 U160 ( .A(n106), .Y(n114) );
  XOR2X1 U161 ( .A(n87), .B(n88), .Y(SUM[27]) );
  NAND2X1 U162 ( .A(n80), .B(n76), .Y(n87) );
  AOI21X1 U163 ( .A0(n77), .A1(n89), .B0(n90), .Y(n88) );
  INVX1 U164 ( .A(n82), .Y(n90) );
  XOR2X1 U165 ( .A(n140), .B(n141), .Y(SUM[18]) );
  NOR2BX1 U166 ( .AN(n127), .B(n128), .Y(n141) );
  XOR2X1 U167 ( .A(n21), .B(n22), .Y(SUM[8]) );
  XOR2X1 U168 ( .A(n145), .B(n147), .Y(SUM[16]) );
  NOR2BX1 U169 ( .AN(n131), .B(n148), .Y(n147) );
  INVX1 U170 ( .A(n146), .Y(n148) );
  NAND2X1 U171 ( .A(n74), .B(n85), .Y(n92) );
  NAND2X1 U172 ( .A(n122), .B(n131), .Y(n143) );
  NAND2X1 U173 ( .A(n98), .B(n109), .Y(n116) );
  OAI21XL U174 ( .A0(n164), .A1(n165), .B0(n166), .Y(n163) );
  AOI21X1 U175 ( .A0(n153), .A1(n154), .B0(n155), .Y(n151) );
  NAND2X1 U176 ( .A(n99), .B(n116), .Y(n115) );
  NAND2X1 U177 ( .A(n91), .B(n86), .Y(n89) );
  NAND2X1 U178 ( .A(n75), .B(n92), .Y(n91) );
  NAND2X1 U179 ( .A(n72), .B(n73), .Y(n68) );
  AOI21X1 U180 ( .A0(n78), .A1(n76), .B0(n79), .Y(n72) );
  NAND4BXL U181 ( .AN(n74), .B(n75), .C(n76), .D(n77), .Y(n73) );
  INVX1 U182 ( .A(n80), .Y(n79) );
  NAND2X1 U183 ( .A(n96), .B(n97), .Y(n94) );
  AOI21X1 U184 ( .A0(n102), .A1(n100), .B0(n103), .Y(n96) );
  NAND4BXL U185 ( .AN(n98), .B(n99), .C(n100), .D(n101), .Y(n97) );
  INVX1 U186 ( .A(n104), .Y(n103) );
  NAND2X1 U187 ( .A(n192), .B(n193), .Y(n161) );
  NOR2X1 U188 ( .A(n194), .B(n195), .Y(n192) );
  NOR2X1 U189 ( .A(n9), .B(n8), .Y(n193) );
  INVX1 U190 ( .A(n48), .Y(n169) );
  NAND2X1 U191 ( .A(n135), .B(n143), .Y(n142) );
  NAND2X1 U192 ( .A(n54), .B(n55), .Y(n53) );
  NAND2X1 U193 ( .A(n65), .B(n64), .Y(n136) );
  NAND2X1 U194 ( .A(n171), .B(n172), .Y(n160) );
  NOR2X1 U195 ( .A(n13), .B(n173), .Y(n172) );
  NOR2X1 U196 ( .A(n12), .B(n11), .Y(n171) );
  INVX1 U197 ( .A(n99), .Y(n108) );
  NAND2X1 U198 ( .A(n105), .B(n106), .Y(n102) );
  NAND2X1 U199 ( .A(n101), .B(n107), .Y(n105) );
  OAI21XL U200 ( .A0(n108), .A1(n109), .B0(n110), .Y(n107) );
  INVX1 U201 ( .A(n75), .Y(n84) );
  NAND2X1 U202 ( .A(n81), .B(n82), .Y(n78) );
  NAND2X1 U203 ( .A(n77), .B(n83), .Y(n81) );
  OAI21XL U204 ( .A0(n84), .A1(n85), .B0(n86), .Y(n83) );
  XOR3X2 U205 ( .A(B[31]), .B(A[31]), .C(n53), .Y(SUM[31]) );
  NAND3X1 U206 ( .A(n210), .B(n64), .C(n211), .Y(n168) );
  OAI2BB1X1 U207 ( .A0N(B[0]), .A1N(A[0]), .B0(n65), .Y(n211) );
  OR2X2 U208 ( .A(A[2]), .B(B[2]), .Y(n66) );
  OR2X2 U209 ( .A(A[7]), .B(B[7]), .Y(n207) );
  NOR2X1 U210 ( .A(A[8]), .B(B[8]), .Y(n9) );
  NOR2X1 U211 ( .A(A[19]), .B(B[19]), .Y(n10) );
  NAND2X1 U212 ( .A(B[16]), .B(A[16]), .Y(n131) );
  NAND2X1 U213 ( .A(B[12]), .B(A[12]), .Y(n157) );
  NAND2X1 U214 ( .A(B[14]), .B(A[14]), .Y(n156) );
  OR2X2 U215 ( .A(A[17]), .B(B[17]), .Y(n135) );
  XOR2X1 U216 ( .A(n17), .B(n136), .Y(SUM[1]) );
  OR2X2 U217 ( .A(A[14]), .B(B[14]), .Y(n153) );
  OR2X2 U218 ( .A(A[11]), .B(B[11]), .Y(n185) );
  OR2X2 U219 ( .A(A[18]), .B(B[18]), .Y(n134) );
  OR2X2 U220 ( .A(A[10]), .B(B[10]), .Y(n189) );
  NOR2X1 U221 ( .A(A[15]), .B(B[15]), .Y(n13) );
  OR2X2 U222 ( .A(A[22]), .B(B[22]), .Y(n101) );
  NAND2X1 U223 ( .A(B[20]), .B(A[20]), .Y(n109) );
  NAND2X1 U224 ( .A(B[18]), .B(A[18]), .Y(n127) );
  NAND2X1 U225 ( .A(B[22]), .B(A[22]), .Y(n106) );
  OR2X2 U226 ( .A(A[23]), .B(B[23]), .Y(n100) );
  NAND2X1 U227 ( .A(B[21]), .B(A[21]), .Y(n110) );
  OR2X2 U228 ( .A(A[21]), .B(B[21]), .Y(n99) );
  NOR2X1 U229 ( .A(n15), .B(n16), .Y(SUM[0]) );
  NAND2X1 U230 ( .A(B[23]), .B(A[23]), .Y(n104) );
  NAND2X1 U231 ( .A(B[19]), .B(A[19]), .Y(n133) );
  OR2X2 U232 ( .A(A[16]), .B(B[16]), .Y(n146) );
  OR2X2 U233 ( .A(A[20]), .B(B[20]), .Y(n119) );
  OR2X2 U234 ( .A(A[26]), .B(B[26]), .Y(n77) );
  NAND2X1 U235 ( .A(B[24]), .B(A[24]), .Y(n85) );
  NAND2X1 U236 ( .A(B[26]), .B(A[26]), .Y(n82) );
  OR2X2 U237 ( .A(A[27]), .B(B[27]), .Y(n76) );
  NAND2X1 U238 ( .A(B[25]), .B(A[25]), .Y(n86) );
  OR2X2 U239 ( .A(A[25]), .B(B[25]), .Y(n75) );
  NAND2X1 U240 ( .A(B[27]), .B(A[27]), .Y(n80) );
  OR2X2 U241 ( .A(A[24]), .B(B[24]), .Y(n95) );
  NAND2X1 U242 ( .A(B[30]), .B(A[30]), .Y(n54) );
  NAND2X1 U243 ( .A(B[29]), .B(A[29]), .Y(n60) );
  NAND2X1 U244 ( .A(B[28]), .B(A[28]), .Y(n71) );
  OR2X2 U245 ( .A(A[28]), .B(B[28]), .Y(n69) );
  OR2X2 U246 ( .A(A[30]), .B(B[30]), .Y(n57) );
  OR2X2 U247 ( .A(A[29]), .B(B[29]), .Y(n61) );
endmodule


module message_schedule_DW01_add_21 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215;

  INVX2 U2 ( .A(n170), .Y(n206) );
  NOR2BX4 U3 ( .AN(n83), .B(n77), .Y(n85) );
  OAI21X2 U4 ( .A0(n82), .A1(n77), .B0(n83), .Y(n80) );
  INVX12 U5 ( .A(n78), .Y(n77) );
  OAI21X4 U6 ( .A0(n44), .A1(n45), .B0(n46), .Y(n43) );
  OR2X4 U7 ( .A(A[27]), .B(B[27]), .Y(n79) );
  NAND2X2 U8 ( .A(n47), .B(n50), .Y(n60) );
  NOR2X4 U9 ( .A(n76), .B(n77), .Y(n68) );
  INVX4 U10 ( .A(n79), .Y(n76) );
  INVX1 U11 ( .A(n181), .Y(n180) );
  OAI21XL U12 ( .A0(n167), .A1(n163), .B0(n168), .Y(n166) );
  OR2X2 U13 ( .A(A[26]), .B(B[26]), .Y(n78) );
  NAND2X1 U14 ( .A(B[27]), .B(A[27]), .Y(n71) );
  OR2X2 U15 ( .A(A[29]), .B(B[29]), .Y(n47) );
  INVX1 U16 ( .A(n202), .Y(n195) );
  OAI2BB1X2 U17 ( .A0N(n187), .A1N(n12), .B0(n168), .Y(n185) );
  NAND2X2 U18 ( .A(n122), .B(n123), .Y(n118) );
  INVX1 U19 ( .A(n178), .Y(n177) );
  AOI21X4 U20 ( .A0(n68), .A1(n69), .B0(n70), .Y(n67) );
  INVX4 U21 ( .A(n54), .Y(n52) );
  NAND3BX1 U22 ( .AN(n72), .B(n78), .C(n79), .Y(n66) );
  AOI21X4 U23 ( .A0(n47), .A1(n42), .B0(n49), .Y(n48) );
  AOI21X4 U24 ( .A0(n41), .A1(n42), .B0(n43), .Y(n40) );
  XOR2X2 U25 ( .A(n60), .B(n61), .Y(SUM[29]) );
  NAND2X2 U26 ( .A(B[28]), .B(A[28]), .Y(n53) );
  XNOR2X2 U27 ( .A(B[31]), .B(A[31]), .Y(n39) );
  XOR2X1 U28 ( .A(B[30]), .B(A[30]), .Y(n1) );
  AOI21X2 U29 ( .A0(n54), .A1(n62), .B0(n63), .Y(n61) );
  XOR2X4 U30 ( .A(n39), .B(n40), .Y(SUM[31]) );
  XNOR2X2 U31 ( .A(n1), .B(n48), .Y(SUM[30]) );
  NAND2X2 U32 ( .A(B[30]), .B(A[30]), .Y(n46) );
  NOR2X2 U33 ( .A(A[30]), .B(B[30]), .Y(n44) );
  NAND2X4 U34 ( .A(n87), .B(n88), .Y(n86) );
  NAND2X4 U35 ( .A(n118), .B(n119), .Y(n95) );
  NAND2X4 U36 ( .A(n65), .B(n90), .Y(n88) );
  OAI21X4 U37 ( .A0(n51), .A1(n52), .B0(n53), .Y(n42) );
  NOR2BX2 U38 ( .AN(n47), .B(n2), .Y(n41) );
  NOR2X2 U39 ( .A(A[30]), .B(B[30]), .Y(n2) );
  NAND2X4 U40 ( .A(n91), .B(n92), .Y(n65) );
  OAI21X4 U41 ( .A0(n95), .A1(n96), .B0(n97), .Y(n91) );
  OAI21X4 U42 ( .A0(n65), .A1(n66), .B0(n67), .Y(n54) );
  NOR2BXL U43 ( .AN(n74), .B(n72), .Y(n89) );
  OAI21X1 U44 ( .A0(n189), .A1(n190), .B0(n191), .Y(n188) );
  INVX2 U45 ( .A(n84), .Y(n82) );
  NAND2X1 U46 ( .A(n86), .B(n74), .Y(n84) );
  INVX1 U47 ( .A(n53), .Y(n63) );
  OAI21XL U48 ( .A0(n180), .A1(n4), .B0(n159), .Y(n178) );
  OR2X2 U49 ( .A(A[10]), .B(B[10]), .Y(n197) );
  NAND2X1 U50 ( .A(B[13]), .B(A[13]), .Y(n159) );
  NAND2X1 U51 ( .A(B[14]), .B(A[14]), .Y(n160) );
  NAND2X1 U52 ( .A(B[9]), .B(A[9]), .Y(n11) );
  NOR2X1 U53 ( .A(A[13]), .B(B[13]), .Y(n4) );
  NAND2X2 U54 ( .A(n152), .B(n153), .Y(n125) );
  INVXL U55 ( .A(n169), .Y(n211) );
  NAND3BXL U56 ( .AN(n102), .B(n108), .C(n109), .Y(n96) );
  INVX2 U57 ( .A(n173), .Y(n162) );
  NAND4BBXL U58 ( .AN(n15), .BN(n5), .C(n197), .D(n192), .Y(n163) );
  NAND4BBXL U59 ( .AN(n6), .BN(n7), .C(n25), .D(n208), .Y(n171) );
  NAND2XL U60 ( .A(n95), .B(n103), .Y(n116) );
  NOR2BXL U61 ( .AN(n101), .B(n106), .Y(n111) );
  NOR2BXL U62 ( .AN(n105), .B(n107), .Y(n114) );
  NOR2BXL U63 ( .AN(n157), .B(n161), .Y(n176) );
  INVX2 U64 ( .A(n71), .Y(n70) );
  NAND2XL U65 ( .A(n205), .B(n14), .Y(n9) );
  NAND2XL U66 ( .A(n12), .B(n198), .Y(n205) );
  INVXL U67 ( .A(n92), .Y(n94) );
  INVXL U68 ( .A(n119), .Y(n121) );
  NOR2BXL U69 ( .AN(n104), .B(n102), .Y(n117) );
  NOR2BXL U70 ( .AN(n133), .B(n3), .Y(n142) );
  NOR2BXL U71 ( .AN(n202), .B(n196), .Y(n203) );
  NOR2BXL U72 ( .AN(n160), .B(n162), .Y(n179) );
  NOR2BXL U73 ( .AN(n137), .B(n127), .Y(n145) );
  NOR2BXL U74 ( .AN(n136), .B(n134), .Y(n148) );
  NAND2XL U75 ( .A(n191), .B(n192), .Y(n199) );
  AOI21XL U76 ( .A0(n197), .A1(n201), .B0(n195), .Y(n200) );
  NAND2XL U77 ( .A(n125), .B(n128), .Y(n149) );
  NAND2XL U78 ( .A(n128), .B(n129), .Y(n124) );
  INVXL U79 ( .A(n172), .Y(n183) );
  NOR2BXL U80 ( .AN(n18), .B(n19), .Y(n17) );
  NOR2BXL U81 ( .AN(n11), .B(n5), .Y(n10) );
  NOR2BXL U82 ( .AN(n27), .B(n6), .Y(n29) );
  INVXL U83 ( .A(n25), .Y(n21) );
  NOR2BXL U84 ( .AN(n34), .B(n8), .Y(n33) );
  NOR2BXL U85 ( .AN(n59), .B(n139), .Y(n138) );
  NAND2XL U86 ( .A(B[11]), .B(A[11]), .Y(n191) );
  NAND2XL U87 ( .A(B[15]), .B(A[15]), .Y(n157) );
  NAND2XL U88 ( .A(B[22]), .B(A[22]), .Y(n105) );
  NAND2XL U89 ( .A(B[19]), .B(A[19]), .Y(n133) );
  NAND2XL U90 ( .A(B[23]), .B(A[23]), .Y(n101) );
  NAND2XL U91 ( .A(B[7]), .B(A[7]), .Y(n18) );
  NAND2XL U92 ( .A(B[3]), .B(A[3]), .Y(n34) );
  OR2XL U93 ( .A(A[2]), .B(B[2]), .Y(n56) );
  NOR2X1 U94 ( .A(n106), .B(n107), .Y(n98) );
  NAND2BX1 U95 ( .AN(n165), .B(n166), .Y(n152) );
  AOI21X1 U96 ( .A0(n154), .A1(n155), .B0(n156), .Y(n153) );
  NOR2X1 U97 ( .A(n161), .B(n162), .Y(n154) );
  AOI21X1 U98 ( .A0(n164), .A1(n169), .B0(n170), .Y(n167) );
  INVX1 U99 ( .A(n171), .Y(n164) );
  OAI21XL U100 ( .A0(n211), .A1(n171), .B0(n206), .Y(n12) );
  INVX1 U101 ( .A(n163), .Y(n187) );
  OAI211X1 U102 ( .A0(n72), .A1(n73), .B0(n74), .C0(n75), .Y(n69) );
  OAI211X1 U103 ( .A0(n102), .A1(n103), .B0(n104), .C0(n105), .Y(n99) );
  INVX1 U104 ( .A(n108), .Y(n107) );
  AOI21X1 U105 ( .A0(n98), .A1(n99), .B0(n100), .Y(n97) );
  INVX1 U106 ( .A(n101), .Y(n100) );
  INVX1 U107 ( .A(n115), .Y(n102) );
  INVX1 U108 ( .A(n109), .Y(n106) );
  AOI21X1 U109 ( .A0(n130), .A1(n131), .B0(n132), .Y(n122) );
  NAND3BX1 U110 ( .AN(n124), .B(n125), .C(n126), .Y(n123) );
  INVX1 U111 ( .A(n133), .Y(n132) );
  NOR2X1 U112 ( .A(n127), .B(n3), .Y(n126) );
  XOR2X1 U113 ( .A(n54), .B(n64), .Y(SUM[28]) );
  NOR2BX1 U114 ( .AN(n53), .B(n51), .Y(n64) );
  XOR2X1 U115 ( .A(n84), .B(n85), .Y(SUM[26]) );
  XOR2X1 U116 ( .A(n88), .B(n89), .Y(SUM[25]) );
  XOR2X1 U117 ( .A(n80), .B(n81), .Y(SUM[27]) );
  NOR2BXL U118 ( .AN(n71), .B(n76), .Y(n81) );
  OAI211X1 U119 ( .A0(n4), .A1(n158), .B0(n159), .C0(n160), .Y(n155) );
  OAI211X1 U120 ( .A0(n134), .A1(n135), .B0(n136), .C0(n137), .Y(n131) );
  INVX1 U121 ( .A(n143), .Y(n127) );
  INVX1 U122 ( .A(n129), .Y(n134) );
  INVX1 U123 ( .A(n174), .Y(n161) );
  NOR2X1 U124 ( .A(n3), .B(n127), .Y(n130) );
  OAI2BB1X1 U125 ( .A0N(n115), .A1N(n116), .B0(n104), .Y(n113) );
  NAND4BXL U126 ( .AN(n4), .B(n172), .C(n173), .D(n174), .Y(n165) );
  XOR2X1 U127 ( .A(n91), .B(n93), .Y(SUM[24]) );
  NOR2BX1 U128 ( .AN(n90), .B(n94), .Y(n93) );
  XOR2X1 U129 ( .A(n113), .B(n114), .Y(SUM[22]) );
  XOR2X1 U130 ( .A(n110), .B(n111), .Y(SUM[23]) );
  OAI21XL U131 ( .A0(n112), .A1(n107), .B0(n105), .Y(n110) );
  INVX1 U132 ( .A(n113), .Y(n112) );
  OAI21XL U133 ( .A0(n207), .A1(n19), .B0(n18), .Y(n170) );
  AOI21X1 U134 ( .A0(n25), .A1(n209), .B0(n210), .Y(n207) );
  INVX1 U135 ( .A(n22), .Y(n210) );
  OAI21XL U136 ( .A0(n6), .A1(n30), .B0(n27), .Y(n209) );
  OAI21XL U137 ( .A0(n146), .A1(n134), .B0(n136), .Y(n144) );
  INVX1 U138 ( .A(n147), .Y(n146) );
  INVX1 U139 ( .A(n197), .Y(n196) );
  INVX1 U140 ( .A(n208), .Y(n19) );
  INVX1 U141 ( .A(n188), .Y(n168) );
  INVX1 U142 ( .A(n192), .Y(n190) );
  AOI21X1 U143 ( .A0(n193), .A1(n194), .B0(n195), .Y(n189) );
  NOR2X1 U144 ( .A(n5), .B(n196), .Y(n193) );
  NAND2X1 U145 ( .A(n149), .B(n135), .Y(n147) );
  NAND2X1 U146 ( .A(n14), .B(n11), .Y(n194) );
  XOR2X1 U147 ( .A(n141), .B(n142), .Y(SUM[19]) );
  OAI2BB1X1 U148 ( .A0N(n143), .A1N(n144), .B0(n137), .Y(n141) );
  XOR2X1 U149 ( .A(n116), .B(n117), .Y(SUM[21]) );
  XOR2X1 U150 ( .A(n118), .B(n120), .Y(SUM[20]) );
  NOR2BX1 U151 ( .AN(n103), .B(n121), .Y(n120) );
  INVX1 U152 ( .A(n157), .Y(n156) );
  XOR2X1 U153 ( .A(n144), .B(n145), .Y(SUM[18]) );
  XOR2X1 U154 ( .A(n147), .B(n148), .Y(SUM[17]) );
  OAI21XL U155 ( .A0(n212), .A1(n8), .B0(n34), .Y(n169) );
  AOI21X1 U156 ( .A0(n56), .A1(n213), .B0(n214), .Y(n212) );
  INVX1 U157 ( .A(n37), .Y(n214) );
  OAI21XL U158 ( .A0(n139), .A1(n140), .B0(n59), .Y(n213) );
  OAI21XL U159 ( .A0(n183), .A1(n184), .B0(n158), .Y(n181) );
  INVX1 U160 ( .A(n185), .Y(n184) );
  INVX1 U161 ( .A(n57), .Y(n139) );
  INVX1 U162 ( .A(n198), .Y(n15) );
  XOR2X1 U163 ( .A(n178), .B(n179), .Y(SUM[14]) );
  XOR2X1 U164 ( .A(n181), .B(n182), .Y(SUM[13]) );
  NOR2BX1 U165 ( .AN(n159), .B(n4), .Y(n182) );
  XOR2X1 U166 ( .A(n125), .B(n150), .Y(SUM[16]) );
  NOR2BX1 U167 ( .AN(n135), .B(n151), .Y(n150) );
  INVX1 U168 ( .A(n128), .Y(n151) );
  XOR2X1 U169 ( .A(n175), .B(n176), .Y(SUM[15]) );
  OAI21XL U170 ( .A0(n177), .A1(n162), .B0(n160), .Y(n175) );
  OAI21XL U171 ( .A0(n204), .A1(n5), .B0(n11), .Y(n201) );
  INVX1 U172 ( .A(n9), .Y(n204) );
  OAI21XL U173 ( .A0(n26), .A1(n6), .B0(n27), .Y(n23) );
  INVX1 U174 ( .A(n28), .Y(n26) );
  OAI21XL U175 ( .A0(n7), .A1(n211), .B0(n30), .Y(n28) );
  XOR2X1 U176 ( .A(n12), .B(n13), .Y(SUM[8]) );
  NOR2BX1 U177 ( .AN(n14), .B(n15), .Y(n13) );
  XOR2X1 U178 ( .A(n201), .B(n203), .Y(SUM[10]) );
  XOR2X1 U179 ( .A(n23), .B(n24), .Y(SUM[6]) );
  NOR2BX1 U180 ( .AN(n22), .B(n21), .Y(n24) );
  XOR2X1 U181 ( .A(n199), .B(n200), .Y(SUM[11]) );
  XOR2X1 U182 ( .A(n9), .B(n10), .Y(SUM[9]) );
  XOR2X1 U183 ( .A(n16), .B(n17), .Y(SUM[7]) );
  OAI21XL U184 ( .A0(n20), .A1(n21), .B0(n22), .Y(n16) );
  INVX1 U185 ( .A(n23), .Y(n20) );
  XOR2X1 U186 ( .A(n185), .B(n186), .Y(SUM[12]) );
  NOR2BX1 U187 ( .AN(n158), .B(n183), .Y(n186) );
  INVX1 U188 ( .A(n56), .Y(n36) );
  XOR2X1 U189 ( .A(n28), .B(n29), .Y(SUM[5]) );
  XOR2X1 U190 ( .A(n169), .B(n31), .Y(SUM[4]) );
  NOR2BX1 U191 ( .AN(n30), .B(n7), .Y(n31) );
  XOR2X1 U192 ( .A(n38), .B(n55), .Y(SUM[2]) );
  NOR2BX1 U193 ( .AN(n37), .B(n36), .Y(n55) );
  XOR2X1 U194 ( .A(n32), .B(n33), .Y(SUM[3]) );
  OAI21XL U195 ( .A0(n35), .A1(n36), .B0(n37), .Y(n32) );
  INVX1 U196 ( .A(n38), .Y(n35) );
  XOR2X1 U197 ( .A(n58), .B(n138), .Y(SUM[1]) );
  OAI2BB1X1 U198 ( .A0N(n57), .A1N(n58), .B0(n59), .Y(n38) );
  INVX1 U199 ( .A(n140), .Y(n58) );
  NOR2X1 U200 ( .A(A[19]), .B(B[19]), .Y(n3) );
  NAND2X1 U201 ( .A(B[25]), .B(A[25]), .Y(n74) );
  NAND2X1 U202 ( .A(A[29]), .B(B[29]), .Y(n45) );
  NAND2X1 U203 ( .A(B[29]), .B(A[29]), .Y(n50) );
  NAND2X1 U204 ( .A(B[24]), .B(A[24]), .Y(n90) );
  NAND2XL U205 ( .A(B[26]), .B(A[26]), .Y(n83) );
  NOR2X1 U206 ( .A(A[25]), .B(B[25]), .Y(n72) );
  OR2X2 U207 ( .A(A[25]), .B(B[25]), .Y(n87) );
  OR2X2 U208 ( .A(A[24]), .B(B[24]), .Y(n92) );
  OR2X2 U209 ( .A(A[23]), .B(B[23]), .Y(n109) );
  OR2X2 U210 ( .A(A[22]), .B(B[22]), .Y(n108) );
  INVX1 U211 ( .A(n50), .Y(n49) );
  NAND2XL U212 ( .A(B[26]), .B(A[26]), .Y(n75) );
  NAND2X1 U213 ( .A(A[24]), .B(B[24]), .Y(n73) );
  OR2X2 U214 ( .A(A[21]), .B(B[21]), .Y(n115) );
  NAND2X1 U215 ( .A(B[20]), .B(A[20]), .Y(n103) );
  NAND2X1 U216 ( .A(B[16]), .B(A[16]), .Y(n135) );
  NAND2X1 U217 ( .A(B[17]), .B(A[17]), .Y(n136) );
  NAND2X1 U218 ( .A(B[18]), .B(A[18]), .Y(n137) );
  NAND2X1 U219 ( .A(B[21]), .B(A[21]), .Y(n104) );
  OR2X2 U220 ( .A(A[16]), .B(B[16]), .Y(n128) );
  OR2X2 U221 ( .A(A[15]), .B(B[15]), .Y(n174) );
  OR2X2 U222 ( .A(A[14]), .B(B[14]), .Y(n173) );
  OR2X2 U223 ( .A(A[17]), .B(B[17]), .Y(n129) );
  OR2X2 U224 ( .A(A[20]), .B(B[20]), .Y(n119) );
  OR2X2 U225 ( .A(A[18]), .B(B[18]), .Y(n143) );
  NOR2X1 U226 ( .A(A[9]), .B(B[9]), .Y(n5) );
  NAND2X1 U227 ( .A(B[12]), .B(A[12]), .Y(n158) );
  OR2X2 U228 ( .A(A[11]), .B(B[11]), .Y(n192) );
  NAND2X1 U229 ( .A(B[10]), .B(A[10]), .Y(n202) );
  OR2X2 U230 ( .A(A[7]), .B(B[7]), .Y(n208) );
  OR2X2 U231 ( .A(A[12]), .B(B[12]), .Y(n172) );
  NOR2X1 U232 ( .A(A[5]), .B(B[5]), .Y(n6) );
  NOR2X1 U233 ( .A(A[4]), .B(B[4]), .Y(n7) );
  NAND2X1 U234 ( .A(B[4]), .B(A[4]), .Y(n30) );
  NAND2X1 U235 ( .A(B[8]), .B(A[8]), .Y(n14) );
  NAND2X1 U236 ( .A(B[5]), .B(A[5]), .Y(n27) );
  NAND2X1 U237 ( .A(B[2]), .B(A[2]), .Y(n37) );
  NAND2X1 U238 ( .A(B[6]), .B(A[6]), .Y(n22) );
  OR2X2 U239 ( .A(A[6]), .B(B[6]), .Y(n25) );
  NOR2X1 U240 ( .A(A[3]), .B(B[3]), .Y(n8) );
  OR2X2 U241 ( .A(A[8]), .B(B[8]), .Y(n198) );
  OR2X2 U242 ( .A(A[1]), .B(B[1]), .Y(n57) );
  NAND2X1 U243 ( .A(B[1]), .B(A[1]), .Y(n59) );
  NAND2X1 U244 ( .A(B[0]), .B(A[0]), .Y(n140) );
  AND2X2 U245 ( .A(n140), .B(n215), .Y(SUM[0]) );
  OR2X2 U246 ( .A(A[0]), .B(B[0]), .Y(n215) );
  CLKINVX3 U247 ( .A(n62), .Y(n51) );
  OR2X4 U248 ( .A(A[28]), .B(B[28]), .Y(n62) );
endmodule


module message_schedule ( clk, reset, data, write_enable, inner_busy, Wt );
  input [7:0] data;
  output [31:0] Wt;
  input clk, reset, write_enable, inner_busy;
  wire   n2228, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451,
         N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462,
         N463, N464, N465, N474, N475, N476, N477, N478, N479, N480, N481,
         N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492,
         N493, N494, N495, N496, N497, N506, N507, N508, N509, N510, N511,
         N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522,
         N523, N524, N525, N526, N527, N528, N529, N538, N539, N540, N541,
         N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552,
         N553, N554, N555, N556, N557, N558, N559, N560, N561, N570, N571,
         N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582,
         N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593,
         N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612,
         N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623,
         N624, N625, N634, N635, N636, N637, N638, N639, N640, N641, N642,
         N643, N644, N645, N646, N647, N648, N649, N650, N651, N652, N653,
         N654, N655, N656, N657, N666, N667, N668, N669, N670, N671, N672,
         N673, N674, N675, N676, N677, N678, N679, N680, N681, N682, N683,
         N684, N685, N686, N687, N688, N689, N698, N699, N700, N701, N702,
         N703, N704, N705, N706, N707, N708, N709, N710, N711, N712, N713,
         N714, N715, N716, N717, N718, N719, N720, N721, N730, N731, N732,
         N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743,
         N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N762,
         N763, N764, N765, N766, N767, N768, N769, N770, N771, N772, N773,
         N774, N775, N776, N777, N778, N779, N780, N781, N782, N783, N784,
         N785, N794, N795, N796, N797, N798, N799, N800, N801, N802, N803,
         N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814,
         N815, N816, N817, N826, N827, N828, N829, N830, N831, N832, N833,
         N834, N835, N836, N837, N838, N839, N840, N841, N842, N843, N844,
         N845, N846, N847, N848, N849, N858, N859, N860, N861, N862, N863,
         N864, N865, N866, N867, N868, N869, N870, N871, N872, N873, N874,
         N875, N876, N877, N878, N879, N880, N881, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N911, N912, N913, N922, N923,
         N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934,
         N935, N936, N937, N938, N939, N940, N941, N942, N943, N944, N945,
         N1462, N1463, N1464, N1465, N1466, N1467, N1468, N2133, N2134, N2135,
         N2136, N2137, N2138, N2139, N2140, N2141, N2142, N2143, N2144, N2145,
         N2146, N2147, N2148, N2149, N2150, N2151, N2152, N2153, N2154, N2155,
         N2156, N2157, N2158, N2159, N2160, N2161, N2162, N2163, N2164, N2171,
         N2172, N2173, N2174, N2175, N2176, N2177, n1056, n1057, n1059, n1060,
         n1061, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1266, n1267, n1268, n1269, n1270, n1271, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1731, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2064, n2065, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, N86, N85, N84, N83, N82,
         N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68,
         N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54,
         N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40,
         N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26,
         N25, N24, N23, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n58, n59, n60, n61, n417, n418, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1058, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1149, n1265, n1272, n1300, n1704, n1705, n1706, n1707,
         n1708, n1717, n1718, n1719, n1730, n1732, n1733, n1734, n1735, n1744,
         n1755, n1766, n1777, n1788, n1799, n1810, n1821, n1832, n1843, n1854,
         n1865, n1876, n1887, n1898, n1909, n1920, n1931, n1942, n1953, n1964,
         n1975, n1986, n1997, n2008, n2019, n2030, n2041, n2052, n2063, n2066,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224;
  wire   [31:0] R14;
  wire   [31:0] sigma0;
  wire   [31:0] R1;
  wire   [31:0] sigma1;
  wire   [31:0] R15;
  wire   [31:0] R6;
  wire   [31:0] logic_result;
  wire   [127:0] buffer;
  wire   [6:0] counter1;
  wire   [6:0] counter2;
  wire   [31:0] R2;
  wire   [31:0] R3;
  wire   [31:0] R4;
  wire   [31:0] R5;
  wire   [31:0] R7;
  wire   [31:0] R8;
  wire   [31:0] R9;
  wire   [31:0] R10;
  wire   [31:0] R11;
  wire   [31:0] R12;
  wire   [31:0] R13;

  DFFHQX4 Wt_reg_15_ ( .D(N2148), .CK(clk), .Q(Wt[15]) );
  DFFHQX4 Wt_reg_14_ ( .D(N2147), .CK(clk), .Q(Wt[14]) );
  DFFHQX4 Wt_reg_12_ ( .D(N2145), .CK(clk), .Q(Wt[12]) );
  DFFHQX4 Wt_reg_11_ ( .D(N2144), .CK(clk), .Q(Wt[11]) );
  DFFHQX4 Wt_reg_10_ ( .D(N2143), .CK(clk), .Q(Wt[10]) );
  DFFHQX4 Wt_reg_9_ ( .D(N2142), .CK(clk), .Q(Wt[9]) );
  DFFHQX4 Wt_reg_8_ ( .D(N2141), .CK(clk), .Q(Wt[8]) );
  DFFHQX4 Wt_reg_7_ ( .D(N2140), .CK(clk), .Q(Wt[7]) );
  DFFHQX4 Wt_reg_6_ ( .D(N2139), .CK(clk), .Q(Wt[6]) );
  DFFHQX4 Wt_reg_5_ ( .D(N2138), .CK(clk), .Q(Wt[5]) );
  DFFHQX4 Wt_reg_4_ ( .D(N2137), .CK(clk), .Q(Wt[4]) );
  DFFHQX4 Wt_reg_3_ ( .D(N2136), .CK(clk), .Q(Wt[3]) );
  DFFHQX4 Wt_reg_2_ ( .D(N2135), .CK(clk), .Q(Wt[2]) );
  DFFHQX4 Wt_reg_1_ ( .D(N2134), .CK(clk), .Q(Wt[1]) );
  DFFHQX4 Wt_reg_0_ ( .D(N2133), .CK(clk), .Q(n2228) );
  DFFTRX4 R6_reg_0_ ( .D(R5[0]), .RN(n550), .CK(clk), .Q(R6[0]) );
  DFFTRX4 R15_reg_0_ ( .D(R14[0]), .RN(n550), .CK(clk), .Q(R15[0]) );
  NOR2X4 U508 ( .A(n1476), .B(reset), .Y(n1477) );
  NOR2X4 U577 ( .A(n1549), .B(reset), .Y(n1550) );
  NOR2X4 U611 ( .A(n1585), .B(reset), .Y(n1586) );
  NOR2X4 U645 ( .A(n1620), .B(reset), .Y(n1621) );
  NOR2X4 U679 ( .A(n615), .B(reset), .Y(n1657) );
  AOI2BB1X4 U680 ( .A0N(n1689), .A1N(n1654), .B0(reset), .Y(n1656) );
  AND3X4 U682 ( .A(n1690), .B(n1440), .C(n1333), .Y(n1583) );
  AND3X4 U686 ( .A(n1153), .B(n1691), .C(write_enable), .Y(n1224) );
  AND2X2 U688 ( .A(n1694), .B(n1261), .Y(n1151) );
  AND2X2 U689 ( .A(n1695), .B(n1262), .Y(n1152) );
  AND2X2 U697 ( .A(n1155), .B(n1154), .Y(n1333) );
  AND2X2 U702 ( .A(n1698), .B(n1702), .Y(n1404) );
  AND2X2 U703 ( .A(n1698), .B(n1700), .Y(n1368) );
  AND2X2 U707 ( .A(n1702), .B(n1703), .Y(n1689) );
  AND2X2 U708 ( .A(n1703), .B(n1700), .Y(n1653) );
  AND2X2 U709 ( .A(n1582), .B(n1618), .Y(n1547) );
  AND2X2 U715 ( .A(n1702), .B(n1701), .Y(n1545) );
  AND2X2 U716 ( .A(n1700), .B(n1701), .Y(n1509) );
  AND2X2 U1102 ( .A(n2072), .B(n2073), .Y(n1714) );
  AND2X2 U1103 ( .A(n2074), .B(n2072), .Y(n1713) );
  AND2X2 U1105 ( .A(n2075), .B(n2073), .Y(n1716) );
  AND2X2 U1106 ( .A(n2074), .B(n2075), .Y(n1715) );
  AND2X2 U1115 ( .A(n2082), .B(n2072), .Y(n1726) );
  AND2X2 U1116 ( .A(n2072), .B(n2083), .Y(n1725) );
  AND2X2 U1119 ( .A(n2075), .B(n2082), .Y(n1728) );
  AND2X2 U1120 ( .A(n2075), .B(n2083), .Y(n1727) );
  AND2X2 U1124 ( .A(n2076), .B(n2083), .Y(n1729) );
  AND2X2 U1129 ( .A(n2083), .B(n2077), .Y(n1731) );
  AND2X2 U1135 ( .A(n2073), .B(n2077), .Y(n1720) );
  message_schedule_DW01_inc_0 add_564 ( .A(counter2), .SUM({N2177, N2176, 
        N2175, N2174, N2173, N2172, N2171}) );
  message_schedule_DW01_inc_1 add_461 ( .A(counter1), .SUM({N1468, N1467, 
        N1466, N1465, N1464, N1463, N1462}) );
  message_schedule_DW01_add_17 add_2_root_add_0_root_add_35_3 ( .A(R15), .B(R6), .SUM({N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, 
        N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, 
        N58, N57, N56, N55}) );
  message_schedule_DW01_add_20 add_1_root_add_0_root_add_35_3 ( .A(sigma1), 
        .B(sigma0), .SUM({N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, 
        N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, 
        N30, N29, N28, N27, N26, N25, N24, N23}) );
  message_schedule_DW01_add_21 add_0_root_add_0_root_add_35_3 ( .A({N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55}), .B({N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23}), .SUM(logic_result) );
  DFFHQXL buffer_reg_14__24_ ( .D(n2160), .CK(clk), .Q(buffer[8]) );
  DFFHQXL buffer_reg_14__25_ ( .D(n2159), .CK(clk), .Q(buffer[9]) );
  DFFHQXL buffer_reg_14__26_ ( .D(n2158), .CK(clk), .Q(buffer[10]) );
  DFFHQXL buffer_reg_14__27_ ( .D(n2157), .CK(clk), .Q(buffer[11]) );
  DFFHQXL buffer_reg_14__28_ ( .D(n2156), .CK(clk), .Q(buffer[12]) );
  DFFHQXL buffer_reg_14__29_ ( .D(n2155), .CK(clk), .Q(buffer[13]) );
  DFFHQXL buffer_reg_14__30_ ( .D(n2154), .CK(clk), .Q(buffer[14]) );
  DFFHQXL buffer_reg_14__31_ ( .D(n2153), .CK(clk), .Q(buffer[15]) );
  DFFHQXL buffer_reg_10__24_ ( .D(n1111), .CK(clk), .Q(buffer[40]) );
  DFFHQXL buffer_reg_10__25_ ( .D(n1110), .CK(clk), .Q(buffer[41]) );
  DFFHQXL buffer_reg_10__26_ ( .D(n1109), .CK(clk), .Q(buffer[42]) );
  DFFHQXL buffer_reg_10__27_ ( .D(n1108), .CK(clk), .Q(buffer[43]) );
  DFFHQXL buffer_reg_10__28_ ( .D(n1107), .CK(clk), .Q(buffer[44]) );
  DFFHQXL buffer_reg_10__29_ ( .D(n1106), .CK(clk), .Q(buffer[45]) );
  DFFHQXL buffer_reg_10__30_ ( .D(n1105), .CK(clk), .Q(buffer[46]) );
  DFFHQXL buffer_reg_10__31_ ( .D(n1104), .CK(clk), .Q(buffer[47]) );
  DFFHQXL buffer_reg_12__24_ ( .D(n2098), .CK(clk), .Q(buffer[24]) );
  DFFHQXL buffer_reg_12__25_ ( .D(n2097), .CK(clk), .Q(buffer[25]) );
  DFFHQXL buffer_reg_12__26_ ( .D(n2096), .CK(clk), .Q(buffer[26]) );
  DFFHQXL buffer_reg_12__27_ ( .D(n2095), .CK(clk), .Q(buffer[27]) );
  DFFHQXL buffer_reg_12__28_ ( .D(n2094), .CK(clk), .Q(buffer[28]) );
  DFFHQXL buffer_reg_12__29_ ( .D(n2093), .CK(clk), .Q(buffer[29]) );
  DFFHQXL buffer_reg_12__30_ ( .D(n2092), .CK(clk), .Q(buffer[30]) );
  DFFHQXL buffer_reg_12__31_ ( .D(n2091), .CK(clk), .Q(buffer[31]) );
  DFFHQXL buffer_reg_8__24_ ( .D(n1044), .CK(clk), .Q(buffer[56]) );
  DFFHQXL buffer_reg_8__25_ ( .D(n1043), .CK(clk), .Q(buffer[57]) );
  DFFHQXL buffer_reg_8__26_ ( .D(n1042), .CK(clk), .Q(buffer[58]) );
  DFFHQXL buffer_reg_8__27_ ( .D(n1041), .CK(clk), .Q(buffer[59]) );
  DFFHQXL buffer_reg_8__28_ ( .D(n1040), .CK(clk), .Q(buffer[60]) );
  DFFHQXL buffer_reg_8__29_ ( .D(n1039), .CK(clk), .Q(buffer[61]) );
  DFFHQXL buffer_reg_8__30_ ( .D(n1038), .CK(clk), .Q(buffer[62]) );
  DFFHQXL buffer_reg_8__31_ ( .D(n1037), .CK(clk), .Q(buffer[63]) );
  DFFHQXL buffer_reg_15__24_ ( .D(n2191), .CK(clk), .Q(buffer[0]) );
  DFFHQXL buffer_reg_15__25_ ( .D(n2190), .CK(clk), .Q(buffer[1]) );
  DFFHQXL buffer_reg_15__26_ ( .D(n2189), .CK(clk), .Q(buffer[2]) );
  DFFHQXL buffer_reg_15__27_ ( .D(n2188), .CK(clk), .Q(buffer[3]) );
  DFFHQXL buffer_reg_15__28_ ( .D(n2187), .CK(clk), .Q(buffer[4]) );
  DFFHQXL buffer_reg_15__29_ ( .D(n2186), .CK(clk), .Q(buffer[5]) );
  DFFHQXL buffer_reg_15__30_ ( .D(n2185), .CK(clk), .Q(buffer[6]) );
  DFFHQXL buffer_reg_15__31_ ( .D(n2184), .CK(clk), .Q(buffer[7]) );
  DFFHQXL buffer_reg_11__24_ ( .D(n1876), .CK(clk), .Q(buffer[32]) );
  DFFHQXL buffer_reg_11__25_ ( .D(n1865), .CK(clk), .Q(buffer[33]) );
  DFFHQXL buffer_reg_11__26_ ( .D(n1854), .CK(clk), .Q(buffer[34]) );
  DFFHQXL buffer_reg_11__27_ ( .D(n1843), .CK(clk), .Q(buffer[35]) );
  DFFHQXL buffer_reg_11__28_ ( .D(n1832), .CK(clk), .Q(buffer[36]) );
  DFFHQXL buffer_reg_11__29_ ( .D(n1821), .CK(clk), .Q(buffer[37]) );
  DFFHQXL buffer_reg_11__30_ ( .D(n1810), .CK(clk), .Q(buffer[38]) );
  DFFHQXL buffer_reg_11__31_ ( .D(n1799), .CK(clk), .Q(buffer[39]) );
  DFFHQXL buffer_reg_13__24_ ( .D(n2129), .CK(clk), .Q(buffer[16]) );
  DFFHQXL buffer_reg_13__25_ ( .D(n2128), .CK(clk), .Q(buffer[17]) );
  DFFHQXL buffer_reg_13__26_ ( .D(n2127), .CK(clk), .Q(buffer[18]) );
  DFFHQXL buffer_reg_13__27_ ( .D(n2126), .CK(clk), .Q(buffer[19]) );
  DFFHQXL buffer_reg_13__28_ ( .D(n2125), .CK(clk), .Q(buffer[20]) );
  DFFHQXL buffer_reg_13__29_ ( .D(n2124), .CK(clk), .Q(buffer[21]) );
  DFFHQXL buffer_reg_13__30_ ( .D(n2123), .CK(clk), .Q(buffer[22]) );
  DFFHQXL buffer_reg_13__31_ ( .D(n2122), .CK(clk), .Q(buffer[23]) );
  DFFHQXL buffer_reg_9__24_ ( .D(n1080), .CK(clk), .Q(buffer[48]) );
  DFFHQXL buffer_reg_9__25_ ( .D(n1079), .CK(clk), .Q(buffer[49]) );
  DFFHQXL buffer_reg_9__26_ ( .D(n1078), .CK(clk), .Q(buffer[50]) );
  DFFHQXL buffer_reg_9__27_ ( .D(n1077), .CK(clk), .Q(buffer[51]) );
  DFFHQXL buffer_reg_9__28_ ( .D(n1076), .CK(clk), .Q(buffer[52]) );
  DFFHQXL buffer_reg_9__29_ ( .D(n1075), .CK(clk), .Q(buffer[53]) );
  DFFHQXL buffer_reg_9__30_ ( .D(n1074), .CK(clk), .Q(buffer[54]) );
  DFFHQXL buffer_reg_9__31_ ( .D(n1073), .CK(clk), .Q(buffer[55]) );
  DFFHQXL buffer_reg_14__0_ ( .D(n2220), .CK(clk), .Q(N890) );
  DFFHQXL buffer_reg_14__1_ ( .D(n2152), .CK(clk), .Q(N891) );
  DFFHQXL buffer_reg_14__2_ ( .D(n2151), .CK(clk), .Q(N892) );
  DFFHQXL buffer_reg_14__3_ ( .D(n2150), .CK(clk), .Q(N893) );
  DFFHQXL buffer_reg_14__4_ ( .D(n2149), .CK(clk), .Q(N894) );
  DFFHQXL buffer_reg_14__5_ ( .D(n2148), .CK(clk), .Q(N895) );
  DFFHQXL buffer_reg_14__6_ ( .D(n2147), .CK(clk), .Q(N896) );
  DFFHQXL buffer_reg_14__7_ ( .D(n2146), .CK(clk), .Q(N897) );
  DFFHQXL buffer_reg_14__8_ ( .D(n2176), .CK(clk), .Q(N898) );
  DFFHQXL buffer_reg_14__9_ ( .D(n2175), .CK(clk), .Q(N899) );
  DFFHQXL buffer_reg_14__10_ ( .D(n2174), .CK(clk), .Q(N900) );
  DFFHQXL buffer_reg_14__11_ ( .D(n2173), .CK(clk), .Q(N901) );
  DFFHQXL buffer_reg_14__12_ ( .D(n2172), .CK(clk), .Q(N902) );
  DFFHQXL buffer_reg_14__13_ ( .D(n2171), .CK(clk), .Q(N903) );
  DFFHQXL buffer_reg_14__14_ ( .D(n2170), .CK(clk), .Q(N904) );
  DFFHQXL buffer_reg_14__15_ ( .D(n2169), .CK(clk), .Q(N905) );
  DFFHQXL buffer_reg_14__16_ ( .D(n2168), .CK(clk), .Q(N906) );
  DFFHQXL buffer_reg_14__17_ ( .D(n2167), .CK(clk), .Q(N907) );
  DFFHQXL buffer_reg_14__18_ ( .D(n2166), .CK(clk), .Q(N908) );
  DFFHQXL buffer_reg_14__19_ ( .D(n2165), .CK(clk), .Q(N909) );
  DFFHQXL buffer_reg_14__20_ ( .D(n2164), .CK(clk), .Q(N910) );
  DFFHQXL buffer_reg_14__21_ ( .D(n2163), .CK(clk), .Q(N911) );
  DFFHQXL buffer_reg_14__22_ ( .D(n2162), .CK(clk), .Q(N912) );
  DFFHQXL buffer_reg_14__23_ ( .D(n2161), .CK(clk), .Q(N913) );
  DFFHQXL buffer_reg_10__0_ ( .D(n2223), .CK(clk), .Q(N762) );
  DFFHQXL buffer_reg_10__1_ ( .D(n1103), .CK(clk), .Q(N763) );
  DFFHQXL buffer_reg_10__2_ ( .D(n1102), .CK(clk), .Q(N764) );
  DFFHQXL buffer_reg_10__3_ ( .D(n1101), .CK(clk), .Q(N765) );
  DFFHQXL buffer_reg_10__4_ ( .D(n1100), .CK(clk), .Q(N766) );
  DFFHQXL buffer_reg_10__5_ ( .D(n1099), .CK(clk), .Q(N767) );
  DFFHQXL buffer_reg_10__6_ ( .D(n1098), .CK(clk), .Q(N768) );
  DFFHQXL buffer_reg_10__7_ ( .D(n1097), .CK(clk), .Q(N769) );
  DFFHQXL buffer_reg_10__8_ ( .D(n1733), .CK(clk), .Q(N770) );
  DFFHQXL buffer_reg_10__9_ ( .D(n1732), .CK(clk), .Q(N771) );
  DFFHQXL buffer_reg_10__10_ ( .D(n1730), .CK(clk), .Q(N772) );
  DFFHQXL buffer_reg_10__11_ ( .D(n1719), .CK(clk), .Q(N773) );
  DFFHQXL buffer_reg_10__12_ ( .D(n1718), .CK(clk), .Q(N774) );
  DFFHQXL buffer_reg_10__13_ ( .D(n1717), .CK(clk), .Q(N775) );
  DFFHQXL buffer_reg_10__14_ ( .D(n1708), .CK(clk), .Q(N776) );
  DFFHQXL buffer_reg_10__15_ ( .D(n1707), .CK(clk), .Q(N777) );
  DFFHQXL buffer_reg_10__16_ ( .D(n1706), .CK(clk), .Q(N778) );
  DFFHQXL buffer_reg_10__17_ ( .D(n1705), .CK(clk), .Q(N779) );
  DFFHQXL buffer_reg_10__18_ ( .D(n1704), .CK(clk), .Q(N780) );
  DFFHQXL buffer_reg_10__19_ ( .D(n1300), .CK(clk), .Q(N781) );
  DFFHQXL buffer_reg_10__20_ ( .D(n1272), .CK(clk), .Q(N782) );
  DFFHQXL buffer_reg_10__21_ ( .D(n1265), .CK(clk), .Q(N783) );
  DFFHQXL buffer_reg_10__22_ ( .D(n1149), .CK(clk), .Q(N784) );
  DFFHQXL buffer_reg_10__23_ ( .D(n1112), .CK(clk), .Q(N785) );
  DFFHQXL buffer_reg_12__0_ ( .D(n2222), .CK(clk), .Q(N826) );
  DFFHQXL buffer_reg_12__1_ ( .D(n2090), .CK(clk), .Q(N827) );
  DFFHQXL buffer_reg_12__2_ ( .D(n2089), .CK(clk), .Q(N828) );
  DFFHQXL buffer_reg_12__3_ ( .D(n2088), .CK(clk), .Q(N829) );
  DFFHQXL buffer_reg_12__4_ ( .D(n2087), .CK(clk), .Q(N830) );
  DFFHQXL buffer_reg_12__5_ ( .D(n2086), .CK(clk), .Q(N831) );
  DFFHQXL buffer_reg_12__6_ ( .D(n2066), .CK(clk), .Q(N832) );
  DFFHQXL buffer_reg_12__7_ ( .D(n2063), .CK(clk), .Q(N833) );
  DFFHQXL buffer_reg_12__8_ ( .D(n2114), .CK(clk), .Q(N834) );
  DFFHQXL buffer_reg_12__9_ ( .D(n2113), .CK(clk), .Q(N835) );
  DFFHQXL buffer_reg_12__10_ ( .D(n2112), .CK(clk), .Q(N836) );
  DFFHQXL buffer_reg_12__11_ ( .D(n2111), .CK(clk), .Q(N837) );
  DFFHQXL buffer_reg_12__12_ ( .D(n2110), .CK(clk), .Q(N838) );
  DFFHQXL buffer_reg_12__13_ ( .D(n2109), .CK(clk), .Q(N839) );
  DFFHQXL buffer_reg_12__14_ ( .D(n2108), .CK(clk), .Q(N840) );
  DFFHQXL buffer_reg_12__15_ ( .D(n2107), .CK(clk), .Q(N841) );
  DFFHQXL buffer_reg_12__16_ ( .D(n2106), .CK(clk), .Q(N842) );
  DFFHQXL buffer_reg_12__17_ ( .D(n2105), .CK(clk), .Q(N843) );
  DFFHQXL buffer_reg_12__18_ ( .D(n2104), .CK(clk), .Q(N844) );
  DFFHQXL buffer_reg_12__19_ ( .D(n2103), .CK(clk), .Q(N845) );
  DFFHQXL buffer_reg_12__20_ ( .D(n2102), .CK(clk), .Q(N846) );
  DFFHQXL buffer_reg_12__21_ ( .D(n2101), .CK(clk), .Q(N847) );
  DFFHQXL buffer_reg_12__22_ ( .D(n2100), .CK(clk), .Q(N848) );
  DFFHQXL buffer_reg_12__23_ ( .D(n2099), .CK(clk), .Q(N849) );
  DFFHQX1 buffer_reg_0__12_ ( .D(n809), .CK(clk), .Q(N454) );
  DFFHQX1 buffer_reg_0__13_ ( .D(n808), .CK(clk), .Q(N455) );
  DFFHQX1 buffer_reg_0__14_ ( .D(n807), .CK(clk), .Q(N456) );
  DFFHQX1 buffer_reg_0__15_ ( .D(n806), .CK(clk), .Q(N457) );
  DFFHQX1 buffer_reg_0__16_ ( .D(n805), .CK(clk), .Q(N458) );
  DFFHQX1 buffer_reg_0__17_ ( .D(n804), .CK(clk), .Q(N459) );
  DFFHQX1 buffer_reg_0__18_ ( .D(n803), .CK(clk), .Q(N460) );
  DFFHQX1 buffer_reg_0__19_ ( .D(n802), .CK(clk), .Q(N461) );
  DFFHQX1 buffer_reg_0__20_ ( .D(n801), .CK(clk), .Q(N462) );
  DFFHQX1 buffer_reg_0__21_ ( .D(n800), .CK(clk), .Q(N463) );
  DFFHQX1 buffer_reg_0__22_ ( .D(n799), .CK(clk), .Q(N464) );
  DFFHQX1 buffer_reg_0__23_ ( .D(n798), .CK(clk), .Q(N465) );
  DFFHQXL buffer_reg_8__0_ ( .D(n2211), .CK(clk), .Q(N698) );
  DFFHQXL buffer_reg_8__1_ ( .D(n1036), .CK(clk), .Q(N699) );
  DFFHQXL buffer_reg_8__2_ ( .D(n1035), .CK(clk), .Q(N700) );
  DFFHQXL buffer_reg_8__3_ ( .D(n1034), .CK(clk), .Q(N701) );
  DFFHQXL buffer_reg_8__4_ ( .D(n1033), .CK(clk), .Q(N702) );
  DFFHQXL buffer_reg_8__5_ ( .D(n1032), .CK(clk), .Q(N703) );
  DFFHQXL buffer_reg_8__6_ ( .D(n1031), .CK(clk), .Q(N704) );
  DFFHQXL buffer_reg_8__7_ ( .D(n1030), .CK(clk), .Q(N705) );
  DFFHQXL buffer_reg_8__8_ ( .D(n1065), .CK(clk), .Q(N706) );
  DFFHQXL buffer_reg_8__9_ ( .D(n1064), .CK(clk), .Q(N707) );
  DFFHQXL buffer_reg_8__10_ ( .D(n1063), .CK(clk), .Q(N708) );
  DFFHQXL buffer_reg_8__11_ ( .D(n1062), .CK(clk), .Q(N709) );
  DFFHQXL buffer_reg_8__12_ ( .D(n1058), .CK(clk), .Q(N710) );
  DFFHQXL buffer_reg_8__13_ ( .D(n1055), .CK(clk), .Q(N711) );
  DFFHQXL buffer_reg_8__14_ ( .D(n1054), .CK(clk), .Q(N712) );
  DFFHQXL buffer_reg_8__15_ ( .D(n1053), .CK(clk), .Q(N713) );
  DFFHQXL buffer_reg_8__16_ ( .D(n1052), .CK(clk), .Q(N714) );
  DFFHQXL buffer_reg_8__17_ ( .D(n1051), .CK(clk), .Q(N715) );
  DFFHQXL buffer_reg_8__18_ ( .D(n1050), .CK(clk), .Q(N716) );
  DFFHQXL buffer_reg_8__19_ ( .D(n1049), .CK(clk), .Q(N717) );
  DFFHQXL buffer_reg_8__20_ ( .D(n1048), .CK(clk), .Q(N718) );
  DFFHQXL buffer_reg_8__21_ ( .D(n1047), .CK(clk), .Q(N719) );
  DFFHQXL buffer_reg_8__22_ ( .D(n1046), .CK(clk), .Q(N720) );
  DFFHQXL buffer_reg_8__23_ ( .D(n1045), .CK(clk), .Q(N721) );
  DFFHQXL buffer_reg_15__0_ ( .D(n2219), .CK(clk), .Q(N922) );
  DFFHQXL buffer_reg_15__1_ ( .D(n2183), .CK(clk), .Q(N923) );
  DFFHQXL buffer_reg_15__2_ ( .D(n2182), .CK(clk), .Q(N924) );
  DFFHQXL buffer_reg_15__3_ ( .D(n2181), .CK(clk), .Q(N925) );
  DFFHQXL buffer_reg_15__4_ ( .D(n2180), .CK(clk), .Q(N926) );
  DFFHQXL buffer_reg_15__5_ ( .D(n2179), .CK(clk), .Q(N927) );
  DFFHQXL buffer_reg_15__6_ ( .D(n2178), .CK(clk), .Q(N928) );
  DFFHQXL buffer_reg_15__7_ ( .D(n2177), .CK(clk), .Q(N929) );
  DFFHQXL buffer_reg_15__8_ ( .D(n2207), .CK(clk), .Q(N930) );
  DFFHQXL buffer_reg_15__9_ ( .D(n2206), .CK(clk), .Q(N931) );
  DFFHQXL buffer_reg_15__10_ ( .D(n2205), .CK(clk), .Q(N932) );
  DFFHQXL buffer_reg_15__11_ ( .D(n2204), .CK(clk), .Q(N933) );
  DFFHQXL buffer_reg_15__12_ ( .D(n2203), .CK(clk), .Q(N934) );
  DFFHQXL buffer_reg_15__13_ ( .D(n2202), .CK(clk), .Q(N935) );
  DFFHQXL buffer_reg_15__14_ ( .D(n2201), .CK(clk), .Q(N936) );
  DFFHQXL buffer_reg_15__15_ ( .D(n2200), .CK(clk), .Q(N937) );
  DFFHQXL buffer_reg_15__16_ ( .D(n2199), .CK(clk), .Q(N938) );
  DFFHQXL buffer_reg_15__17_ ( .D(n2198), .CK(clk), .Q(N939) );
  DFFHQXL buffer_reg_15__18_ ( .D(n2197), .CK(clk), .Q(N940) );
  DFFHQXL buffer_reg_15__19_ ( .D(n2196), .CK(clk), .Q(N941) );
  DFFHQXL buffer_reg_15__20_ ( .D(n2195), .CK(clk), .Q(N942) );
  DFFHQXL buffer_reg_15__21_ ( .D(n2194), .CK(clk), .Q(N943) );
  DFFHQXL buffer_reg_15__22_ ( .D(n2193), .CK(clk), .Q(N944) );
  DFFHQXL buffer_reg_15__23_ ( .D(n2192), .CK(clk), .Q(N945) );
  DFFHQXL buffer_reg_11__0_ ( .D(n2224), .CK(clk), .Q(N794) );
  DFFHQXL buffer_reg_11__1_ ( .D(n1788), .CK(clk), .Q(N795) );
  DFFHQXL buffer_reg_11__2_ ( .D(n1777), .CK(clk), .Q(N796) );
  DFFHQXL buffer_reg_11__3_ ( .D(n1766), .CK(clk), .Q(N797) );
  DFFHQXL buffer_reg_11__4_ ( .D(n1755), .CK(clk), .Q(N798) );
  DFFHQXL buffer_reg_11__5_ ( .D(n1744), .CK(clk), .Q(N799) );
  DFFHQXL buffer_reg_11__6_ ( .D(n1735), .CK(clk), .Q(N800) );
  DFFHQXL buffer_reg_11__7_ ( .D(n1734), .CK(clk), .Q(N801) );
  DFFHQXL buffer_reg_11__8_ ( .D(n2052), .CK(clk), .Q(N802) );
  DFFHQXL buffer_reg_11__9_ ( .D(n2041), .CK(clk), .Q(N803) );
  DFFHQXL buffer_reg_11__10_ ( .D(n2030), .CK(clk), .Q(N804) );
  DFFHQXL buffer_reg_11__11_ ( .D(n2019), .CK(clk), .Q(N805) );
  DFFHQXL buffer_reg_11__12_ ( .D(n2008), .CK(clk), .Q(N806) );
  DFFHQXL buffer_reg_11__13_ ( .D(n1997), .CK(clk), .Q(N807) );
  DFFHQXL buffer_reg_11__14_ ( .D(n1986), .CK(clk), .Q(N808) );
  DFFHQXL buffer_reg_11__15_ ( .D(n1975), .CK(clk), .Q(N809) );
  DFFHQXL buffer_reg_11__16_ ( .D(n1964), .CK(clk), .Q(N810) );
  DFFHQXL buffer_reg_11__17_ ( .D(n1953), .CK(clk), .Q(N811) );
  DFFHQXL buffer_reg_11__18_ ( .D(n1942), .CK(clk), .Q(N812) );
  DFFHQXL buffer_reg_11__19_ ( .D(n1931), .CK(clk), .Q(N813) );
  DFFHQXL buffer_reg_11__20_ ( .D(n1920), .CK(clk), .Q(N814) );
  DFFHQXL buffer_reg_11__21_ ( .D(n1909), .CK(clk), .Q(N815) );
  DFFHQXL buffer_reg_11__22_ ( .D(n1898), .CK(clk), .Q(N816) );
  DFFHQXL buffer_reg_11__23_ ( .D(n1887), .CK(clk), .Q(N817) );
  DFFHQXL buffer_reg_13__0_ ( .D(n2221), .CK(clk), .Q(N858) );
  DFFHQXL buffer_reg_13__1_ ( .D(n2121), .CK(clk), .Q(N859) );
  DFFHQXL buffer_reg_13__2_ ( .D(n2120), .CK(clk), .Q(N860) );
  DFFHQXL buffer_reg_13__3_ ( .D(n2119), .CK(clk), .Q(N861) );
  DFFHQXL buffer_reg_13__4_ ( .D(n2118), .CK(clk), .Q(N862) );
  DFFHQXL buffer_reg_13__5_ ( .D(n2117), .CK(clk), .Q(N863) );
  DFFHQXL buffer_reg_13__6_ ( .D(n2116), .CK(clk), .Q(N864) );
  DFFHQXL buffer_reg_13__7_ ( .D(n2115), .CK(clk), .Q(N865) );
  DFFHQXL buffer_reg_13__8_ ( .D(n2145), .CK(clk), .Q(N866) );
  DFFHQXL buffer_reg_13__9_ ( .D(n2144), .CK(clk), .Q(N867) );
  DFFHQXL buffer_reg_13__10_ ( .D(n2143), .CK(clk), .Q(N868) );
  DFFHQXL buffer_reg_13__11_ ( .D(n2142), .CK(clk), .Q(N869) );
  DFFHQXL buffer_reg_13__12_ ( .D(n2141), .CK(clk), .Q(N870) );
  DFFHQXL buffer_reg_13__13_ ( .D(n2140), .CK(clk), .Q(N871) );
  DFFHQXL buffer_reg_13__14_ ( .D(n2139), .CK(clk), .Q(N872) );
  DFFHQXL buffer_reg_13__15_ ( .D(n2138), .CK(clk), .Q(N873) );
  DFFHQXL buffer_reg_13__16_ ( .D(n2137), .CK(clk), .Q(N874) );
  DFFHQXL buffer_reg_13__17_ ( .D(n2136), .CK(clk), .Q(N875) );
  DFFHQXL buffer_reg_13__18_ ( .D(n2135), .CK(clk), .Q(N876) );
  DFFHQXL buffer_reg_13__19_ ( .D(n2134), .CK(clk), .Q(N877) );
  DFFHQXL buffer_reg_13__20_ ( .D(n2133), .CK(clk), .Q(N878) );
  DFFHQXL buffer_reg_13__21_ ( .D(n2132), .CK(clk), .Q(N879) );
  DFFHQXL buffer_reg_13__22_ ( .D(n2131), .CK(clk), .Q(N880) );
  DFFHQXL buffer_reg_13__23_ ( .D(n2130), .CK(clk), .Q(N881) );
  DFFHQXL buffer_reg_9__0_ ( .D(n2210), .CK(clk), .Q(N730) );
  DFFHQXL buffer_reg_9__1_ ( .D(n1072), .CK(clk), .Q(N731) );
  DFFHQXL buffer_reg_9__2_ ( .D(n1071), .CK(clk), .Q(N732) );
  DFFHQXL buffer_reg_9__3_ ( .D(n1070), .CK(clk), .Q(N733) );
  DFFHQXL buffer_reg_9__4_ ( .D(n1069), .CK(clk), .Q(N734) );
  DFFHQXL buffer_reg_9__5_ ( .D(n1068), .CK(clk), .Q(N735) );
  DFFHQXL buffer_reg_9__6_ ( .D(n1067), .CK(clk), .Q(N736) );
  DFFHQXL buffer_reg_9__7_ ( .D(n1066), .CK(clk), .Q(N737) );
  DFFHQXL buffer_reg_9__8_ ( .D(n1096), .CK(clk), .Q(N738) );
  DFFHQXL buffer_reg_9__9_ ( .D(n1095), .CK(clk), .Q(N739) );
  DFFHQXL buffer_reg_9__10_ ( .D(n1094), .CK(clk), .Q(N740) );
  DFFHQXL buffer_reg_9__11_ ( .D(n1093), .CK(clk), .Q(N741) );
  DFFHQXL buffer_reg_9__12_ ( .D(n1092), .CK(clk), .Q(N742) );
  DFFHQXL buffer_reg_9__13_ ( .D(n1091), .CK(clk), .Q(N743) );
  DFFHQXL buffer_reg_9__14_ ( .D(n1090), .CK(clk), .Q(N744) );
  DFFHQXL buffer_reg_9__15_ ( .D(n1089), .CK(clk), .Q(N745) );
  DFFHQXL buffer_reg_9__16_ ( .D(n1088), .CK(clk), .Q(N746) );
  DFFHQXL buffer_reg_9__17_ ( .D(n1087), .CK(clk), .Q(N747) );
  DFFHQXL buffer_reg_9__18_ ( .D(n1086), .CK(clk), .Q(N748) );
  DFFHQXL buffer_reg_9__19_ ( .D(n1085), .CK(clk), .Q(N749) );
  DFFHQXL buffer_reg_9__20_ ( .D(n1084), .CK(clk), .Q(N750) );
  DFFHQXL buffer_reg_9__21_ ( .D(n1083), .CK(clk), .Q(N751) );
  DFFHQXL buffer_reg_9__22_ ( .D(n1082), .CK(clk), .Q(N752) );
  DFFHQXL buffer_reg_9__23_ ( .D(n1081), .CK(clk), .Q(N753) );
  DFFTRX1 R15_reg_31_ ( .D(R14[31]), .RN(n581), .CK(clk), .Q(R15[31]) );
  DFFTRX1 R15_reg_29_ ( .D(R14[29]), .RN(n583), .CK(clk), .Q(R15[29]) );
  DFFTRX1 R15_reg_30_ ( .D(R14[30]), .RN(n584), .CK(clk), .Q(R15[30]) );
  DFFTRX1 counter1_reg_1_ ( .D(N1463), .RN(n2085), .CK(clk), .Q(counter1[1])
         );
  DFFTRX1 counter1_reg_0_ ( .D(N1462), .RN(n2085), .CK(clk), .Q(counter1[0])
         );
  DFFTRX1 R6_reg_31_ ( .D(R5[31]), .RN(n585), .CK(clk), .Q(R6[31]) );
  DFFTRX1 R6_reg_29_ ( .D(R5[29]), .RN(n584), .CK(clk), .Q(R6[29]) );
  DFFTRX1 R6_reg_30_ ( .D(R5[30]), .RN(n580), .CK(clk), .Q(R6[30]) );
  DFFTRX1 counter2_reg_4_ ( .D(N2175), .RN(n582), .CK(clk), .Q(counter2[4]) );
  DFFTRX1 counter2_reg_6_ ( .D(N2177), .RN(n585), .CK(clk), .Q(counter2[6]) );
  DFFTRX1 counter2_reg_5_ ( .D(N2176), .RN(n585), .CK(clk), .Q(counter2[5]) );
  DFFTRX1 R15_reg_28_ ( .D(R14[28]), .RN(n582), .CK(clk), .Q(R15[28]) );
  DFFTRX1 R15_reg_27_ ( .D(R14[27]), .RN(n585), .CK(clk), .Q(R15[27]) );
  DFFTRX1 R15_reg_26_ ( .D(R14[26]), .RN(n580), .CK(clk), .Q(R15[26]) );
  DFFTRX1 R6_reg_28_ ( .D(R5[28]), .RN(n582), .CK(clk), .Q(R6[28]) );
  DFFTRX1 R6_reg_27_ ( .D(R5[27]), .RN(n581), .CK(clk), .Q(R6[27]) );
  DFFTRX1 R6_reg_26_ ( .D(R5[26]), .RN(n584), .CK(clk), .Q(R6[26]) );
  DFFTRX1 counter1_reg_6_ ( .D(N1468), .RN(n2085), .CK(clk), .Q(counter1[6])
         );
  DFFTRX1 counter2_reg_1_ ( .D(N2172), .RN(n580), .CK(clk), .Q(counter2[1]), 
        .QN(n1060) );
  DFFTRX1 counter2_reg_3_ ( .D(N2174), .RN(n584), .CK(clk), .Q(counter2[3]), 
        .QN(n1059) );
  DFFTRX1 counter2_reg_0_ ( .D(N2171), .RN(n584), .CK(clk), .Q(counter2[0]), 
        .QN(n1061) );
  DFFTRX1 R15_reg_25_ ( .D(R14[25]), .RN(n579), .CK(clk), .Q(R15[25]) );
  DFFTRX1 R15_reg_24_ ( .D(R14[24]), .RN(n578), .CK(clk), .Q(R15[24]) );
  DFFTRX1 R15_reg_23_ ( .D(R14[23]), .RN(n576), .CK(clk), .Q(R15[23]) );
  DFFTRX1 R15_reg_22_ ( .D(R14[22]), .RN(n575), .CK(clk), .Q(R15[22]) );
  DFFTRX1 R6_reg_25_ ( .D(R5[25]), .RN(n580), .CK(clk), .Q(R6[25]) );
  DFFTRX1 R6_reg_24_ ( .D(R5[24]), .RN(n578), .CK(clk), .Q(R6[24]) );
  DFFTRX1 R6_reg_23_ ( .D(R5[23]), .RN(n577), .CK(clk), .Q(R6[23]) );
  DFFTRX1 R6_reg_22_ ( .D(R5[22]), .RN(n576), .CK(clk), .Q(R6[22]) );
  DFFTRX1 R6_reg_21_ ( .D(R5[21]), .RN(n575), .CK(clk), .Q(R6[21]) );
  DFFHQXL Wt_reg_31_ ( .D(N2164), .CK(clk), .Q(Wt[31]) );
  DFFTRX1 counter2_reg_2_ ( .D(N2173), .RN(n583), .CK(clk), .Q(counter2[2]) );
  DFFTRX1 R15_reg_21_ ( .D(R14[21]), .RN(n574), .CK(clk), .Q(R15[21]) );
  DFFTRX1 R15_reg_20_ ( .D(R14[20]), .RN(n573), .CK(clk), .Q(R15[20]) );
  DFFTRX1 R15_reg_19_ ( .D(R14[19]), .RN(n571), .CK(clk), .Q(R15[19]) );
  DFFTRX1 R15_reg_18_ ( .D(R14[18]), .RN(n570), .CK(clk), .Q(R15[18]) );
  DFFTRX1 counter1_reg_2_ ( .D(N1464), .RN(n2085), .CK(clk), .Q(counter1[2]), 
        .QN(n1057) );
  DFFTRX1 R6_reg_20_ ( .D(R5[20]), .RN(n573), .CK(clk), .Q(R6[20]) );
  DFFTRX1 R6_reg_19_ ( .D(R5[19]), .RN(n572), .CK(clk), .Q(R6[19]) );
  DFFTRX1 R6_reg_18_ ( .D(R5[18]), .RN(n571), .CK(clk), .Q(R6[18]) );
  DFFTRX1 R14_reg_2_ ( .D(R13[2]), .RN(n551), .CK(clk), .Q(R14[2]) );
  DFFTRX1 R1_reg_9_ ( .D(Wt[9]), .RN(n560), .CK(clk), .Q(R1[9]) );
  DFFTRX1 R1_reg_6_ ( .D(Wt[6]), .RN(n556), .CK(clk), .Q(R1[6]) );
  DFFTRX1 R1_reg_5_ ( .D(Wt[5]), .RN(n555), .CK(clk), .Q(R1[5]) );
  DFFTRX1 R1_reg_8_ ( .D(Wt[8]), .RN(n559), .CK(clk), .Q(R1[8]) );
  DFFTRX1 R1_reg_7_ ( .D(Wt[7]), .RN(n558), .CK(clk), .Q(R1[7]) );
  DFFHQXL Wt_reg_30_ ( .D(N2163), .CK(clk), .Q(Wt[30]) );
  DFFHQX1 Wt_reg_29_ ( .D(N2162), .CK(clk), .Q(Wt[29]) );
  DFFTRX1 counter1_reg_5_ ( .D(N1467), .RN(n2085), .CK(clk), .Q(counter1[5]), 
        .QN(n1056) );
  DFFTRX1 counter1_reg_3_ ( .D(N1465), .RN(n2085), .CK(clk), .Q(counter1[3])
         );
  DFFTRX1 counter1_reg_4_ ( .D(N1466), .RN(n2085), .CK(clk), .Q(counter1[4])
         );
  DFFTRX1 R15_reg_16_ ( .D(R14[16]), .RN(n568), .CK(clk), .Q(R15[16]) );
  DFFTRX1 R15_reg_15_ ( .D(R14[15]), .RN(n566), .CK(clk), .Q(R15[15]) );
  DFFTRX1 R15_reg_14_ ( .D(R14[14]), .RN(n565), .CK(clk), .Q(R15[14]) );
  DFFTRX1 R15_reg_17_ ( .D(R14[17]), .RN(n550), .CK(clk), .Q(R15[17]) );
  DFFTRX1 R6_reg_17_ ( .D(R5[17]), .RN(n570), .CK(clk), .Q(R6[17]) );
  DFFTRX1 R6_reg_16_ ( .D(R5[16]), .RN(n568), .CK(clk), .Q(R6[16]) );
  DFFTRX1 R6_reg_15_ ( .D(R5[15]), .RN(n567), .CK(clk), .Q(R6[15]) );
  DFFTRX1 R6_reg_14_ ( .D(R5[14]), .RN(n566), .CK(clk), .Q(R6[14]) );
  DFFTRX1 R14_reg_1_ ( .D(R13[1]), .RN(n547), .CK(clk), .Q(R14[1]) );
  DFFTRX1 R14_reg_0_ ( .D(R13[0]), .RN(n550), .CK(clk), .Q(R14[0]) );
  DFFTRX1 R1_reg_4_ ( .D(Wt[4]), .RN(n554), .CK(clk), .Q(R1[4]) );
  DFFHQX1 Wt_reg_28_ ( .D(N2161), .CK(clk), .Q(Wt[28]) );
  DFFTRX1 R1_reg_29_ ( .D(Wt[29]), .RN(n584), .CK(clk), .Q(R1[29]) );
  DFFTRX1 R1_reg_27_ ( .D(Wt[27]), .RN(n581), .CK(clk), .Q(R1[27]) );
  DFFTRX1 R14_reg_26_ ( .D(R13[26]), .RN(n580), .CK(clk), .Q(R14[26]) );
  DFFTRX1 R1_reg_31_ ( .D(Wt[31]), .RN(n585), .CK(clk), .Q(R1[31]) );
  DFFTRX1 R1_reg_30_ ( .D(Wt[30]), .RN(n547), .CK(clk), .Q(R1[30]) );
  DFFTRX1 R14_reg_28_ ( .D(R13[28]), .RN(n582), .CK(clk), .Q(R14[28]) );
  DFFTRX1 R14_reg_15_ ( .D(R13[15]), .RN(n566), .CK(clk), .Q(R14[15]) );
  DFFTRX1 R14_reg_17_ ( .D(R13[17]), .RN(n569), .CK(clk), .Q(R14[17]) );
  DFFTRX1 R14_reg_31_ ( .D(R13[31]), .RN(n584), .CK(clk), .Q(R14[31]) );
  DFFTRX1 R14_reg_30_ ( .D(R13[30]), .RN(n584), .CK(clk), .Q(R14[30]) );
  DFFTRX1 R14_reg_29_ ( .D(R13[29]), .RN(n583), .CK(clk), .Q(R14[29]) );
  DFFTRX1 R1_reg_0_ ( .D(Wt[0]), .RN(n585), .CK(clk), .Q(R1[0]) );
  DFFTRX1 R1_reg_3_ ( .D(Wt[3]), .RN(n553), .CK(clk), .Q(R1[3]) );
  DFFTRX1 R1_reg_2_ ( .D(Wt[2]), .RN(n551), .CK(clk), .Q(R1[2]) );
  DFFTRX1 R15_reg_13_ ( .D(R14[13]), .RN(n564), .CK(clk), .Q(R15[13]) );
  DFFTRX1 R15_reg_12_ ( .D(R14[12]), .RN(n563), .CK(clk), .Q(R15[12]) );
  DFFTRX1 R15_reg_11_ ( .D(R14[11]), .RN(n561), .CK(clk), .Q(R15[11]) );
  DFFTRX1 R15_reg_10_ ( .D(R14[10]), .RN(n560), .CK(clk), .Q(R15[10]) );
  DFFTRX1 R6_reg_13_ ( .D(R5[13]), .RN(n565), .CK(clk), .Q(R6[13]) );
  DFFTRX1 R6_reg_12_ ( .D(R5[12]), .RN(n563), .CK(clk), .Q(R6[12]) );
  DFFTRX1 R6_reg_11_ ( .D(R5[11]), .RN(n562), .CK(clk), .Q(R6[11]) );
  DFFTRX1 R6_reg_10_ ( .D(R5[10]), .RN(n561), .CK(clk), .Q(R6[10]) );
  DFFTRX1 R14_reg_21_ ( .D(R13[21]), .RN(n574), .CK(clk), .Q(R14[21]) );
  DFFTRX1 R14_reg_20_ ( .D(R13[20]), .RN(n573), .CK(clk), .Q(R14[20]) );
  DFFTRX1 R14_reg_19_ ( .D(R13[19]), .RN(n571), .CK(clk), .Q(R14[19]) );
  DFFTRX1 R14_reg_18_ ( .D(R13[18]), .RN(n570), .CK(clk), .Q(R14[18]) );
  DFFHQX1 Wt_reg_24_ ( .D(N2157), .CK(clk), .Q(Wt[24]) );
  DFFHQX1 Wt_reg_23_ ( .D(N2156), .CK(clk), .Q(Wt[23]) );
  DFFTRX1 R1_reg_20_ ( .D(Wt[20]), .RN(n574), .CK(clk), .Q(R1[20]) );
  DFFTRX1 R1_reg_19_ ( .D(Wt[19]), .RN(n572), .CK(clk), .Q(R1[19]) );
  DFFTRX1 R14_reg_3_ ( .D(R13[3]), .RN(n552), .CK(clk), .Q(R14[3]) );
  DFFTRX1 R14_reg_6_ ( .D(R13[6]), .RN(n555), .CK(clk), .Q(R14[6]) );
  DFFTRX1 R14_reg_5_ ( .D(R13[5]), .RN(n554), .CK(clk), .Q(R14[5]) );
  DFFTRX1 R14_reg_4_ ( .D(R13[4]), .RN(n553), .CK(clk), .Q(R14[4]) );
  DFFTRX1 R1_reg_28_ ( .D(Wt[28]), .RN(n583), .CK(clk), .Q(R1[28]) );
  DFFTRX1 R14_reg_27_ ( .D(R13[27]), .RN(n581), .CK(clk), .Q(R14[27]) );
  DFFTRX1 R1_reg_26_ ( .D(Wt[26]), .RN(n580), .CK(clk), .Q(R1[26]) );
  DFFTRX1 R1_reg_25_ ( .D(Wt[25]), .RN(n580), .CK(clk), .Q(R1[25]) );
  DFFTRX1 R14_reg_25_ ( .D(R13[25]), .RN(n579), .CK(clk), .Q(R14[25]) );
  DFFTRX1 R1_reg_24_ ( .D(Wt[24]), .RN(n579), .CK(clk), .Q(R1[24]) );
  DFFTRX1 R14_reg_24_ ( .D(R13[24]), .RN(n578), .CK(clk), .Q(R14[24]) );
  DFFTRX1 R14_reg_14_ ( .D(R13[14]), .RN(n565), .CK(clk), .Q(R14[14]) );
  DFFTRX1 R14_reg_13_ ( .D(R13[13]), .RN(n564), .CK(clk), .Q(R14[13]) );
  DFFTRX1 R14_reg_11_ ( .D(R13[11]), .RN(n561), .CK(clk), .Q(R14[11]) );
  DFFTRX1 R1_reg_16_ ( .D(Wt[16]), .RN(n569), .CK(clk), .Q(R1[16]) );
  DFFTRX1 R1_reg_15_ ( .D(Wt[15]), .RN(n568), .CK(clk), .Q(R1[15]) );
  DFFTRX1 R1_reg_14_ ( .D(Wt[14]), .RN(n566), .CK(clk), .Q(R1[14]) );
  DFFTRX1 R1_reg_13_ ( .D(Wt[13]), .RN(n565), .CK(clk), .Q(R1[13]) );
  DFFTRX1 R1_reg_12_ ( .D(Wt[12]), .RN(n564), .CK(clk), .Q(R1[12]) );
  DFFTRX1 R1_reg_11_ ( .D(Wt[11]), .RN(n563), .CK(clk), .Q(R1[11]) );
  DFFTRX1 R1_reg_10_ ( .D(Wt[10]), .RN(n561), .CK(clk), .Q(R1[10]) );
  DFFTRX1 R14_reg_10_ ( .D(R13[10]), .RN(n560), .CK(clk), .Q(R14[10]) );
  DFFTRX1 R14_reg_9_ ( .D(R13[9]), .RN(n559), .CK(clk), .Q(R14[9]) );
  DFFTRX1 R14_reg_8_ ( .D(R13[8]), .RN(n558), .CK(clk), .Q(R14[8]) );
  DFFTRX1 R14_reg_7_ ( .D(R13[7]), .RN(n556), .CK(clk), .Q(R14[7]) );
  DFFTRX1 R1_reg_17_ ( .D(Wt[17]), .RN(n570), .CK(clk), .Q(R1[17]) );
  DFFTRX1 R14_reg_16_ ( .D(R13[16]), .RN(n568), .CK(clk), .Q(R14[16]) );
  DFFTRX1 R15_reg_9_ ( .D(R14[9]), .RN(n559), .CK(clk), .Q(R15[9]) );
  DFFTRX1 R15_reg_8_ ( .D(R14[8]), .RN(n558), .CK(clk), .Q(R15[8]) );
  DFFTRX1 R15_reg_7_ ( .D(R14[7]), .RN(n556), .CK(clk), .Q(R15[7]) );
  DFFTRX1 R15_reg_6_ ( .D(R14[6]), .RN(n555), .CK(clk), .Q(R15[6]) );
  DFFTRX1 R6_reg_9_ ( .D(R5[9]), .RN(n560), .CK(clk), .Q(R6[9]) );
  DFFTRX1 R6_reg_8_ ( .D(R5[8]), .RN(n558), .CK(clk), .Q(R6[8]) );
  DFFTRX1 R6_reg_7_ ( .D(R5[7]), .RN(n557), .CK(clk), .Q(R6[7]) );
  DFFTRX1 R6_reg_6_ ( .D(R5[6]), .RN(n556), .CK(clk), .Q(R6[6]) );
  DFFHQX1 Wt_reg_22_ ( .D(N2155), .CK(clk), .Q(Wt[22]) );
  DFFHQX1 Wt_reg_20_ ( .D(N2153), .CK(clk), .Q(Wt[20]) );
  DFFTRX1 R15_reg_5_ ( .D(R14[5]), .RN(n554), .CK(clk), .Q(R15[5]) );
  DFFTRX1 R15_reg_4_ ( .D(R14[4]), .RN(n553), .CK(clk), .Q(R15[4]) );
  DFFTRX1 R15_reg_3_ ( .D(R14[3]), .RN(n550), .CK(clk), .Q(R15[3]) );
  DFFTRX1 R6_reg_5_ ( .D(R5[5]), .RN(n555), .CK(clk), .Q(R6[5]) );
  DFFTRX1 R6_reg_4_ ( .D(R5[4]), .RN(n553), .CK(clk), .Q(R6[4]) );
  DFFTRX1 R6_reg_3_ ( .D(R5[3]), .RN(n552), .CK(clk), .Q(R6[3]) );
  DFFHQX1 Wt_reg_19_ ( .D(N2152), .CK(clk), .Q(Wt[19]) );
  DFFHQX1 Wt_reg_16_ ( .D(N2149), .CK(clk), .Q(Wt[16]) );
  DFFTRX1 R2_reg_31_ ( .D(R1[31]), .RN(n585), .CK(clk), .Q(R2[31]) );
  DFFTRX1 R3_reg_31_ ( .D(R2[31]), .RN(n585), .CK(clk), .Q(R3[31]) );
  DFFTRX1 R4_reg_31_ ( .D(R3[31]), .RN(n585), .CK(clk), .Q(R4[31]) );
  DFFTRX1 R5_reg_31_ ( .D(R4[31]), .RN(n585), .CK(clk), .Q(R5[31]) );
  DFFTRX1 R7_reg_31_ ( .D(R6[31]), .RN(n585), .CK(clk), .Q(R7[31]) );
  DFFTRX1 R8_reg_31_ ( .D(R7[31]), .RN(n585), .CK(clk), .Q(R8[31]) );
  DFFTRX1 R9_reg_31_ ( .D(R8[31]), .RN(n585), .CK(clk), .Q(R9[31]) );
  DFFTRX1 R10_reg_31_ ( .D(R9[31]), .RN(n585), .CK(clk), .Q(R10[31]) );
  DFFTRX1 R11_reg_31_ ( .D(R10[31]), .RN(n585), .CK(clk), .Q(R11[31]) );
  DFFTRX1 R12_reg_31_ ( .D(R11[31]), .RN(n585), .CK(clk), .Q(R12[31]) );
  DFFTRX1 R13_reg_31_ ( .D(R12[31]), .RN(n585), .CK(clk), .Q(R13[31]) );
  DFFTRX1 R2_reg_30_ ( .D(R1[30]), .RN(n545), .CK(clk), .Q(R2[30]) );
  DFFTRX1 R3_reg_30_ ( .D(R2[30]), .RN(n585), .CK(clk), .Q(R3[30]) );
  DFFTRX1 R4_reg_30_ ( .D(R3[30]), .RN(n584), .CK(clk), .Q(R4[30]) );
  DFFTRX1 R5_reg_30_ ( .D(R4[30]), .RN(n581), .CK(clk), .Q(R5[30]) );
  DFFTRX1 R7_reg_30_ ( .D(R6[30]), .RN(n551), .CK(clk), .Q(R7[30]) );
  DFFTRX1 R8_reg_30_ ( .D(R7[30]), .RN(n552), .CK(clk), .Q(R8[30]) );
  DFFTRX1 R9_reg_30_ ( .D(R8[30]), .RN(n552), .CK(clk), .Q(R9[30]) );
  DFFTRX1 R10_reg_30_ ( .D(R9[30]), .RN(n584), .CK(clk), .Q(R10[30]) );
  DFFTRX1 R11_reg_30_ ( .D(R10[30]), .RN(n584), .CK(clk), .Q(R11[30]) );
  DFFTRX1 R12_reg_30_ ( .D(R11[30]), .RN(n584), .CK(clk), .Q(R12[30]) );
  DFFTRX1 R13_reg_30_ ( .D(R12[30]), .RN(n584), .CK(clk), .Q(R13[30]) );
  DFFTRX1 R2_reg_29_ ( .D(R1[29]), .RN(n584), .CK(clk), .Q(R2[29]) );
  DFFTRX1 R3_reg_29_ ( .D(R2[29]), .RN(n584), .CK(clk), .Q(R3[29]) );
  DFFTRX1 R4_reg_29_ ( .D(R3[29]), .RN(n584), .CK(clk), .Q(R4[29]) );
  DFFTRX1 R5_reg_29_ ( .D(R4[29]), .RN(n584), .CK(clk), .Q(R5[29]) );
  DFFTRX1 R7_reg_29_ ( .D(R6[29]), .RN(n583), .CK(clk), .Q(R7[29]) );
  DFFTRX1 R8_reg_29_ ( .D(R7[29]), .RN(n583), .CK(clk), .Q(R8[29]) );
  DFFTRX1 R9_reg_29_ ( .D(R8[29]), .RN(n583), .CK(clk), .Q(R9[29]) );
  DFFTRX1 R10_reg_29_ ( .D(R9[29]), .RN(n583), .CK(clk), .Q(R10[29]) );
  DFFTRX1 R11_reg_29_ ( .D(R10[29]), .RN(n583), .CK(clk), .Q(R11[29]) );
  DFFTRX1 R12_reg_29_ ( .D(R11[29]), .RN(n583), .CK(clk), .Q(R12[29]) );
  DFFTRX1 R13_reg_29_ ( .D(R12[29]), .RN(n583), .CK(clk), .Q(R13[29]) );
  DFFTRX1 R2_reg_28_ ( .D(R1[28]), .RN(n583), .CK(clk), .Q(R2[28]) );
  DFFTRX1 R3_reg_28_ ( .D(R2[28]), .RN(n583), .CK(clk), .Q(R3[28]) );
  DFFTRX1 R4_reg_28_ ( .D(R3[28]), .RN(n582), .CK(clk), .Q(R4[28]) );
  DFFTRX1 R5_reg_28_ ( .D(R4[28]), .RN(n582), .CK(clk), .Q(R5[28]) );
  DFFTRX1 R7_reg_28_ ( .D(R6[28]), .RN(n582), .CK(clk), .Q(R7[28]) );
  DFFTRX1 R8_reg_28_ ( .D(R7[28]), .RN(n582), .CK(clk), .Q(R8[28]) );
  DFFTRX1 R9_reg_28_ ( .D(R8[28]), .RN(n582), .CK(clk), .Q(R9[28]) );
  DFFTRX1 R10_reg_28_ ( .D(R9[28]), .RN(n582), .CK(clk), .Q(R10[28]) );
  DFFTRX1 R11_reg_28_ ( .D(R10[28]), .RN(n582), .CK(clk), .Q(R11[28]) );
  DFFTRX1 R12_reg_28_ ( .D(R11[28]), .RN(n582), .CK(clk), .Q(R12[28]) );
  DFFTRX1 R13_reg_28_ ( .D(R12[28]), .RN(n582), .CK(clk), .Q(R13[28]) );
  DFFTRX1 R8_reg_0_ ( .D(R7[0]), .RN(n550), .CK(clk), .Q(R8[0]) );
  DFFTRX1 R9_reg_0_ ( .D(R8[0]), .RN(n550), .CK(clk), .Q(R9[0]) );
  DFFTRX1 R10_reg_0_ ( .D(R9[0]), .RN(n550), .CK(clk), .Q(R10[0]) );
  DFFTRX1 R11_reg_0_ ( .D(R10[0]), .RN(n550), .CK(clk), .Q(R11[0]) );
  DFFTRX1 R12_reg_0_ ( .D(R11[0]), .RN(n550), .CK(clk), .Q(R12[0]) );
  DFFTRX1 R13_reg_0_ ( .D(R12[0]), .RN(n550), .CK(clk), .Q(R13[0]) );
  DFFTRX1 R2_reg_27_ ( .D(R1[27]), .RN(n581), .CK(clk), .Q(R2[27]) );
  DFFTRX1 R3_reg_27_ ( .D(R2[27]), .RN(n581), .CK(clk), .Q(R3[27]) );
  DFFTRX1 R4_reg_27_ ( .D(R3[27]), .RN(n581), .CK(clk), .Q(R4[27]) );
  DFFTRX1 R5_reg_27_ ( .D(R4[27]), .RN(n581), .CK(clk), .Q(R5[27]) );
  DFFTRX1 R7_reg_27_ ( .D(R6[27]), .RN(n581), .CK(clk), .Q(R7[27]) );
  DFFTRX1 R8_reg_27_ ( .D(R7[27]), .RN(n581), .CK(clk), .Q(R8[27]) );
  DFFTRX1 R9_reg_27_ ( .D(R8[27]), .RN(n581), .CK(clk), .Q(R9[27]) );
  DFFTRX1 R10_reg_27_ ( .D(R9[27]), .RN(n581), .CK(clk), .Q(R10[27]) );
  DFFTRX1 R11_reg_27_ ( .D(R10[27]), .RN(n581), .CK(clk), .Q(R11[27]) );
  DFFTRX1 R12_reg_27_ ( .D(R11[27]), .RN(n581), .CK(clk), .Q(R12[27]) );
  DFFTRX1 R13_reg_27_ ( .D(R12[27]), .RN(n585), .CK(clk), .Q(R13[27]) );
  DFFTRX1 R2_reg_26_ ( .D(R1[26]), .RN(n584), .CK(clk), .Q(R2[26]) );
  DFFTRX1 R3_reg_26_ ( .D(R2[26]), .RN(n581), .CK(clk), .Q(R3[26]) );
  DFFTRX1 R4_reg_26_ ( .D(R3[26]), .RN(n580), .CK(clk), .Q(R4[26]) );
  DFFTRX1 R5_reg_26_ ( .D(R4[26]), .RN(n581), .CK(clk), .Q(R5[26]) );
  DFFTRX1 R7_reg_26_ ( .D(R6[26]), .RN(n580), .CK(clk), .Q(R7[26]) );
  DFFTRX1 R8_reg_26_ ( .D(R7[26]), .RN(n581), .CK(clk), .Q(R8[26]) );
  DFFTRX1 R9_reg_26_ ( .D(R8[26]), .RN(n580), .CK(clk), .Q(R9[26]) );
  DFFTRX1 R10_reg_26_ ( .D(R9[26]), .RN(n580), .CK(clk), .Q(R10[26]) );
  DFFTRX1 R11_reg_26_ ( .D(R10[26]), .RN(n580), .CK(clk), .Q(R11[26]) );
  DFFTRX1 R12_reg_26_ ( .D(R11[26]), .RN(n580), .CK(clk), .Q(R12[26]) );
  DFFTRX1 R13_reg_26_ ( .D(R12[26]), .RN(n580), .CK(clk), .Q(R13[26]) );
  DFFTRX1 R2_reg_25_ ( .D(R1[25]), .RN(n580), .CK(clk), .Q(R2[25]) );
  DFFTRX1 R3_reg_25_ ( .D(R2[25]), .RN(n580), .CK(clk), .Q(R3[25]) );
  DFFTRX1 R4_reg_25_ ( .D(R3[25]), .RN(n580), .CK(clk), .Q(R4[25]) );
  DFFTRX1 R5_reg_25_ ( .D(R4[25]), .RN(n580), .CK(clk), .Q(R5[25]) );
  DFFTRX1 R7_reg_25_ ( .D(R6[25]), .RN(n579), .CK(clk), .Q(R7[25]) );
  DFFTRX1 R8_reg_25_ ( .D(R7[25]), .RN(n579), .CK(clk), .Q(R8[25]) );
  DFFTRX1 R9_reg_25_ ( .D(R8[25]), .RN(n579), .CK(clk), .Q(R9[25]) );
  DFFTRX1 R10_reg_25_ ( .D(R9[25]), .RN(n579), .CK(clk), .Q(R10[25]) );
  DFFTRX1 R11_reg_25_ ( .D(R10[25]), .RN(n579), .CK(clk), .Q(R11[25]) );
  DFFTRX1 R12_reg_25_ ( .D(R11[25]), .RN(n579), .CK(clk), .Q(R12[25]) );
  DFFTRX1 R13_reg_25_ ( .D(R12[25]), .RN(n579), .CK(clk), .Q(R13[25]) );
  DFFTRX1 R2_reg_24_ ( .D(R1[24]), .RN(n579), .CK(clk), .Q(R2[24]) );
  DFFTRX1 R3_reg_24_ ( .D(R2[24]), .RN(n579), .CK(clk), .Q(R3[24]) );
  DFFTRX1 R4_reg_24_ ( .D(R3[24]), .RN(n578), .CK(clk), .Q(R4[24]) );
  DFFTRX1 R5_reg_24_ ( .D(R4[24]), .RN(n578), .CK(clk), .Q(R5[24]) );
  DFFTRX1 R7_reg_24_ ( .D(R6[24]), .RN(n578), .CK(clk), .Q(R7[24]) );
  DFFTRX1 R8_reg_24_ ( .D(R7[24]), .RN(n578), .CK(clk), .Q(R8[24]) );
  DFFTRX1 R9_reg_24_ ( .D(R8[24]), .RN(n578), .CK(clk), .Q(R9[24]) );
  DFFTRX1 R10_reg_24_ ( .D(R9[24]), .RN(n578), .CK(clk), .Q(R10[24]) );
  DFFTRX1 R11_reg_24_ ( .D(R10[24]), .RN(n578), .CK(clk), .Q(R11[24]) );
  DFFTRX1 R12_reg_24_ ( .D(R11[24]), .RN(n578), .CK(clk), .Q(R12[24]) );
  DFFTRX1 R13_reg_24_ ( .D(R12[24]), .RN(n578), .CK(clk), .Q(R13[24]) );
  DFFTRX1 R2_reg_23_ ( .D(R1[23]), .RN(n577), .CK(clk), .Q(R2[23]) );
  DFFTRX1 R3_reg_23_ ( .D(R2[23]), .RN(n577), .CK(clk), .Q(R3[23]) );
  DFFTRX1 R4_reg_23_ ( .D(R3[23]), .RN(n577), .CK(clk), .Q(R4[23]) );
  DFFTRX1 R5_reg_23_ ( .D(R4[23]), .RN(n577), .CK(clk), .Q(R5[23]) );
  DFFTRX1 R7_reg_23_ ( .D(R6[23]), .RN(n577), .CK(clk), .Q(R7[23]) );
  DFFTRX1 R8_reg_23_ ( .D(R7[23]), .RN(n577), .CK(clk), .Q(R8[23]) );
  DFFTRX1 R9_reg_23_ ( .D(R8[23]), .RN(n577), .CK(clk), .Q(R9[23]) );
  DFFTRX1 R10_reg_23_ ( .D(R9[23]), .RN(n577), .CK(clk), .Q(R10[23]) );
  DFFTRX1 R11_reg_23_ ( .D(R10[23]), .RN(n577), .CK(clk), .Q(R11[23]) );
  DFFTRX1 R12_reg_23_ ( .D(R11[23]), .RN(n577), .CK(clk), .Q(R12[23]) );
  DFFTRX1 R13_reg_23_ ( .D(R12[23]), .RN(n576), .CK(clk), .Q(R13[23]) );
  DFFTRX1 R2_reg_22_ ( .D(R1[22]), .RN(n576), .CK(clk), .Q(R2[22]) );
  DFFTRX1 R3_reg_22_ ( .D(R2[22]), .RN(n576), .CK(clk), .Q(R3[22]) );
  DFFTRX1 R4_reg_22_ ( .D(R3[22]), .RN(n576), .CK(clk), .Q(R4[22]) );
  DFFTRX1 R5_reg_22_ ( .D(R4[22]), .RN(n576), .CK(clk), .Q(R5[22]) );
  DFFTRX1 R7_reg_22_ ( .D(R6[22]), .RN(n576), .CK(clk), .Q(R7[22]) );
  DFFTRX1 R8_reg_22_ ( .D(R7[22]), .RN(n576), .CK(clk), .Q(R8[22]) );
  DFFTRX1 R9_reg_22_ ( .D(R8[22]), .RN(n576), .CK(clk), .Q(R9[22]) );
  DFFTRX1 R10_reg_22_ ( .D(R9[22]), .RN(n575), .CK(clk), .Q(R10[22]) );
  DFFTRX1 R11_reg_22_ ( .D(R10[22]), .RN(n575), .CK(clk), .Q(R11[22]) );
  DFFTRX1 R12_reg_22_ ( .D(R11[22]), .RN(n575), .CK(clk), .Q(R12[22]) );
  DFFTRX1 R13_reg_22_ ( .D(R12[22]), .RN(n575), .CK(clk), .Q(R13[22]) );
  DFFTRX1 R2_reg_21_ ( .D(R1[21]), .RN(n575), .CK(clk), .Q(R2[21]) );
  DFFTRX1 R3_reg_21_ ( .D(R2[21]), .RN(n575), .CK(clk), .Q(R3[21]) );
  DFFTRX1 R4_reg_21_ ( .D(R3[21]), .RN(n575), .CK(clk), .Q(R4[21]) );
  DFFTRX1 R5_reg_21_ ( .D(R4[21]), .RN(n575), .CK(clk), .Q(R5[21]) );
  DFFTRX1 R7_reg_21_ ( .D(R6[21]), .RN(n574), .CK(clk), .Q(R7[21]) );
  DFFTRX1 R8_reg_21_ ( .D(R7[21]), .RN(n574), .CK(clk), .Q(R8[21]) );
  DFFTRX1 R9_reg_21_ ( .D(R8[21]), .RN(n574), .CK(clk), .Q(R9[21]) );
  DFFTRX1 R10_reg_21_ ( .D(R9[21]), .RN(n574), .CK(clk), .Q(R10[21]) );
  DFFTRX1 R11_reg_21_ ( .D(R10[21]), .RN(n574), .CK(clk), .Q(R11[21]) );
  DFFTRX1 R12_reg_21_ ( .D(R11[21]), .RN(n574), .CK(clk), .Q(R12[21]) );
  DFFTRX1 R13_reg_21_ ( .D(R12[21]), .RN(n574), .CK(clk), .Q(R13[21]) );
  DFFTRX1 R2_reg_20_ ( .D(R1[20]), .RN(n574), .CK(clk), .Q(R2[20]) );
  DFFTRX1 R3_reg_20_ ( .D(R2[20]), .RN(n574), .CK(clk), .Q(R3[20]) );
  DFFTRX1 R4_reg_20_ ( .D(R3[20]), .RN(n573), .CK(clk), .Q(R4[20]) );
  DFFTRX1 R5_reg_20_ ( .D(R4[20]), .RN(n573), .CK(clk), .Q(R5[20]) );
  DFFTRX1 R7_reg_20_ ( .D(R6[20]), .RN(n573), .CK(clk), .Q(R7[20]) );
  DFFTRX1 R8_reg_20_ ( .D(R7[20]), .RN(n573), .CK(clk), .Q(R8[20]) );
  DFFTRX1 R9_reg_20_ ( .D(R8[20]), .RN(n573), .CK(clk), .Q(R9[20]) );
  DFFTRX1 R10_reg_20_ ( .D(R9[20]), .RN(n573), .CK(clk), .Q(R10[20]) );
  DFFTRX1 R11_reg_20_ ( .D(R10[20]), .RN(n573), .CK(clk), .Q(R11[20]) );
  DFFTRX1 R12_reg_20_ ( .D(R11[20]), .RN(n573), .CK(clk), .Q(R12[20]) );
  DFFTRX1 R13_reg_20_ ( .D(R12[20]), .RN(n573), .CK(clk), .Q(R13[20]) );
  DFFTRX1 R2_reg_19_ ( .D(R1[19]), .RN(n572), .CK(clk), .Q(R2[19]) );
  DFFTRX1 R3_reg_19_ ( .D(R2[19]), .RN(n572), .CK(clk), .Q(R3[19]) );
  DFFTRX1 R4_reg_19_ ( .D(R3[19]), .RN(n572), .CK(clk), .Q(R4[19]) );
  DFFTRX1 R5_reg_19_ ( .D(R4[19]), .RN(n572), .CK(clk), .Q(R5[19]) );
  DFFTRX1 R7_reg_19_ ( .D(R6[19]), .RN(n572), .CK(clk), .Q(R7[19]) );
  DFFTRX1 R8_reg_19_ ( .D(R7[19]), .RN(n572), .CK(clk), .Q(R8[19]) );
  DFFTRX1 R9_reg_19_ ( .D(R8[19]), .RN(n572), .CK(clk), .Q(R9[19]) );
  DFFTRX1 R10_reg_19_ ( .D(R9[19]), .RN(n572), .CK(clk), .Q(R10[19]) );
  DFFTRX1 R11_reg_19_ ( .D(R10[19]), .RN(n572), .CK(clk), .Q(R11[19]) );
  DFFTRX1 R12_reg_19_ ( .D(R11[19]), .RN(n572), .CK(clk), .Q(R12[19]) );
  DFFTRX1 R13_reg_19_ ( .D(R12[19]), .RN(n571), .CK(clk), .Q(R13[19]) );
  DFFTRX1 R2_reg_18_ ( .D(R1[18]), .RN(n571), .CK(clk), .Q(R2[18]) );
  DFFTRX1 R3_reg_18_ ( .D(R2[18]), .RN(n571), .CK(clk), .Q(R3[18]) );
  DFFTRX1 R4_reg_18_ ( .D(R3[18]), .RN(n571), .CK(clk), .Q(R4[18]) );
  DFFTRX1 R5_reg_18_ ( .D(R4[18]), .RN(n571), .CK(clk), .Q(R5[18]) );
  DFFTRX1 R7_reg_18_ ( .D(R6[18]), .RN(n571), .CK(clk), .Q(R7[18]) );
  DFFTRX1 R8_reg_18_ ( .D(R7[18]), .RN(n571), .CK(clk), .Q(R8[18]) );
  DFFTRX1 R9_reg_18_ ( .D(R8[18]), .RN(n571), .CK(clk), .Q(R9[18]) );
  DFFTRX1 R10_reg_18_ ( .D(R9[18]), .RN(n570), .CK(clk), .Q(R10[18]) );
  DFFTRX1 R11_reg_18_ ( .D(R10[18]), .RN(n570), .CK(clk), .Q(R11[18]) );
  DFFTRX1 R12_reg_18_ ( .D(R11[18]), .RN(n570), .CK(clk), .Q(R12[18]) );
  DFFTRX1 R13_reg_18_ ( .D(R12[18]), .RN(n570), .CK(clk), .Q(R13[18]) );
  DFFTRX1 R2_reg_17_ ( .D(R1[17]), .RN(n570), .CK(clk), .Q(R2[17]) );
  DFFTRX1 R3_reg_17_ ( .D(R2[17]), .RN(n570), .CK(clk), .Q(R3[17]) );
  DFFTRX1 R4_reg_17_ ( .D(R3[17]), .RN(n570), .CK(clk), .Q(R4[17]) );
  DFFTRX1 R5_reg_17_ ( .D(R4[17]), .RN(n570), .CK(clk), .Q(R5[17]) );
  DFFTRX1 R7_reg_17_ ( .D(R6[17]), .RN(n569), .CK(clk), .Q(R7[17]) );
  DFFTRX1 R8_reg_17_ ( .D(R7[17]), .RN(n569), .CK(clk), .Q(R8[17]) );
  DFFTRX1 R9_reg_17_ ( .D(R8[17]), .RN(n569), .CK(clk), .Q(R9[17]) );
  DFFTRX1 R10_reg_17_ ( .D(R9[17]), .RN(n569), .CK(clk), .Q(R10[17]) );
  DFFTRX1 R11_reg_17_ ( .D(R10[17]), .RN(n569), .CK(clk), .Q(R11[17]) );
  DFFTRX1 R12_reg_17_ ( .D(R11[17]), .RN(n569), .CK(clk), .Q(R12[17]) );
  DFFTRX1 R13_reg_17_ ( .D(R12[17]), .RN(n569), .CK(clk), .Q(R13[17]) );
  DFFTRX1 R2_reg_16_ ( .D(R1[16]), .RN(n569), .CK(clk), .Q(R2[16]) );
  DFFTRX1 R3_reg_16_ ( .D(R2[16]), .RN(n569), .CK(clk), .Q(R3[16]) );
  DFFTRX1 R4_reg_16_ ( .D(R3[16]), .RN(n569), .CK(clk), .Q(R4[16]) );
  DFFTRX1 R5_reg_16_ ( .D(R4[16]), .RN(n568), .CK(clk), .Q(R5[16]) );
  DFFTRX1 R7_reg_16_ ( .D(R6[16]), .RN(n568), .CK(clk), .Q(R7[16]) );
  DFFTRX1 R8_reg_16_ ( .D(R7[16]), .RN(n568), .CK(clk), .Q(R8[16]) );
  DFFTRX1 R9_reg_16_ ( .D(R8[16]), .RN(n568), .CK(clk), .Q(R9[16]) );
  DFFTRX1 R10_reg_16_ ( .D(R9[16]), .RN(n568), .CK(clk), .Q(R10[16]) );
  DFFTRX1 R11_reg_16_ ( .D(R10[16]), .RN(n568), .CK(clk), .Q(R11[16]) );
  DFFTRX1 R12_reg_16_ ( .D(R11[16]), .RN(n568), .CK(clk), .Q(R12[16]) );
  DFFTRX1 R13_reg_16_ ( .D(R12[16]), .RN(n568), .CK(clk), .Q(R13[16]) );
  DFFTRX1 R2_reg_15_ ( .D(R1[15]), .RN(n567), .CK(clk), .Q(R2[15]) );
  DFFTRX1 R3_reg_15_ ( .D(R2[15]), .RN(n567), .CK(clk), .Q(R3[15]) );
  DFFTRX1 R4_reg_15_ ( .D(R3[15]), .RN(n567), .CK(clk), .Q(R4[15]) );
  DFFTRX1 R5_reg_15_ ( .D(R4[15]), .RN(n567), .CK(clk), .Q(R5[15]) );
  DFFTRX1 R7_reg_15_ ( .D(R6[15]), .RN(n567), .CK(clk), .Q(R7[15]) );
  DFFTRX1 R8_reg_15_ ( .D(R7[15]), .RN(n567), .CK(clk), .Q(R8[15]) );
  DFFTRX1 R9_reg_15_ ( .D(R8[15]), .RN(n567), .CK(clk), .Q(R9[15]) );
  DFFTRX1 R10_reg_15_ ( .D(R9[15]), .RN(n567), .CK(clk), .Q(R10[15]) );
  DFFTRX1 R11_reg_15_ ( .D(R10[15]), .RN(n567), .CK(clk), .Q(R11[15]) );
  DFFTRX1 R12_reg_15_ ( .D(R11[15]), .RN(n567), .CK(clk), .Q(R12[15]) );
  DFFTRX1 R13_reg_15_ ( .D(R12[15]), .RN(n567), .CK(clk), .Q(R13[15]) );
  DFFTRX1 R2_reg_14_ ( .D(R1[14]), .RN(n566), .CK(clk), .Q(R2[14]) );
  DFFTRX1 R3_reg_14_ ( .D(R2[14]), .RN(n566), .CK(clk), .Q(R3[14]) );
  DFFTRX1 R4_reg_14_ ( .D(R3[14]), .RN(n566), .CK(clk), .Q(R4[14]) );
  DFFTRX1 R5_reg_14_ ( .D(R4[14]), .RN(n566), .CK(clk), .Q(R5[14]) );
  DFFTRX1 R7_reg_14_ ( .D(R6[14]), .RN(n566), .CK(clk), .Q(R7[14]) );
  DFFTRX1 R8_reg_14_ ( .D(R7[14]), .RN(n566), .CK(clk), .Q(R8[14]) );
  DFFTRX1 R9_reg_14_ ( .D(R8[14]), .RN(n566), .CK(clk), .Q(R9[14]) );
  DFFTRX1 R10_reg_14_ ( .D(R9[14]), .RN(n566), .CK(clk), .Q(R10[14]) );
  DFFTRX1 R11_reg_14_ ( .D(R10[14]), .RN(n565), .CK(clk), .Q(R11[14]) );
  DFFTRX1 R12_reg_14_ ( .D(R11[14]), .RN(n565), .CK(clk), .Q(R12[14]) );
  DFFTRX1 R13_reg_14_ ( .D(R12[14]), .RN(n565), .CK(clk), .Q(R13[14]) );
  DFFTRX1 R2_reg_13_ ( .D(R1[13]), .RN(n565), .CK(clk), .Q(R2[13]) );
  DFFTRX1 R3_reg_13_ ( .D(R2[13]), .RN(n565), .CK(clk), .Q(R3[13]) );
  DFFTRX1 R4_reg_13_ ( .D(R3[13]), .RN(n565), .CK(clk), .Q(R4[13]) );
  DFFTRX1 R5_reg_13_ ( .D(R4[13]), .RN(n565), .CK(clk), .Q(R5[13]) );
  DFFTRX1 R7_reg_13_ ( .D(R6[13]), .RN(n565), .CK(clk), .Q(R7[13]) );
  DFFTRX1 R8_reg_13_ ( .D(R7[13]), .RN(n564), .CK(clk), .Q(R8[13]) );
  DFFTRX1 R9_reg_13_ ( .D(R8[13]), .RN(n564), .CK(clk), .Q(R9[13]) );
  DFFTRX1 R10_reg_13_ ( .D(R9[13]), .RN(n564), .CK(clk), .Q(R10[13]) );
  DFFTRX1 R11_reg_13_ ( .D(R10[13]), .RN(n564), .CK(clk), .Q(R11[13]) );
  DFFTRX1 R12_reg_13_ ( .D(R11[13]), .RN(n564), .CK(clk), .Q(R12[13]) );
  DFFTRX1 R13_reg_13_ ( .D(R12[13]), .RN(n564), .CK(clk), .Q(R13[13]) );
  DFFTRX1 R2_reg_12_ ( .D(R1[12]), .RN(n564), .CK(clk), .Q(R2[12]) );
  DFFTRX1 R3_reg_12_ ( .D(R2[12]), .RN(n564), .CK(clk), .Q(R3[12]) );
  DFFTRX1 R4_reg_12_ ( .D(R3[12]), .RN(n564), .CK(clk), .Q(R4[12]) );
  DFFTRX1 R5_reg_12_ ( .D(R4[12]), .RN(n563), .CK(clk), .Q(R5[12]) );
  DFFTRX1 R7_reg_12_ ( .D(R6[12]), .RN(n563), .CK(clk), .Q(R7[12]) );
  DFFTRX1 R8_reg_12_ ( .D(R7[12]), .RN(n563), .CK(clk), .Q(R8[12]) );
  DFFTRX1 R9_reg_12_ ( .D(R8[12]), .RN(n563), .CK(clk), .Q(R9[12]) );
  DFFTRX1 R10_reg_12_ ( .D(R9[12]), .RN(n563), .CK(clk), .Q(R10[12]) );
  DFFTRX1 R11_reg_12_ ( .D(R10[12]), .RN(n563), .CK(clk), .Q(R11[12]) );
  DFFTRX1 R12_reg_12_ ( .D(R11[12]), .RN(n563), .CK(clk), .Q(R12[12]) );
  DFFTRX1 R13_reg_12_ ( .D(R12[12]), .RN(n563), .CK(clk), .Q(R13[12]) );
  DFFTRX1 R2_reg_11_ ( .D(R1[11]), .RN(n562), .CK(clk), .Q(R2[11]) );
  DFFTRX1 R3_reg_11_ ( .D(R2[11]), .RN(n562), .CK(clk), .Q(R3[11]) );
  DFFTRX1 R4_reg_11_ ( .D(R3[11]), .RN(n562), .CK(clk), .Q(R4[11]) );
  DFFTRX1 R5_reg_11_ ( .D(R4[11]), .RN(n562), .CK(clk), .Q(R5[11]) );
  DFFTRX1 R7_reg_11_ ( .D(R6[11]), .RN(n562), .CK(clk), .Q(R7[11]) );
  DFFTRX1 R8_reg_11_ ( .D(R7[11]), .RN(n562), .CK(clk), .Q(R8[11]) );
  DFFTRX1 R9_reg_11_ ( .D(R8[11]), .RN(n562), .CK(clk), .Q(R9[11]) );
  DFFTRX1 R10_reg_11_ ( .D(R9[11]), .RN(n562), .CK(clk), .Q(R10[11]) );
  DFFTRX1 R11_reg_11_ ( .D(R10[11]), .RN(n562), .CK(clk), .Q(R11[11]) );
  DFFTRX1 R12_reg_11_ ( .D(R11[11]), .RN(n562), .CK(clk), .Q(R12[11]) );
  DFFTRX1 R13_reg_11_ ( .D(R12[11]), .RN(n562), .CK(clk), .Q(R13[11]) );
  DFFTRX1 R2_reg_10_ ( .D(R1[10]), .RN(n561), .CK(clk), .Q(R2[10]) );
  DFFTRX1 R3_reg_10_ ( .D(R2[10]), .RN(n561), .CK(clk), .Q(R3[10]) );
  DFFTRX1 R4_reg_10_ ( .D(R3[10]), .RN(n561), .CK(clk), .Q(R4[10]) );
  DFFTRX1 R5_reg_10_ ( .D(R4[10]), .RN(n561), .CK(clk), .Q(R5[10]) );
  DFFTRX1 R7_reg_10_ ( .D(R6[10]), .RN(n561), .CK(clk), .Q(R7[10]) );
  DFFTRX1 R8_reg_10_ ( .D(R7[10]), .RN(n561), .CK(clk), .Q(R8[10]) );
  DFFTRX1 R9_reg_10_ ( .D(R8[10]), .RN(n561), .CK(clk), .Q(R9[10]) );
  DFFTRX1 R10_reg_10_ ( .D(R9[10]), .RN(n561), .CK(clk), .Q(R10[10]) );
  DFFTRX1 R11_reg_10_ ( .D(R10[10]), .RN(n560), .CK(clk), .Q(R11[10]) );
  DFFTRX1 R12_reg_10_ ( .D(R11[10]), .RN(n560), .CK(clk), .Q(R12[10]) );
  DFFTRX1 R13_reg_10_ ( .D(R12[10]), .RN(n560), .CK(clk), .Q(R13[10]) );
  DFFTRX1 R2_reg_9_ ( .D(R1[9]), .RN(n560), .CK(clk), .Q(R2[9]) );
  DFFTRX1 R3_reg_9_ ( .D(R2[9]), .RN(n560), .CK(clk), .Q(R3[9]) );
  DFFTRX1 R4_reg_9_ ( .D(R3[9]), .RN(n560), .CK(clk), .Q(R4[9]) );
  DFFTRX1 R5_reg_9_ ( .D(R4[9]), .RN(n560), .CK(clk), .Q(R5[9]) );
  DFFTRX1 R7_reg_9_ ( .D(R6[9]), .RN(n560), .CK(clk), .Q(R7[9]) );
  DFFTRX1 R8_reg_9_ ( .D(R7[9]), .RN(n559), .CK(clk), .Q(R8[9]) );
  DFFTRX1 R9_reg_9_ ( .D(R8[9]), .RN(n559), .CK(clk), .Q(R9[9]) );
  DFFTRX1 R10_reg_9_ ( .D(R9[9]), .RN(n559), .CK(clk), .Q(R10[9]) );
  DFFTRX1 R11_reg_9_ ( .D(R10[9]), .RN(n559), .CK(clk), .Q(R11[9]) );
  DFFTRX1 R12_reg_9_ ( .D(R11[9]), .RN(n559), .CK(clk), .Q(R12[9]) );
  DFFTRX1 R13_reg_9_ ( .D(R12[9]), .RN(n559), .CK(clk), .Q(R13[9]) );
  DFFTRX1 R2_reg_8_ ( .D(R1[8]), .RN(n559), .CK(clk), .Q(R2[8]) );
  DFFTRX1 R3_reg_8_ ( .D(R2[8]), .RN(n559), .CK(clk), .Q(R3[8]) );
  DFFTRX1 R4_reg_8_ ( .D(R3[8]), .RN(n559), .CK(clk), .Q(R4[8]) );
  DFFTRX1 R5_reg_8_ ( .D(R4[8]), .RN(n558), .CK(clk), .Q(R5[8]) );
  DFFTRX1 R7_reg_8_ ( .D(R6[8]), .RN(n558), .CK(clk), .Q(R7[8]) );
  DFFTRX1 R8_reg_8_ ( .D(R7[8]), .RN(n558), .CK(clk), .Q(R8[8]) );
  DFFTRX1 R9_reg_8_ ( .D(R8[8]), .RN(n558), .CK(clk), .Q(R9[8]) );
  DFFTRX1 R10_reg_8_ ( .D(R9[8]), .RN(n558), .CK(clk), .Q(R10[8]) );
  DFFTRX1 R11_reg_8_ ( .D(R10[8]), .RN(n558), .CK(clk), .Q(R11[8]) );
  DFFTRX1 R12_reg_8_ ( .D(R11[8]), .RN(n558), .CK(clk), .Q(R12[8]) );
  DFFTRX1 R13_reg_8_ ( .D(R12[8]), .RN(n558), .CK(clk), .Q(R13[8]) );
  DFFTRX1 R2_reg_7_ ( .D(R1[7]), .RN(n557), .CK(clk), .Q(R2[7]) );
  DFFTRX1 R3_reg_7_ ( .D(R2[7]), .RN(n557), .CK(clk), .Q(R3[7]) );
  DFFTRX1 R4_reg_7_ ( .D(R3[7]), .RN(n557), .CK(clk), .Q(R4[7]) );
  DFFTRX1 R5_reg_7_ ( .D(R4[7]), .RN(n557), .CK(clk), .Q(R5[7]) );
  DFFTRX1 R7_reg_7_ ( .D(R6[7]), .RN(n557), .CK(clk), .Q(R7[7]) );
  DFFTRX1 R8_reg_7_ ( .D(R7[7]), .RN(n557), .CK(clk), .Q(R8[7]) );
  DFFTRX1 R9_reg_7_ ( .D(R8[7]), .RN(n557), .CK(clk), .Q(R9[7]) );
  DFFTRX1 R10_reg_7_ ( .D(R9[7]), .RN(n557), .CK(clk), .Q(R10[7]) );
  DFFTRX1 R11_reg_7_ ( .D(R10[7]), .RN(n557), .CK(clk), .Q(R11[7]) );
  DFFTRX1 R12_reg_7_ ( .D(R11[7]), .RN(n557), .CK(clk), .Q(R12[7]) );
  DFFTRX1 R13_reg_7_ ( .D(R12[7]), .RN(n557), .CK(clk), .Q(R13[7]) );
  DFFTRX1 R2_reg_6_ ( .D(R1[6]), .RN(n556), .CK(clk), .Q(R2[6]) );
  DFFTRX1 R3_reg_6_ ( .D(R2[6]), .RN(n556), .CK(clk), .Q(R3[6]) );
  DFFTRX1 R4_reg_6_ ( .D(R3[6]), .RN(n556), .CK(clk), .Q(R4[6]) );
  DFFTRX1 R5_reg_6_ ( .D(R4[6]), .RN(n556), .CK(clk), .Q(R5[6]) );
  DFFTRX1 R7_reg_6_ ( .D(R6[6]), .RN(n556), .CK(clk), .Q(R7[6]) );
  DFFTRX1 R8_reg_6_ ( .D(R7[6]), .RN(n556), .CK(clk), .Q(R8[6]) );
  DFFTRX1 R9_reg_6_ ( .D(R8[6]), .RN(n556), .CK(clk), .Q(R9[6]) );
  DFFTRX1 R10_reg_6_ ( .D(R9[6]), .RN(n556), .CK(clk), .Q(R10[6]) );
  DFFTRX1 R11_reg_6_ ( .D(R10[6]), .RN(n555), .CK(clk), .Q(R11[6]) );
  DFFTRX1 R12_reg_6_ ( .D(R11[6]), .RN(n555), .CK(clk), .Q(R12[6]) );
  DFFTRX1 R13_reg_6_ ( .D(R12[6]), .RN(n555), .CK(clk), .Q(R13[6]) );
  DFFTRX1 R2_reg_5_ ( .D(R1[5]), .RN(n555), .CK(clk), .Q(R2[5]) );
  DFFTRX1 R3_reg_5_ ( .D(R2[5]), .RN(n555), .CK(clk), .Q(R3[5]) );
  DFFTRX1 R4_reg_5_ ( .D(R3[5]), .RN(n555), .CK(clk), .Q(R4[5]) );
  DFFTRX1 R5_reg_5_ ( .D(R4[5]), .RN(n555), .CK(clk), .Q(R5[5]) );
  DFFTRX1 R7_reg_5_ ( .D(R6[5]), .RN(n555), .CK(clk), .Q(R7[5]) );
  DFFTRX1 R8_reg_5_ ( .D(R7[5]), .RN(n554), .CK(clk), .Q(R8[5]) );
  DFFTRX1 R9_reg_5_ ( .D(R8[5]), .RN(n554), .CK(clk), .Q(R9[5]) );
  DFFTRX1 R10_reg_5_ ( .D(R9[5]), .RN(n554), .CK(clk), .Q(R10[5]) );
  DFFTRX1 R11_reg_5_ ( .D(R10[5]), .RN(n554), .CK(clk), .Q(R11[5]) );
  DFFTRX1 R12_reg_5_ ( .D(R11[5]), .RN(n554), .CK(clk), .Q(R12[5]) );
  DFFTRX1 R13_reg_5_ ( .D(R12[5]), .RN(n554), .CK(clk), .Q(R13[5]) );
  DFFTRX1 R2_reg_4_ ( .D(R1[4]), .RN(n554), .CK(clk), .Q(R2[4]) );
  DFFTRX1 R3_reg_4_ ( .D(R2[4]), .RN(n554), .CK(clk), .Q(R3[4]) );
  DFFTRX1 R4_reg_4_ ( .D(R3[4]), .RN(n554), .CK(clk), .Q(R4[4]) );
  DFFTRX1 R5_reg_4_ ( .D(R4[4]), .RN(n553), .CK(clk), .Q(R5[4]) );
  DFFTRX1 R7_reg_4_ ( .D(R6[4]), .RN(n553), .CK(clk), .Q(R7[4]) );
  DFFTRX1 R8_reg_4_ ( .D(R7[4]), .RN(n553), .CK(clk), .Q(R8[4]) );
  DFFTRX1 R9_reg_4_ ( .D(R8[4]), .RN(n553), .CK(clk), .Q(R9[4]) );
  DFFTRX1 R10_reg_4_ ( .D(R9[4]), .RN(n553), .CK(clk), .Q(R10[4]) );
  DFFTRX1 R11_reg_4_ ( .D(R10[4]), .RN(n553), .CK(clk), .Q(R11[4]) );
  DFFTRX1 R12_reg_4_ ( .D(R11[4]), .RN(n553), .CK(clk), .Q(R12[4]) );
  DFFTRX1 R13_reg_4_ ( .D(R12[4]), .RN(n553), .CK(clk), .Q(R13[4]) );
  DFFTRX1 R2_reg_3_ ( .D(R1[3]), .RN(n552), .CK(clk), .Q(R2[3]) );
  DFFTRX1 R3_reg_3_ ( .D(R2[3]), .RN(n552), .CK(clk), .Q(R3[3]) );
  DFFTRX1 R4_reg_3_ ( .D(R3[3]), .RN(n552), .CK(clk), .Q(R4[3]) );
  DFFTRX1 R5_reg_3_ ( .D(R4[3]), .RN(n552), .CK(clk), .Q(R5[3]) );
  DFFTRX1 R7_reg_3_ ( .D(R6[3]), .RN(n552), .CK(clk), .Q(R7[3]) );
  DFFTRX1 R8_reg_3_ ( .D(R7[3]), .RN(n552), .CK(clk), .Q(R8[3]) );
  DFFTRX1 R9_reg_3_ ( .D(R8[3]), .RN(n552), .CK(clk), .Q(R9[3]) );
  DFFTRX1 R10_reg_3_ ( .D(R9[3]), .RN(n552), .CK(clk), .Q(R10[3]) );
  DFFTRX1 R11_reg_3_ ( .D(R10[3]), .RN(n552), .CK(clk), .Q(R11[3]) );
  DFFTRX1 R12_reg_3_ ( .D(R11[3]), .RN(n552), .CK(clk), .Q(R12[3]) );
  DFFTRX1 R13_reg_3_ ( .D(R12[3]), .RN(n552), .CK(clk), .Q(R13[3]) );
  DFFTRX1 R2_reg_2_ ( .D(R1[2]), .RN(n551), .CK(clk), .Q(R2[2]) );
  DFFTRX1 R3_reg_2_ ( .D(R2[2]), .RN(n552), .CK(clk), .Q(R3[2]) );
  DFFTRX1 R4_reg_2_ ( .D(R3[2]), .RN(n550), .CK(clk), .Q(R4[2]) );
  DFFTRX1 R5_reg_2_ ( .D(R4[2]), .RN(n551), .CK(clk), .Q(R5[2]) );
  DFFTRX1 R7_reg_2_ ( .D(R6[2]), .RN(n552), .CK(clk), .Q(R7[2]) );
  DFFTRX1 R8_reg_2_ ( .D(R7[2]), .RN(n550), .CK(clk), .Q(R8[2]) );
  DFFTRX1 R9_reg_2_ ( .D(R8[2]), .RN(n551), .CK(clk), .Q(R9[2]) );
  DFFTRX1 R10_reg_2_ ( .D(R9[2]), .RN(n552), .CK(clk), .Q(R10[2]) );
  DFFTRX1 R11_reg_2_ ( .D(R10[2]), .RN(n551), .CK(clk), .Q(R11[2]) );
  DFFTRX1 R12_reg_2_ ( .D(R11[2]), .RN(n551), .CK(clk), .Q(R12[2]) );
  DFFTRX1 R13_reg_2_ ( .D(R12[2]), .RN(n551), .CK(clk), .Q(R13[2]) );
  DFFTRX1 R2_reg_1_ ( .D(R1[1]), .RN(n551), .CK(clk), .Q(R2[1]) );
  DFFTRX1 R3_reg_1_ ( .D(R2[1]), .RN(n551), .CK(clk), .Q(R3[1]) );
  DFFTRX1 R4_reg_1_ ( .D(R3[1]), .RN(n551), .CK(clk), .Q(R4[1]) );
  DFFTRX1 R5_reg_1_ ( .D(R4[1]), .RN(n551), .CK(clk), .Q(R5[1]) );
  DFFTRX1 R7_reg_1_ ( .D(R6[1]), .RN(n551), .CK(clk), .Q(R7[1]) );
  DFFTRX1 R8_reg_1_ ( .D(R7[1]), .RN(n584), .CK(clk), .Q(R8[1]) );
  DFFTRX1 R9_reg_1_ ( .D(R8[1]), .RN(n581), .CK(clk), .Q(R9[1]) );
  DFFTRX1 R10_reg_1_ ( .D(R9[1]), .RN(n580), .CK(clk), .Q(R10[1]) );
  DFFTRX1 R11_reg_1_ ( .D(R10[1]), .RN(n547), .CK(clk), .Q(R11[1]) );
  DFFTRX1 R12_reg_1_ ( .D(R11[1]), .RN(n550), .CK(clk), .Q(R12[1]) );
  DFFTRX1 R13_reg_1_ ( .D(R12[1]), .RN(n585), .CK(clk), .Q(R13[1]) );
  DFFTRX1 R2_reg_0_ ( .D(R1[0]), .RN(n584), .CK(clk), .Q(R2[0]) );
  DFFTRX1 R3_reg_0_ ( .D(R2[0]), .RN(n581), .CK(clk), .Q(R3[0]) );
  DFFTRX1 R4_reg_0_ ( .D(R3[0]), .RN(n580), .CK(clk), .Q(R4[0]) );
  DFFTRX1 R5_reg_0_ ( .D(R4[0]), .RN(n550), .CK(clk), .Q(R5[0]) );
  DFFHQXL Wt_reg_25_ ( .D(N2158), .CK(clk), .Q(Wt[25]) );
  DFFHQX1 Wt_reg_21_ ( .D(N2154), .CK(clk), .Q(Wt[21]) );
  DFFHQXL buffer_reg_0__27_ ( .D(n794), .CK(clk), .Q(buffer[123]) );
  DFFHQXL buffer_reg_0__28_ ( .D(n793), .CK(clk), .Q(buffer[124]) );
  DFFHQXL buffer_reg_0__29_ ( .D(n792), .CK(clk), .Q(buffer[125]) );
  DFFHQXL buffer_reg_0__30_ ( .D(n791), .CK(clk), .Q(buffer[126]) );
  DFFHQXL buffer_reg_0__31_ ( .D(n790), .CK(clk), .Q(buffer[127]) );
  DFFHQXL buffer_reg_2__24_ ( .D(n859), .CK(clk), .Q(buffer[104]) );
  DFFHQXL buffer_reg_2__25_ ( .D(n858), .CK(clk), .Q(buffer[105]) );
  DFFHQXL buffer_reg_2__26_ ( .D(n857), .CK(clk), .Q(buffer[106]) );
  DFFHQXL buffer_reg_2__27_ ( .D(n856), .CK(clk), .Q(buffer[107]) );
  DFFHQXL buffer_reg_2__28_ ( .D(n855), .CK(clk), .Q(buffer[108]) );
  DFFHQXL buffer_reg_2__29_ ( .D(n854), .CK(clk), .Q(buffer[109]) );
  DFFHQXL buffer_reg_2__30_ ( .D(n853), .CK(clk), .Q(buffer[110]) );
  DFFHQXL buffer_reg_2__31_ ( .D(n852), .CK(clk), .Q(buffer[111]) );
  DFFHQXL buffer_reg_4__24_ ( .D(n28), .CK(clk), .Q(buffer[88]) );
  DFFHQXL buffer_reg_4__25_ ( .D(n920), .CK(clk), .Q(buffer[89]) );
  DFFHQXL buffer_reg_4__26_ ( .D(n919), .CK(clk), .Q(buffer[90]) );
  DFFHQXL buffer_reg_4__27_ ( .D(n918), .CK(clk), .Q(buffer[91]) );
  DFFHQXL buffer_reg_4__28_ ( .D(n917), .CK(clk), .Q(buffer[92]) );
  DFFHQXL buffer_reg_4__29_ ( .D(n916), .CK(clk), .Q(buffer[93]) );
  DFFHQXL buffer_reg_4__30_ ( .D(n915), .CK(clk), .Q(buffer[94]) );
  DFFHQXL buffer_reg_4__31_ ( .D(n914), .CK(clk), .Q(buffer[95]) );
  DFFHQXL buffer_reg_6__24_ ( .D(n982), .CK(clk), .Q(buffer[72]) );
  DFFHQXL buffer_reg_6__25_ ( .D(n981), .CK(clk), .Q(buffer[73]) );
  DFFHQXL buffer_reg_6__26_ ( .D(n980), .CK(clk), .Q(buffer[74]) );
  DFFHQXL buffer_reg_6__27_ ( .D(n979), .CK(clk), .Q(buffer[75]) );
  DFFHQXL buffer_reg_6__28_ ( .D(n978), .CK(clk), .Q(buffer[76]) );
  DFFHQXL buffer_reg_6__29_ ( .D(n977), .CK(clk), .Q(buffer[77]) );
  DFFHQXL buffer_reg_6__30_ ( .D(n976), .CK(clk), .Q(buffer[78]) );
  DFFHQXL buffer_reg_6__31_ ( .D(n975), .CK(clk), .Q(buffer[79]) );
  DFFHQXL buffer_reg_0__24_ ( .D(n797), .CK(clk), .Q(buffer[120]) );
  DFFHQXL buffer_reg_0__25_ ( .D(n796), .CK(clk), .Q(buffer[121]) );
  DFFHQXL buffer_reg_0__26_ ( .D(n795), .CK(clk), .Q(buffer[122]) );
  DFFHQXL buffer_reg_3__24_ ( .D(n890), .CK(clk), .Q(buffer[96]) );
  DFFHQXL buffer_reg_3__25_ ( .D(n889), .CK(clk), .Q(buffer[97]) );
  DFFHQXL buffer_reg_3__26_ ( .D(n888), .CK(clk), .Q(buffer[98]) );
  DFFHQXL buffer_reg_3__27_ ( .D(n887), .CK(clk), .Q(buffer[99]) );
  DFFHQXL buffer_reg_3__28_ ( .D(n886), .CK(clk), .Q(buffer[100]) );
  DFFHQXL buffer_reg_3__29_ ( .D(n885), .CK(clk), .Q(buffer[101]) );
  DFFHQXL buffer_reg_3__30_ ( .D(n884), .CK(clk), .Q(buffer[102]) );
  DFFHQXL buffer_reg_3__31_ ( .D(n883), .CK(clk), .Q(buffer[103]) );
  DFFHQXL buffer_reg_5__24_ ( .D(n951), .CK(clk), .Q(buffer[80]) );
  DFFHQXL buffer_reg_5__25_ ( .D(n950), .CK(clk), .Q(buffer[81]) );
  DFFHQXL buffer_reg_5__26_ ( .D(n949), .CK(clk), .Q(buffer[82]) );
  DFFHQXL buffer_reg_5__27_ ( .D(n948), .CK(clk), .Q(buffer[83]) );
  DFFHQXL buffer_reg_5__28_ ( .D(n947), .CK(clk), .Q(buffer[84]) );
  DFFHQXL buffer_reg_5__29_ ( .D(n946), .CK(clk), .Q(buffer[85]) );
  DFFHQXL buffer_reg_5__30_ ( .D(n945), .CK(clk), .Q(buffer[86]) );
  DFFHQXL buffer_reg_5__31_ ( .D(n944), .CK(clk), .Q(buffer[87]) );
  DFFHQXL buffer_reg_7__24_ ( .D(n1013), .CK(clk), .Q(buffer[64]) );
  DFFHQXL buffer_reg_7__25_ ( .D(n1012), .CK(clk), .Q(buffer[65]) );
  DFFHQXL buffer_reg_7__26_ ( .D(n1011), .CK(clk), .Q(buffer[66]) );
  DFFHQXL buffer_reg_7__27_ ( .D(n1010), .CK(clk), .Q(buffer[67]) );
  DFFHQXL buffer_reg_7__28_ ( .D(n1009), .CK(clk), .Q(buffer[68]) );
  DFFHQXL buffer_reg_7__29_ ( .D(n1008), .CK(clk), .Q(buffer[69]) );
  DFFHQXL buffer_reg_7__30_ ( .D(n1007), .CK(clk), .Q(buffer[70]) );
  DFFHQXL buffer_reg_7__31_ ( .D(n1006), .CK(clk), .Q(buffer[71]) );
  DFFHQXL buffer_reg_1__27_ ( .D(n825), .CK(clk), .Q(buffer[115]) );
  DFFHQXL buffer_reg_1__28_ ( .D(n824), .CK(clk), .Q(buffer[116]) );
  DFFHQXL buffer_reg_1__29_ ( .D(n823), .CK(clk), .Q(buffer[117]) );
  DFFHQXL buffer_reg_1__30_ ( .D(n822), .CK(clk), .Q(buffer[118]) );
  DFFHQXL buffer_reg_1__31_ ( .D(n821), .CK(clk), .Q(buffer[119]) );
  DFFHQXL buffer_reg_1__24_ ( .D(n828), .CK(clk), .Q(buffer[112]) );
  DFFHQXL buffer_reg_1__25_ ( .D(n827), .CK(clk), .Q(buffer[113]) );
  DFFHQXL buffer_reg_1__26_ ( .D(n826), .CK(clk), .Q(buffer[114]) );
  DFFHQXL buffer_reg_0__0_ ( .D(n2218), .CK(clk), .Q(N442) );
  DFFHQXL buffer_reg_0__1_ ( .D(n789), .CK(clk), .Q(N443) );
  DFFHQXL buffer_reg_0__2_ ( .D(n788), .CK(clk), .Q(N444) );
  DFFHQXL buffer_reg_0__3_ ( .D(n787), .CK(clk), .Q(N445) );
  DFFHQXL buffer_reg_2__3_ ( .D(n849), .CK(clk), .Q(N509) );
  DFFHQXL buffer_reg_4__0_ ( .D(n2215), .CK(clk), .Q(N570) );
  DFFHQXL buffer_reg_4__1_ ( .D(n913), .CK(clk), .Q(N571) );
  DFFHQXL buffer_reg_4__2_ ( .D(n912), .CK(clk), .Q(N572) );
  DFFHQXL buffer_reg_4__3_ ( .D(n911), .CK(clk), .Q(N573) );
  DFFHQXL buffer_reg_4__4_ ( .D(n910), .CK(clk), .Q(N574) );
  DFFHQXL buffer_reg_4__5_ ( .D(n909), .CK(clk), .Q(N575) );
  DFFHQXL buffer_reg_4__6_ ( .D(n908), .CK(clk), .Q(N576) );
  DFFHQXL buffer_reg_4__7_ ( .D(n907), .CK(clk), .Q(N577) );
  DFFHQXL buffer_reg_6__0_ ( .D(n2213), .CK(clk), .Q(N634) );
  DFFHQXL buffer_reg_6__1_ ( .D(n974), .CK(clk), .Q(N635) );
  DFFHQXL buffer_reg_6__2_ ( .D(n973), .CK(clk), .Q(N636) );
  DFFHQXL buffer_reg_6__4_ ( .D(n971), .CK(clk), .Q(N638) );
  DFFHQXL buffer_reg_6__5_ ( .D(n970), .CK(clk), .Q(N639) );
  DFFHQXL buffer_reg_6__6_ ( .D(n969), .CK(clk), .Q(N640) );
  DFFHQXL buffer_reg_6__7_ ( .D(n968), .CK(clk), .Q(N641) );
  DFFHQXL buffer_reg_2__0_ ( .D(n2217), .CK(clk), .Q(N506) );
  DFFHQXL buffer_reg_2__1_ ( .D(n851), .CK(clk), .Q(N507) );
  DFFHQXL buffer_reg_2__2_ ( .D(n850), .CK(clk), .Q(N508) );
  DFFHQXL buffer_reg_2__4_ ( .D(n848), .CK(clk), .Q(N510) );
  DFFHQXL buffer_reg_2__5_ ( .D(n847), .CK(clk), .Q(N511) );
  DFFHQXL buffer_reg_2__6_ ( .D(n846), .CK(clk), .Q(N512) );
  DFFHQXL buffer_reg_2__7_ ( .D(n845), .CK(clk), .Q(N513) );
  DFFHQXL buffer_reg_6__3_ ( .D(n972), .CK(clk), .Q(N637) );
  DFFHQXL buffer_reg_0__4_ ( .D(n786), .CK(clk), .Q(N446) );
  DFFHQXL buffer_reg_0__5_ ( .D(n785), .CK(clk), .Q(N447) );
  DFFHQXL buffer_reg_0__6_ ( .D(n784), .CK(clk), .Q(N448) );
  DFFHQXL buffer_reg_0__7_ ( .D(n783), .CK(clk), .Q(N449) );
  DFFHQXL buffer_reg_3__3_ ( .D(n880), .CK(clk), .Q(N541) );
  DFFHQXL buffer_reg_5__0_ ( .D(n2214), .CK(clk), .Q(N602) );
  DFFHQXL buffer_reg_5__1_ ( .D(n943), .CK(clk), .Q(N603) );
  DFFHQXL buffer_reg_5__2_ ( .D(n942), .CK(clk), .Q(N604) );
  DFFHQXL buffer_reg_5__3_ ( .D(n941), .CK(clk), .Q(N605) );
  DFFHQXL buffer_reg_5__4_ ( .D(n940), .CK(clk), .Q(N606) );
  DFFHQXL buffer_reg_5__5_ ( .D(n939), .CK(clk), .Q(N607) );
  DFFHQXL buffer_reg_5__6_ ( .D(n938), .CK(clk), .Q(N608) );
  DFFHQXL buffer_reg_5__7_ ( .D(n937), .CK(clk), .Q(N609) );
  DFFHQXL buffer_reg_7__0_ ( .D(n2212), .CK(clk), .Q(N666) );
  DFFHQXL buffer_reg_7__1_ ( .D(n1005), .CK(clk), .Q(N667) );
  DFFHQXL buffer_reg_7__2_ ( .D(n1004), .CK(clk), .Q(N668) );
  DFFHQXL buffer_reg_7__4_ ( .D(n1002), .CK(clk), .Q(N670) );
  DFFHQXL buffer_reg_7__5_ ( .D(n1001), .CK(clk), .Q(N671) );
  DFFHQXL buffer_reg_7__6_ ( .D(n1000), .CK(clk), .Q(N672) );
  DFFHQXL buffer_reg_7__7_ ( .D(n999), .CK(clk), .Q(N673) );
  DFFHQXL buffer_reg_1__0_ ( .D(n2209), .CK(clk), .Q(N474) );
  DFFHQXL buffer_reg_1__1_ ( .D(n820), .CK(clk), .Q(N475) );
  DFFHQXL buffer_reg_1__2_ ( .D(n819), .CK(clk), .Q(N476) );
  DFFHQXL buffer_reg_1__3_ ( .D(n818), .CK(clk), .Q(N477) );
  DFFHQXL buffer_reg_1__4_ ( .D(n817), .CK(clk), .Q(N478) );
  DFFHQXL buffer_reg_1__5_ ( .D(n816), .CK(clk), .Q(N479) );
  DFFHQXL buffer_reg_1__6_ ( .D(n815), .CK(clk), .Q(N480) );
  DFFHQXL buffer_reg_1__7_ ( .D(n814), .CK(clk), .Q(N481) );
  DFFHQXL buffer_reg_3__0_ ( .D(n2216), .CK(clk), .Q(N538) );
  DFFHQXL buffer_reg_3__1_ ( .D(n882), .CK(clk), .Q(N539) );
  DFFHQXL buffer_reg_3__2_ ( .D(n881), .CK(clk), .Q(N540) );
  DFFHQXL buffer_reg_3__4_ ( .D(n879), .CK(clk), .Q(N542) );
  DFFHQXL buffer_reg_3__5_ ( .D(n878), .CK(clk), .Q(N543) );
  DFFHQXL buffer_reg_3__6_ ( .D(n877), .CK(clk), .Q(N544) );
  DFFHQXL buffer_reg_3__7_ ( .D(n876), .CK(clk), .Q(N545) );
  DFFHQXL buffer_reg_7__3_ ( .D(n1003), .CK(clk), .Q(N669) );
  DFFHQXL buffer_reg_2__19_ ( .D(n864), .CK(clk), .Q(N525) );
  DFFHQXL buffer_reg_2__20_ ( .D(n863), .CK(clk), .Q(N526) );
  DFFHQXL buffer_reg_2__21_ ( .D(n862), .CK(clk), .Q(N527) );
  DFFHQXL buffer_reg_2__22_ ( .D(n861), .CK(clk), .Q(N528) );
  DFFHQXL buffer_reg_2__23_ ( .D(n860), .CK(clk), .Q(N529) );
  DFFHQXL buffer_reg_4__8_ ( .D(n936), .CK(clk), .Q(N578) );
  DFFHQXL buffer_reg_4__9_ ( .D(n935), .CK(clk), .Q(N579) );
  DFFHQXL buffer_reg_4__10_ ( .D(n934), .CK(clk), .Q(N580) );
  DFFHQXL buffer_reg_4__11_ ( .D(n933), .CK(clk), .Q(N581) );
  DFFHQXL buffer_reg_4__12_ ( .D(n932), .CK(clk), .Q(N582) );
  DFFHQXL buffer_reg_4__13_ ( .D(n931), .CK(clk), .Q(N583) );
  DFFHQXL buffer_reg_4__14_ ( .D(n930), .CK(clk), .Q(N584) );
  DFFHQXL buffer_reg_4__15_ ( .D(n929), .CK(clk), .Q(N585) );
  DFFHQXL buffer_reg_4__16_ ( .D(n928), .CK(clk), .Q(N586) );
  DFFHQXL buffer_reg_4__17_ ( .D(n927), .CK(clk), .Q(N587) );
  DFFHQXL buffer_reg_4__18_ ( .D(n926), .CK(clk), .Q(N588) );
  DFFHQXL buffer_reg_4__19_ ( .D(n925), .CK(clk), .Q(N589) );
  DFFHQXL buffer_reg_4__20_ ( .D(n924), .CK(clk), .Q(N590) );
  DFFHQXL buffer_reg_4__21_ ( .D(n923), .CK(clk), .Q(N591) );
  DFFHQXL buffer_reg_4__22_ ( .D(n922), .CK(clk), .Q(N592) );
  DFFHQXL buffer_reg_4__23_ ( .D(n921), .CK(clk), .Q(N593) );
  DFFHQXL buffer_reg_6__8_ ( .D(n998), .CK(clk), .Q(N642) );
  DFFHQXL buffer_reg_6__9_ ( .D(n997), .CK(clk), .Q(N643) );
  DFFHQXL buffer_reg_6__10_ ( .D(n996), .CK(clk), .Q(N644) );
  DFFHQXL buffer_reg_6__11_ ( .D(n995), .CK(clk), .Q(N645) );
  DFFHQXL buffer_reg_6__12_ ( .D(n994), .CK(clk), .Q(N646) );
  DFFHQXL buffer_reg_6__13_ ( .D(n993), .CK(clk), .Q(N647) );
  DFFHQXL buffer_reg_6__14_ ( .D(n992), .CK(clk), .Q(N648) );
  DFFHQXL buffer_reg_6__15_ ( .D(n991), .CK(clk), .Q(N649) );
  DFFHQXL buffer_reg_6__16_ ( .D(n990), .CK(clk), .Q(N650) );
  DFFHQXL buffer_reg_6__17_ ( .D(n989), .CK(clk), .Q(N651) );
  DFFHQXL buffer_reg_6__18_ ( .D(n988), .CK(clk), .Q(N652) );
  DFFHQXL buffer_reg_6__19_ ( .D(n987), .CK(clk), .Q(N653) );
  DFFHQXL buffer_reg_6__20_ ( .D(n986), .CK(clk), .Q(N654) );
  DFFHQXL buffer_reg_6__21_ ( .D(n985), .CK(clk), .Q(N655) );
  DFFHQXL buffer_reg_6__22_ ( .D(n984), .CK(clk), .Q(N656) );
  DFFHQXL buffer_reg_6__23_ ( .D(n983), .CK(clk), .Q(N657) );
  DFFHQXL buffer_reg_2__8_ ( .D(n875), .CK(clk), .Q(N514) );
  DFFHQXL buffer_reg_2__9_ ( .D(n874), .CK(clk), .Q(N515) );
  DFFHQXL buffer_reg_2__10_ ( .D(n873), .CK(clk), .Q(N516) );
  DFFHQXL buffer_reg_2__11_ ( .D(n872), .CK(clk), .Q(N517) );
  DFFHQXL buffer_reg_2__12_ ( .D(n871), .CK(clk), .Q(N518) );
  DFFHQXL buffer_reg_2__13_ ( .D(n870), .CK(clk), .Q(N519) );
  DFFHQXL buffer_reg_2__14_ ( .D(n869), .CK(clk), .Q(N520) );
  DFFHQXL buffer_reg_2__15_ ( .D(n868), .CK(clk), .Q(N521) );
  DFFHQXL buffer_reg_2__16_ ( .D(n867), .CK(clk), .Q(N522) );
  DFFHQXL buffer_reg_2__17_ ( .D(n866), .CK(clk), .Q(N523) );
  DFFHQXL buffer_reg_2__18_ ( .D(n865), .CK(clk), .Q(N524) );
  DFFHQXL buffer_reg_0__8_ ( .D(n813), .CK(clk), .Q(N450) );
  DFFHQXL buffer_reg_0__9_ ( .D(n812), .CK(clk), .Q(N451) );
  DFFHQXL buffer_reg_0__10_ ( .D(n811), .CK(clk), .Q(N452) );
  DFFHQXL buffer_reg_0__11_ ( .D(n810), .CK(clk), .Q(N453) );
  DFFHQXL buffer_reg_3__19_ ( .D(n895), .CK(clk), .Q(N557) );
  DFFHQXL buffer_reg_3__20_ ( .D(n894), .CK(clk), .Q(N558) );
  DFFHQXL buffer_reg_3__21_ ( .D(n893), .CK(clk), .Q(N559) );
  DFFHQXL buffer_reg_3__22_ ( .D(n892), .CK(clk), .Q(N560) );
  DFFHQXL buffer_reg_3__23_ ( .D(n891), .CK(clk), .Q(N561) );
  DFFHQXL buffer_reg_5__8_ ( .D(n967), .CK(clk), .Q(N610) );
  DFFHQXL buffer_reg_5__9_ ( .D(n966), .CK(clk), .Q(N611) );
  DFFHQXL buffer_reg_5__10_ ( .D(n965), .CK(clk), .Q(N612) );
  DFFHQXL buffer_reg_5__11_ ( .D(n964), .CK(clk), .Q(N613) );
  DFFHQXL buffer_reg_5__12_ ( .D(n963), .CK(clk), .Q(N614) );
  DFFHQXL buffer_reg_5__13_ ( .D(n962), .CK(clk), .Q(N615) );
  DFFHQXL buffer_reg_5__14_ ( .D(n961), .CK(clk), .Q(N616) );
  DFFHQXL buffer_reg_5__15_ ( .D(n960), .CK(clk), .Q(N617) );
  DFFHQXL buffer_reg_5__16_ ( .D(n959), .CK(clk), .Q(N618) );
  DFFHQXL buffer_reg_5__17_ ( .D(n958), .CK(clk), .Q(N619) );
  DFFHQXL buffer_reg_5__18_ ( .D(n957), .CK(clk), .Q(N620) );
  DFFHQXL buffer_reg_5__19_ ( .D(n956), .CK(clk), .Q(N621) );
  DFFHQXL buffer_reg_5__20_ ( .D(n955), .CK(clk), .Q(N622) );
  DFFHQXL buffer_reg_5__21_ ( .D(n954), .CK(clk), .Q(N623) );
  DFFHQXL buffer_reg_5__22_ ( .D(n953), .CK(clk), .Q(N624) );
  DFFHQXL buffer_reg_5__23_ ( .D(n952), .CK(clk), .Q(N625) );
  DFFHQXL buffer_reg_7__8_ ( .D(n1029), .CK(clk), .Q(N674) );
  DFFHQXL buffer_reg_7__9_ ( .D(n1028), .CK(clk), .Q(N675) );
  DFFHQXL buffer_reg_7__10_ ( .D(n1027), .CK(clk), .Q(N676) );
  DFFHQXL buffer_reg_7__11_ ( .D(n1026), .CK(clk), .Q(N677) );
  DFFHQXL buffer_reg_7__12_ ( .D(n1025), .CK(clk), .Q(N678) );
  DFFHQXL buffer_reg_7__13_ ( .D(n1024), .CK(clk), .Q(N679) );
  DFFHQXL buffer_reg_7__14_ ( .D(n1023), .CK(clk), .Q(N680) );
  DFFHQXL buffer_reg_7__15_ ( .D(n1022), .CK(clk), .Q(N681) );
  DFFHQXL buffer_reg_7__16_ ( .D(n1021), .CK(clk), .Q(N682) );
  DFFHQXL buffer_reg_7__17_ ( .D(n1020), .CK(clk), .Q(N683) );
  DFFHQXL buffer_reg_7__18_ ( .D(n1019), .CK(clk), .Q(N684) );
  DFFHQXL buffer_reg_7__19_ ( .D(n1018), .CK(clk), .Q(N685) );
  DFFHQXL buffer_reg_7__20_ ( .D(n1017), .CK(clk), .Q(N686) );
  DFFHQXL buffer_reg_7__21_ ( .D(n1016), .CK(clk), .Q(N687) );
  DFFHQXL buffer_reg_7__22_ ( .D(n1015), .CK(clk), .Q(N688) );
  DFFHQXL buffer_reg_7__23_ ( .D(n1014), .CK(clk), .Q(N689) );
  DFFHQXL buffer_reg_1__8_ ( .D(n844), .CK(clk), .Q(N482) );
  DFFHQXL buffer_reg_1__9_ ( .D(n843), .CK(clk), .Q(N483) );
  DFFHQXL buffer_reg_1__10_ ( .D(n842), .CK(clk), .Q(N484) );
  DFFHQXL buffer_reg_1__11_ ( .D(n841), .CK(clk), .Q(N485) );
  DFFHQXL buffer_reg_1__12_ ( .D(n840), .CK(clk), .Q(N486) );
  DFFHQXL buffer_reg_1__13_ ( .D(n839), .CK(clk), .Q(N487) );
  DFFHQXL buffer_reg_1__14_ ( .D(n838), .CK(clk), .Q(N488) );
  DFFHQXL buffer_reg_1__15_ ( .D(n837), .CK(clk), .Q(N489) );
  DFFHQXL buffer_reg_1__16_ ( .D(n836), .CK(clk), .Q(N490) );
  DFFHQXL buffer_reg_1__17_ ( .D(n835), .CK(clk), .Q(N491) );
  DFFHQXL buffer_reg_1__18_ ( .D(n834), .CK(clk), .Q(N492) );
  DFFHQXL buffer_reg_1__19_ ( .D(n833), .CK(clk), .Q(N493) );
  DFFHQXL buffer_reg_1__20_ ( .D(n832), .CK(clk), .Q(N494) );
  DFFHQXL buffer_reg_1__21_ ( .D(n831), .CK(clk), .Q(N495) );
  DFFHQXL buffer_reg_1__22_ ( .D(n830), .CK(clk), .Q(N496) );
  DFFHQXL buffer_reg_1__23_ ( .D(n829), .CK(clk), .Q(N497) );
  DFFHQXL buffer_reg_3__8_ ( .D(n906), .CK(clk), .Q(N546) );
  DFFHQXL buffer_reg_3__9_ ( .D(n905), .CK(clk), .Q(N547) );
  DFFHQXL buffer_reg_3__10_ ( .D(n904), .CK(clk), .Q(N548) );
  DFFHQXL buffer_reg_3__11_ ( .D(n903), .CK(clk), .Q(N549) );
  DFFHQXL buffer_reg_3__12_ ( .D(n902), .CK(clk), .Q(N550) );
  DFFHQXL buffer_reg_3__13_ ( .D(n901), .CK(clk), .Q(N551) );
  DFFHQXL buffer_reg_3__14_ ( .D(n900), .CK(clk), .Q(N552) );
  DFFHQXL buffer_reg_3__15_ ( .D(n899), .CK(clk), .Q(N553) );
  DFFHQXL buffer_reg_3__16_ ( .D(n898), .CK(clk), .Q(N554) );
  DFFHQXL buffer_reg_3__17_ ( .D(n897), .CK(clk), .Q(N555) );
  DFFHQXL buffer_reg_3__18_ ( .D(n896), .CK(clk), .Q(N556) );
  DFFTRX1 R1_reg_23_ ( .D(Wt[23]), .RN(n577), .CK(clk), .Q(R1[23]) );
  DFFHQXL Wt_reg_27_ ( .D(N2160), .CK(clk), .Q(Wt[27]) );
  DFFHQXL Wt_reg_26_ ( .D(N2159), .CK(clk), .Q(Wt[26]) );
  DFFTRX1 R15_reg_2_ ( .D(R14[2]), .RN(n551), .CK(clk), .Q(R15[2]) );
  DFFTRX1 R6_reg_2_ ( .D(R5[2]), .RN(n551), .CK(clk), .Q(R6[2]) );
  DFFHQX2 Wt_reg_18_ ( .D(N2151), .CK(clk), .Q(Wt[18]) );
  DFFTRX4 R15_reg_1_ ( .D(R14[1]), .RN(n550), .CK(clk), .Q(R15[1]) );
  DFFTRX4 R6_reg_1_ ( .D(R5[1]), .RN(n551), .CK(clk), .Q(R6[1]) );
  DFFTRX1 R14_reg_12_ ( .D(R13[12]), .RN(n563), .CK(clk), .Q(R14[12]) );
  DFFTRX1 R1_reg_18_ ( .D(Wt[18]), .RN(n571), .CK(clk), .Q(R1[18]) );
  DFFTRX1 R1_reg_1_ ( .D(Wt[1]), .RN(n551), .CK(clk), .Q(R1[1]) );
  DFFTRX2 R7_reg_0_ ( .D(R6[0]), .RN(n550), .CK(clk), .Q(R7[0]) );
  DFFTRX2 R14_reg_22_ ( .D(R13[22]), .RN(n575), .CK(clk), .Q(R14[22]) );
  DFFTRX2 R1_reg_21_ ( .D(Wt[21]), .RN(n575), .CK(clk), .Q(R1[21]) );
  DFFTRX2 R14_reg_23_ ( .D(R13[23]), .RN(n576), .CK(clk), .Q(R14[23]) );
  DFFTRX2 R1_reg_22_ ( .D(Wt[22]), .RN(n576), .CK(clk), .Q(R1[22]) );
  DFFHQX2 Wt_reg_17_ ( .D(N2150), .CK(clk), .Q(Wt[17]) );
  DFFHQX4 Wt_reg_13_ ( .D(N2146), .CK(clk), .Q(Wt[13]) );
  INVX2 U3 ( .A(logic_result[15]), .Y(n742) );
  INVX4 U4 ( .A(n22), .Y(n675) );
  NAND2XL U5 ( .A(n697), .B(N474), .Y(n1) );
  NAND2X1 U6 ( .A(data[0]), .B(n690), .Y(n2) );
  AND2X2 U7 ( .A(n1), .B(n2), .Y(n1696) );
  CLKINVX3 U8 ( .A(n698), .Y(n697) );
  INVX4 U9 ( .A(n694), .Y(n690) );
  CLKINVX3 U10 ( .A(n1696), .Y(n2209) );
  BUFX16 U11 ( .A(n2228), .Y(Wt[0]) );
  INVX12 U12 ( .A(n640), .Y(n639) );
  NOR2X4 U13 ( .A(n1512), .B(reset), .Y(n1513) );
  INVX4 U14 ( .A(n1657), .Y(n612) );
  INVX8 U15 ( .A(n612), .Y(n611) );
  NOR2X2 U16 ( .A(n660), .B(reset), .Y(n1408) );
  CLKINVX8 U17 ( .A(n661), .Y(n660) );
  INVX2 U18 ( .A(n1416), .Y(n1045) );
  INVX2 U19 ( .A(n1417), .Y(n1046) );
  INVX2 U20 ( .A(n1418), .Y(n1047) );
  INVX2 U21 ( .A(n1419), .Y(n1048) );
  INVX2 U22 ( .A(n1420), .Y(n1049) );
  INVX2 U23 ( .A(n1421), .Y(n1050) );
  INVX2 U24 ( .A(n1422), .Y(n1051) );
  INVX2 U25 ( .A(n1423), .Y(n1052) );
  INVX2 U26 ( .A(n1424), .Y(n1053) );
  INVX2 U27 ( .A(n1425), .Y(n1054) );
  INVX2 U28 ( .A(n1426), .Y(n1055) );
  INVX2 U29 ( .A(n1427), .Y(n1058) );
  AOI31X4 U30 ( .A0(n1546), .A1(n1582), .A2(n1583), .B0(reset), .Y(n1549) );
  CLKINVX3 U31 ( .A(n1549), .Y(n638) );
  INVX16 U32 ( .A(n657), .Y(n655) );
  INVX1 U33 ( .A(n618), .Y(n3) );
  BUFX3 U34 ( .A(n3), .Y(n4) );
  INVX1 U35 ( .A(n619), .Y(n5) );
  BUFX3 U36 ( .A(n5), .Y(n6) );
  CLKINVX2 U37 ( .A(n1621), .Y(n7) );
  CLKINVX2 U38 ( .A(n1621), .Y(n8) );
  CLKINVX3 U39 ( .A(n7), .Y(n9) );
  INVX2 U40 ( .A(n7), .Y(n10) );
  CLKINVX3 U41 ( .A(n8), .Y(n11) );
  INVX4 U42 ( .A(n8), .Y(n12) );
  CLKINVX3 U43 ( .A(n1621), .Y(n618) );
  CLKINVX2 U44 ( .A(n1621), .Y(n619) );
  INVX16 U45 ( .A(n657), .Y(n656) );
  XOR3X4 U46 ( .A(R1[20]), .B(R1[22]), .C(R1[13]), .Y(sigma1[3]) );
  XOR3X4 U47 ( .A(R1[19]), .B(R1[21]), .C(R1[12]), .Y(sigma1[2]) );
  INVX1 U48 ( .A(n1299), .Y(n673) );
  INVX12 U49 ( .A(n693), .Y(n691) );
  XOR3X2 U50 ( .A(R14[21]), .B(R14[10]), .C(R14[6]), .Y(sigma0[3]) );
  NOR2X2 U51 ( .A(n668), .B(reset), .Y(n1336) );
  CLKINVX3 U52 ( .A(n1656), .Y(n616) );
  NAND3BX2 U53 ( .AN(counter1[6]), .B(n1583), .C(n1547), .Y(n1654) );
  AOI31X1 U54 ( .A0(n29), .A1(n1154), .A2(n1440), .B0(reset), .Y(n1442) );
  INVX1 U55 ( .A(n1513), .Y(n640) );
  INVX1 U56 ( .A(n1408), .Y(n657) );
  INVX1 U57 ( .A(n689), .Y(n686) );
  INVX12 U58 ( .A(n693), .Y(n692) );
  CLKINVX3 U59 ( .A(n688), .Y(n687) );
  CLKINVX3 U60 ( .A(n650), .Y(n648) );
  CLKINVX3 U61 ( .A(n643), .Y(n641) );
  INVX1 U62 ( .A(n1177), .Y(n840) );
  AOI22X1 U63 ( .A0(n672), .A1(N609), .B0(data[7]), .B1(n46), .Y(n1324) );
  AOI22X1 U64 ( .A0(n672), .A1(N607), .B0(data[5]), .B1(n45), .Y(n1326) );
  AOI22X1 U65 ( .A0(n672), .A1(N606), .B0(data[4]), .B1(n46), .Y(n1327) );
  AOI22X1 U66 ( .A0(n672), .A1(N605), .B0(data[3]), .B1(n46), .Y(n1328) );
  AOI22X1 U67 ( .A0(n672), .A1(N604), .B0(data[2]), .B1(n44), .Y(n1329) );
  AOI22X1 U68 ( .A0(n672), .A1(N603), .B0(data[1]), .B1(n44), .Y(n1330) );
  AOI22X1 U69 ( .A0(n672), .A1(N602), .B0(data[0]), .B1(n44), .Y(n1331) );
  AOI22X1 U70 ( .A0(n668), .A1(N637), .B0(data[3]), .B1(n61), .Y(n1364) );
  AOI22X1 U71 ( .A0(n668), .A1(N641), .B0(data[7]), .B1(n61), .Y(n1360) );
  AOI22X1 U72 ( .A0(n668), .A1(N639), .B0(data[5]), .B1(n61), .Y(n1362) );
  AOI22X1 U73 ( .A0(n668), .A1(N638), .B0(data[4]), .B1(n61), .Y(n1363) );
  NAND2X2 U74 ( .A(n777), .B(n776), .Y(N2163) );
  NAND2X2 U75 ( .A(logic_result[30]), .B(n417), .Y(n776) );
  INVX1 U76 ( .A(n1431), .Y(n1065) );
  INVX4 U77 ( .A(n622), .Y(n621) );
  INVX1 U78 ( .A(n1620), .Y(n622) );
  INVXL U79 ( .A(n1264), .Y(n678) );
  OR2X2 U80 ( .A(n672), .B(reset), .Y(n21) );
  NOR2X2 U81 ( .A(n664), .B(reset), .Y(n1372) );
  CLKINVX3 U82 ( .A(n1372), .Y(n52) );
  OR2X2 U83 ( .A(n1264), .B(reset), .Y(n22) );
  INVX1 U84 ( .A(n1585), .Y(n630) );
  AOI31X1 U85 ( .A0(n1697), .A1(n29), .A2(n1223), .B0(reset), .Y(n1157) );
  CLKINVX3 U86 ( .A(n56), .Y(n59) );
  CLKINVX3 U87 ( .A(n56), .Y(n60) );
  CLKINVX3 U88 ( .A(n52), .Y(n53) );
  NAND2X1 U89 ( .A(n2082), .B(n2077), .Y(n23) );
  NAND2X1 U90 ( .A(n2074), .B(n2077), .Y(n24) );
  NAND2X1 U91 ( .A(n2074), .B(n2076), .Y(n25) );
  NAND2X1 U92 ( .A(n2076), .B(n2073), .Y(n26) );
  NAND2X1 U93 ( .A(n2076), .B(n2082), .Y(n27) );
  CLKINVX3 U94 ( .A(n681), .Y(n680) );
  AOI2BB1X2 U95 ( .A0N(n1509), .A1N(n1510), .B0(reset), .Y(n1476) );
  CLKINVX3 U96 ( .A(n21), .Y(n45) );
  CLKINVX3 U97 ( .A(n21), .Y(n46) );
  CLKINVX3 U98 ( .A(n21), .Y(n44) );
  CLKINVX3 U99 ( .A(n58), .Y(n61) );
  CLKINVX3 U100 ( .A(n52), .Y(n54) );
  CLKINVX3 U101 ( .A(n1443), .Y(n650) );
  INVX4 U102 ( .A(n650), .Y(n649) );
  AOI2BB1X2 U103 ( .A0N(n1404), .A1N(n1369), .B0(reset), .Y(n1371) );
  AOI2BB1X2 U104 ( .A0N(n1653), .A1N(n1654), .B0(reset), .Y(n1620) );
  INVX1 U105 ( .A(n1335), .Y(n669) );
  INVX2 U106 ( .A(n1586), .Y(n626) );
  INVX4 U107 ( .A(n627), .Y(n624) );
  INVX2 U108 ( .A(n1550), .Y(n634) );
  INVX4 U109 ( .A(n635), .Y(n632) );
  AOI2BB1X2 U110 ( .A0N(n1545), .A1N(n1510), .B0(reset), .Y(n1512) );
  INVX1 U111 ( .A(n1512), .Y(n35) );
  OR2X2 U112 ( .A(n32), .B(n33), .Y(n28) );
  AND3X2 U113 ( .A(n1690), .B(n1547), .C(n1546), .Y(n29) );
  NAND4X1 U114 ( .A(n1333), .B(n1546), .C(n1547), .D(n1440), .Y(n1510) );
  INVX1 U115 ( .A(n702), .Y(n701) );
  CLKINVX3 U116 ( .A(n702), .Y(n700) );
  CLKINVX3 U117 ( .A(n1115), .Y(n702) );
  CLKINVX3 U118 ( .A(n643), .Y(n642) );
  CLKINVX3 U119 ( .A(n661), .Y(n659) );
  CLKINVX3 U120 ( .A(n1407), .Y(n661) );
  INVX4 U121 ( .A(n658), .Y(n654) );
  INVX1 U122 ( .A(n1408), .Y(n658) );
  CLKINVX3 U123 ( .A(n623), .Y(n620) );
  INVXL U124 ( .A(n1620), .Y(n623) );
  NAND2X4 U125 ( .A(n782), .B(n781), .Y(N2164) );
  NOR2X1 U126 ( .A(n652), .B(reset), .Y(n1443) );
  NAND2X4 U127 ( .A(logic_result[31]), .B(n417), .Y(n781) );
  INVXL U128 ( .A(n1191), .Y(n688) );
  CLKINVX3 U129 ( .A(n653), .Y(n651) );
  INVX2 U130 ( .A(n703), .Y(n699) );
  AOI22XL U131 ( .A0(n705), .A1(N453), .B0(N445), .B1(n699), .Y(n1135) );
  CLKINVX3 U132 ( .A(n673), .Y(n672) );
  AOI22X1 U133 ( .A0(n672), .A1(N608), .B0(data[6]), .B1(n46), .Y(n1325) );
  CLKINVX3 U134 ( .A(n1477), .Y(n643) );
  CLKINVX2 U135 ( .A(n616), .Y(n614) );
  INVXL U136 ( .A(n1158), .Y(n693) );
  AND3X2 U137 ( .A(n1297), .B(n1262), .C(n1150), .Y(n1332) );
  CLKINVX3 U138 ( .A(n665), .Y(n664) );
  AOI22X1 U139 ( .A0(n668), .A1(N640), .B0(data[6]), .B1(n60), .Y(n1361) );
  INVX4 U140 ( .A(n669), .Y(n668) );
  INVX2 U141 ( .A(n1442), .Y(n653) );
  AOI31X4 U142 ( .A0(n1260), .A1(n1297), .A2(n29), .B0(reset), .Y(n1264) );
  AND2X4 U143 ( .A(n1152), .B(n1297), .Y(n1405) );
  AOI31X4 U144 ( .A0(n1223), .A1(n1224), .A2(n29), .B0(reset), .Y(n1190) );
  AND2X4 U145 ( .A(n1151), .B(n1224), .Y(n1297) );
  INVX8 U146 ( .A(n685), .Y(n684) );
  AND2X2 U147 ( .A(n676), .B(buffer[88]), .Y(n32) );
  AND2X1 U148 ( .A(N586), .B(n675), .Y(n33) );
  AND3X1 U149 ( .A(n29), .B(n1155), .C(n1440), .Y(n34) );
  NOR2X4 U150 ( .A(n34), .B(reset), .Y(n1407) );
  AND2X4 U151 ( .A(n1150), .B(n1405), .Y(n1440) );
  INVXL U152 ( .A(n35), .Y(n36) );
  INVX1 U153 ( .A(n35), .Y(n37) );
  INVX1 U154 ( .A(n39), .Y(n38) );
  INVX1 U155 ( .A(n1512), .Y(n39) );
  INVX1 U156 ( .A(n39), .Y(n40) );
  INVX1 U157 ( .A(n39), .Y(n41) );
  INVX1 U158 ( .A(n630), .Y(n42) );
  INVX1 U159 ( .A(n630), .Y(n43) );
  AOI31X4 U160 ( .A0(n1546), .A1(n1618), .A2(n1583), .B0(reset), .Y(n1585) );
  INVXL U161 ( .A(n1585), .Y(n631) );
  INVX1 U162 ( .A(n638), .Y(n47) );
  INVX1 U163 ( .A(n638), .Y(n48) );
  INVX12 U164 ( .A(n647), .Y(n49) );
  INVX12 U165 ( .A(n647), .Y(n646) );
  INVX12 U166 ( .A(n647), .Y(n644) );
  INVX12 U167 ( .A(n647), .Y(n645) );
  INVXL U168 ( .A(n1476), .Y(n647) );
  INVX1 U169 ( .A(n52), .Y(n50) );
  BUFX3 U170 ( .A(n50), .Y(n51) );
  INVX1 U171 ( .A(n58), .Y(n55) );
  CLKINVX2 U172 ( .A(n1336), .Y(n56) );
  CLKINVX2 U173 ( .A(n1336), .Y(n58) );
  CLKINVX3 U174 ( .A(n417), .Y(n751) );
  NAND3X2 U175 ( .A(n29), .B(n1405), .C(n1333), .Y(n1369) );
  OAI22XL U176 ( .A0(n733), .A1(n543), .B0(n751), .B1(n732), .Y(N2143) );
  OAI22XL U177 ( .A0(n735), .A1(n543), .B0(n751), .B1(n734), .Y(N2144) );
  OAI22XL U178 ( .A0(n739), .A1(n543), .B0(n751), .B1(n738), .Y(N2146) );
  INVX2 U179 ( .A(n617), .Y(n613) );
  INVXL U180 ( .A(n1586), .Y(n627) );
  INVXL U181 ( .A(n1550), .Y(n635) );
  OAI22XL U182 ( .A0(n713), .A1(n543), .B0(n751), .B1(n712), .Y(N2133) );
  OAI22XL U183 ( .A0(n715), .A1(n543), .B0(n751), .B1(n714), .Y(N2134) );
  OAI22XL U184 ( .A0(n717), .A1(n543), .B0(n751), .B1(n716), .Y(N2135) );
  OAI22XL U185 ( .A0(n721), .A1(n543), .B0(n751), .B1(n720), .Y(N2137) );
  OAI22XL U186 ( .A0(n723), .A1(n543), .B0(n751), .B1(n722), .Y(N2138) );
  OAI22XL U187 ( .A0(n725), .A1(n543), .B0(n751), .B1(n724), .Y(N2139) );
  OAI22XL U188 ( .A0(n727), .A1(n543), .B0(n751), .B1(n726), .Y(N2140) );
  OAI22XL U189 ( .A0(n729), .A1(n543), .B0(n751), .B1(n728), .Y(N2141) );
  OAI22XL U190 ( .A0(n731), .A1(n543), .B0(n751), .B1(n730), .Y(N2142) );
  OAI22XL U191 ( .A0(n737), .A1(n543), .B0(n751), .B1(n736), .Y(N2145) );
  OAI22XL U192 ( .A0(n745), .A1(n543), .B0(n751), .B1(n744), .Y(N2149) );
  NAND3BX1 U193 ( .AN(reset), .B(inner_busy), .C(n2084), .Y(n2067) );
  XOR2X1 U194 ( .A(R1[13]), .B(R1[15]), .Y(sigma1[28]) );
  INVX8 U195 ( .A(n616), .Y(n615) );
  INVX4 U196 ( .A(n653), .Y(n652) );
  INVX2 U197 ( .A(n1226), .Y(n685) );
  INVXL U198 ( .A(n1299), .Y(n674) );
  INVXL U199 ( .A(n1656), .Y(n617) );
  INVX2 U200 ( .A(n1114), .Y(n707) );
  NOR2X4 U201 ( .A(n684), .B(reset), .Y(n1227) );
  NOR2X4 U202 ( .A(n1190), .B(reset), .Y(n1191) );
  AOI22XL U203 ( .A0(n613), .A1(N945), .B0(N937), .B1(n611), .Y(n1665) );
  AOI22XL U204 ( .A0(n621), .A1(N913), .B0(N905), .B1(n9), .Y(n1629) );
  AOI22XL U205 ( .A0(n629), .A1(N881), .B0(N873), .B1(n624), .Y(n1594) );
  AOI22XL U206 ( .A0(n637), .A1(N849), .B0(N841), .B1(n632), .Y(n1558) );
  AOI22XL U207 ( .A0(n37), .A1(N817), .B0(N809), .B1(n639), .Y(n1521) );
  AOI22XL U208 ( .A0(n49), .A1(N785), .B0(N777), .B1(n642), .Y(n1485) );
  AOI22XL U209 ( .A0(n651), .A1(N753), .B0(N745), .B1(n649), .Y(n1451) );
  AOI22XL U210 ( .A0(n659), .A1(N721), .B0(N713), .B1(n655), .Y(n1416) );
  AOI22XL U211 ( .A0(n614), .A1(N933), .B0(N925), .B1(n611), .Y(n1677) );
  AOI22XL U212 ( .A0(n621), .A1(N901), .B0(N893), .B1(n6), .Y(n1641) );
  AOI22XL U213 ( .A0(n42), .A1(N869), .B0(N861), .B1(n624), .Y(n1606) );
  AOI22XL U214 ( .A0(n48), .A1(N837), .B0(N829), .B1(n632), .Y(n1570) );
  AOI22XL U215 ( .A0(n38), .A1(N805), .B0(N797), .B1(n639), .Y(n1533) );
  AOI22XL U216 ( .A0(n49), .A1(N773), .B0(N765), .B1(n641), .Y(n1497) );
  AOI22XL U217 ( .A0(n651), .A1(N741), .B0(N733), .B1(n648), .Y(n1463) );
  AOI22XL U218 ( .A0(n659), .A1(N709), .B0(N701), .B1(n654), .Y(n1428) );
  AOI22XL U219 ( .A0(n664), .A1(N673), .B0(data[7]), .B1(n51), .Y(n1396) );
  AOI22XL U220 ( .A0(n664), .A1(N672), .B0(data[6]), .B1(n53), .Y(n1397) );
  AOI22XL U221 ( .A0(n664), .A1(N671), .B0(data[5]), .B1(n54), .Y(n1398) );
  AOI22XL U222 ( .A0(n664), .A1(N670), .B0(data[4]), .B1(n54), .Y(n1399) );
  AOI22XL U223 ( .A0(n664), .A1(N669), .B0(data[3]), .B1(n54), .Y(n1400) );
  AOI22XL U224 ( .A0(n664), .A1(N668), .B0(data[2]), .B1(n53), .Y(n1401) );
  AOI22XL U225 ( .A0(n664), .A1(N667), .B0(data[1]), .B1(n53), .Y(n1402) );
  AOI22XL U226 ( .A0(n664), .A1(N666), .B0(data[0]), .B1(n53), .Y(n1403) );
  AOI22XL U227 ( .A0(n668), .A1(N636), .B0(data[2]), .B1(n59), .Y(n1365) );
  AOI22XL U228 ( .A0(n668), .A1(N635), .B0(data[1]), .B1(n59), .Y(n1366) );
  AOI22XL U229 ( .A0(n668), .A1(N634), .B0(data[0]), .B1(n60), .Y(n1367) );
  AOI22XL U230 ( .A0(n677), .A1(N577), .B0(data[7]), .B1(n675), .Y(n1289) );
  AOI22XL U231 ( .A0(n1264), .A1(N576), .B0(data[6]), .B1(n675), .Y(n1290) );
  AOI22XL U232 ( .A0(n1264), .A1(N575), .B0(data[5]), .B1(n675), .Y(n1291) );
  AOI22XL U233 ( .A0(n1264), .A1(N574), .B0(data[4]), .B1(n675), .Y(n1292) );
  AOI22XL U234 ( .A0(n1264), .A1(N573), .B0(data[3]), .B1(n675), .Y(n1293) );
  AOI22XL U235 ( .A0(n1264), .A1(N572), .B0(data[2]), .B1(n675), .Y(n1294) );
  AOI22XL U236 ( .A0(n1264), .A1(N571), .B0(data[1]), .B1(n675), .Y(n1295) );
  AOI22XL U237 ( .A0(n1264), .A1(N570), .B0(data[0]), .B1(n675), .Y(n1296) );
  AOI22XL U238 ( .A0(n684), .A1(N545), .B0(data[7]), .B1(n679), .Y(n1251) );
  AOI22XL U239 ( .A0(n684), .A1(N544), .B0(data[6]), .B1(n679), .Y(n1252) );
  AOI22XL U240 ( .A0(n684), .A1(N543), .B0(data[5]), .B1(n679), .Y(n1253) );
  AOI22XL U241 ( .A0(n684), .A1(N542), .B0(data[4]), .B1(n679), .Y(n1254) );
  AOI22XL U242 ( .A0(n684), .A1(N541), .B0(data[3]), .B1(n679), .Y(n1255) );
  AOI22XL U243 ( .A0(n684), .A1(N540), .B0(data[2]), .B1(n679), .Y(n1256) );
  AOI22XL U244 ( .A0(n684), .A1(N539), .B0(data[1]), .B1(n679), .Y(n1257) );
  AOI22XL U245 ( .A0(n684), .A1(N538), .B0(data[0]), .B1(n679), .Y(n1258) );
  NOR2X4 U246 ( .A(n697), .B(reset), .Y(n1158) );
  NOR2X4 U247 ( .A(n706), .B(reset), .Y(n1115) );
  AOI22XL U248 ( .A0(n613), .A1(buffer[7]), .B0(N945), .B1(n611), .Y(n1655) );
  AOI22XL U249 ( .A0(n620), .A1(buffer[15]), .B0(N913), .B1(n6), .Y(n1619) );
  AOI22XL U250 ( .A0(n629), .A1(buffer[23]), .B0(N881), .B1(n625), .Y(n1584)
         );
  AOI22XL U251 ( .A0(n636), .A1(buffer[31]), .B0(N849), .B1(n633), .Y(n1548)
         );
  AOI22XL U252 ( .A0(n40), .A1(buffer[39]), .B0(N817), .B1(n639), .Y(n1511) );
  AOI22XL U253 ( .A0(n646), .A1(buffer[47]), .B0(N785), .B1(n642), .Y(n1475)
         );
  AOI22XL U254 ( .A0(n651), .A1(buffer[55]), .B0(N753), .B1(n649), .Y(n1441)
         );
  AOI22XL U255 ( .A0(n659), .A1(buffer[63]), .B0(N721), .B1(n656), .Y(n1406)
         );
  AOI22XL U256 ( .A0(n1190), .A1(N513), .B0(data[7]), .B1(n686), .Y(n1215) );
  AOI22XL U257 ( .A0(n1190), .A1(N512), .B0(data[6]), .B1(n686), .Y(n1216) );
  AOI22XL U258 ( .A0(n1190), .A1(N511), .B0(data[5]), .B1(n686), .Y(n1217) );
  AOI22XL U259 ( .A0(n1190), .A1(N510), .B0(data[4]), .B1(n686), .Y(n1218) );
  AOI22XL U260 ( .A0(n1190), .A1(N509), .B0(data[3]), .B1(n686), .Y(n1219) );
  AOI22XL U261 ( .A0(n1190), .A1(N508), .B0(data[2]), .B1(n686), .Y(n1220) );
  AOI22XL U262 ( .A0(n1190), .A1(N507), .B0(data[1]), .B1(n686), .Y(n1221) );
  AOI22XL U263 ( .A0(n1190), .A1(N506), .B0(data[0]), .B1(n686), .Y(n1222) );
  AOI22XL U264 ( .A0(n697), .A1(N481), .B0(data[7]), .B1(n690), .Y(n1182) );
  AOI22XL U265 ( .A0(n697), .A1(N480), .B0(data[6]), .B1(n690), .Y(n1183) );
  AOI22XL U266 ( .A0(n697), .A1(N479), .B0(data[5]), .B1(n690), .Y(n1184) );
  AOI22XL U267 ( .A0(n697), .A1(N478), .B0(data[4]), .B1(n690), .Y(n1185) );
  AOI22XL U268 ( .A0(n697), .A1(N477), .B0(data[3]), .B1(n690), .Y(n1186) );
  AOI22XL U269 ( .A0(n697), .A1(N476), .B0(data[2]), .B1(n690), .Y(n1187) );
  AOI22XL U270 ( .A0(n697), .A1(N475), .B0(data[1]), .B1(n690), .Y(n1188) );
  AOI22XL U271 ( .A0(n706), .A1(N449), .B0(data[7]), .B1(n699), .Y(n1139) );
  AOI22XL U272 ( .A0(n706), .A1(N448), .B0(data[6]), .B1(n699), .Y(n1140) );
  AOI22XL U273 ( .A0(n706), .A1(N447), .B0(data[5]), .B1(n699), .Y(n1141) );
  AOI22XL U274 ( .A0(n706), .A1(N446), .B0(data[4]), .B1(n699), .Y(n1142) );
  AOI22XL U275 ( .A0(n706), .A1(N445), .B0(data[3]), .B1(n699), .Y(n1143) );
  AOI22XL U276 ( .A0(n706), .A1(N444), .B0(data[2]), .B1(n699), .Y(n1144) );
  AOI22XL U277 ( .A0(n706), .A1(N443), .B0(data[1]), .B1(n699), .Y(n1145) );
  AOI22XL U278 ( .A0(n706), .A1(N442), .B0(data[0]), .B1(n699), .Y(n1146) );
  XOR2XL U279 ( .A(R1[10]), .B(R1[12]), .Y(sigma1[25]) );
  XOR2XL U280 ( .A(R1[8]), .B(R1[10]), .Y(sigma1[23]) );
  XOR2XL U281 ( .A(R1[9]), .B(R1[11]), .Y(sigma1[24]) );
  XOR2XL U282 ( .A(R1[11]), .B(R1[13]), .Y(sigma1[26]) );
  XOR2XL U283 ( .A(R1[16]), .B(R1[18]), .Y(sigma1[31]) );
  INVX1 U284 ( .A(n600), .Y(n551) );
  INVX1 U285 ( .A(n600), .Y(n552) );
  INVX1 U286 ( .A(n599), .Y(n554) );
  INVX1 U287 ( .A(n598), .Y(n555) );
  INVX1 U288 ( .A(n598), .Y(n556) );
  INVX1 U289 ( .A(n597), .Y(n557) );
  INVX1 U290 ( .A(n597), .Y(n558) );
  INVX1 U291 ( .A(n596), .Y(n559) );
  INVX1 U292 ( .A(n596), .Y(n560) );
  INVX1 U293 ( .A(n595), .Y(n561) );
  INVX1 U294 ( .A(n595), .Y(n562) );
  INVX1 U295 ( .A(n594), .Y(n563) );
  INVX1 U296 ( .A(n594), .Y(n564) );
  INVX1 U297 ( .A(n593), .Y(n565) );
  INVX1 U298 ( .A(n593), .Y(n566) );
  INVX1 U299 ( .A(n592), .Y(n567) );
  INVX1 U300 ( .A(n592), .Y(n568) );
  INVX1 U301 ( .A(n591), .Y(n569) );
  INVX1 U302 ( .A(n591), .Y(n570) );
  INVX1 U303 ( .A(n590), .Y(n571) );
  INVX1 U304 ( .A(n590), .Y(n572) );
  INVX1 U305 ( .A(n589), .Y(n573) );
  INVX1 U306 ( .A(n589), .Y(n574) );
  INVX1 U307 ( .A(n588), .Y(n575) );
  INVX1 U308 ( .A(n588), .Y(n576) );
  INVX1 U309 ( .A(n587), .Y(n577) );
  INVX1 U310 ( .A(n587), .Y(n578) );
  INVX1 U311 ( .A(n587), .Y(n579) );
  INVX1 U312 ( .A(n549), .Y(n580) );
  INVX1 U313 ( .A(n549), .Y(n581) );
  INVX1 U314 ( .A(n599), .Y(n553) );
  INVX1 U315 ( .A(n600), .Y(n550) );
  INVX1 U316 ( .A(n586), .Y(n582) );
  INVX1 U317 ( .A(n586), .Y(n583) );
  INVX1 U318 ( .A(n549), .Y(n584) );
  INVX1 U319 ( .A(n549), .Y(n585) );
  INVX1 U320 ( .A(n2208), .Y(n600) );
  INVX1 U321 ( .A(n547), .Y(n599) );
  INVX1 U322 ( .A(n547), .Y(n598) );
  INVX1 U323 ( .A(n547), .Y(n597) );
  INVX1 U324 ( .A(n546), .Y(n596) );
  INVX1 U325 ( .A(n546), .Y(n595) );
  INVX1 U326 ( .A(n546), .Y(n594) );
  INVX1 U327 ( .A(n545), .Y(n593) );
  INVX1 U328 ( .A(n545), .Y(n592) );
  INVX1 U329 ( .A(n545), .Y(n591) );
  INVX1 U330 ( .A(n544), .Y(n590) );
  INVX1 U331 ( .A(n544), .Y(n589) );
  INVX1 U332 ( .A(n544), .Y(n588) );
  INVX1 U333 ( .A(n544), .Y(n587) );
  INVX1 U334 ( .A(n548), .Y(n547) );
  INVX1 U335 ( .A(n548), .Y(n546) );
  INVX1 U336 ( .A(n548), .Y(n545) );
  INVX1 U337 ( .A(n548), .Y(n544) );
  INVX1 U338 ( .A(n546), .Y(n586) );
  INVX1 U339 ( .A(n24), .Y(n606) );
  INVX1 U340 ( .A(n27), .Y(n604) );
  INVX1 U341 ( .A(n23), .Y(n602) );
  INVX1 U342 ( .A(n26), .Y(n608) );
  INVX1 U343 ( .A(n25), .Y(n610) );
  INVX1 U344 ( .A(n665), .Y(n663) );
  INVX1 U345 ( .A(n669), .Y(n667) );
  INVX1 U346 ( .A(n638), .Y(n636) );
  INVX1 U347 ( .A(n630), .Y(n629) );
  INVX1 U348 ( .A(n638), .Y(n637) );
  INVX1 U349 ( .A(n626), .Y(n625) );
  INVX1 U350 ( .A(n634), .Y(n633) );
  INVX1 U351 ( .A(n698), .Y(n696) );
  INVX1 U352 ( .A(n673), .Y(n671) );
  INVX1 U353 ( .A(n678), .Y(n677) );
  INVX1 U354 ( .A(n685), .Y(n683) );
  INVX1 U355 ( .A(n707), .Y(n705) );
  INVX1 U356 ( .A(n707), .Y(n706) );
  INVX1 U357 ( .A(n543), .Y(n778) );
  INVX1 U358 ( .A(n2208), .Y(n549) );
  INVX1 U359 ( .A(n2208), .Y(n548) );
  NOR2X1 U360 ( .A(n1368), .B(n1404), .Y(n1150) );
  AND3X2 U361 ( .A(n1150), .B(n1695), .C(n1333), .Y(n1260) );
  NOR2X1 U362 ( .A(n1509), .B(n1545), .Y(n1690) );
  AND3X2 U363 ( .A(n1260), .B(n1694), .C(n1262), .Y(n1223) );
  INVX1 U364 ( .A(n25), .Y(n609) );
  INVX1 U365 ( .A(n24), .Y(n605) );
  INVX1 U366 ( .A(n26), .Y(n607) );
  INVX1 U367 ( .A(n27), .Y(n603) );
  INVX1 U368 ( .A(n23), .Y(n601) );
  INVX1 U369 ( .A(n665), .Y(n662) );
  INVX1 U370 ( .A(n1371), .Y(n665) );
  INVX1 U371 ( .A(n669), .Y(n666) );
  INVX1 U372 ( .A(n631), .Y(n628) );
  INVX1 U373 ( .A(n682), .Y(n679) );
  INVX1 U374 ( .A(n1227), .Y(n682) );
  INVX1 U375 ( .A(n1191), .Y(n689) );
  NAND2X1 U376 ( .A(n771), .B(n770), .Y(N2161) );
  OAI21XL U377 ( .A0(n1757), .A1(n1756), .B0(n778), .Y(n771) );
  NAND2X1 U378 ( .A(logic_result[28]), .B(n417), .Y(n770) );
  NAND4X1 U379 ( .A(n1758), .B(n1759), .C(n1760), .D(n1761), .Y(n1757) );
  NAND2X1 U380 ( .A(n773), .B(n772), .Y(N2162) );
  OAI21XL U381 ( .A0(n1746), .A1(n1745), .B0(n778), .Y(n773) );
  NAND2X1 U382 ( .A(logic_result[29]), .B(n417), .Y(n772) );
  NAND4X1 U383 ( .A(n1747), .B(n1748), .C(n1749), .D(n1750), .Y(n1746) );
  OAI21XL U384 ( .A0(n775), .A1(n774), .B0(n778), .Y(n777) );
  NAND4X1 U385 ( .A(n1738), .B(n1739), .C(n1736), .D(n1737), .Y(n775) );
  OAI21XL U386 ( .A0(n780), .A1(n779), .B0(n778), .Y(n782) );
  NAND4X1 U387 ( .A(n1711), .B(n1712), .C(n1709), .D(n1710), .Y(n780) );
  NAND2X1 U388 ( .A(n765), .B(n764), .Y(N2158) );
  OAI21XL U389 ( .A0(n1790), .A1(n1789), .B0(n778), .Y(n765) );
  NAND2X1 U390 ( .A(logic_result[25]), .B(n417), .Y(n764) );
  NAND4X1 U391 ( .A(n1795), .B(n1796), .C(n1797), .D(n1798), .Y(n1789) );
  NAND2X1 U392 ( .A(n767), .B(n766), .Y(N2159) );
  OAI21XL U393 ( .A0(n1779), .A1(n1778), .B0(n778), .Y(n767) );
  NAND2X1 U394 ( .A(logic_result[26]), .B(n417), .Y(n766) );
  NAND4X1 U395 ( .A(n1784), .B(n1785), .C(n1786), .D(n1787), .Y(n1778) );
  NAND2X1 U396 ( .A(n769), .B(n768), .Y(N2160) );
  OAI21XL U397 ( .A0(n1768), .A1(n1767), .B0(n778), .Y(n769) );
  NAND2X1 U398 ( .A(logic_result[27]), .B(n417), .Y(n768) );
  NAND4X1 U399 ( .A(n1769), .B(n1770), .C(n1771), .D(n1772), .Y(n1768) );
  INVX1 U400 ( .A(n1227), .Y(n681) );
  INVX1 U401 ( .A(n708), .Y(n704) );
  INVX1 U402 ( .A(n1114), .Y(n708) );
  INVX1 U403 ( .A(n1158), .Y(n694) );
  INVX1 U404 ( .A(n1115), .Y(n703) );
  NAND2X1 U405 ( .A(n763), .B(n762), .Y(N2157) );
  OAI21XL U406 ( .A0(n1801), .A1(n1800), .B0(n778), .Y(n763) );
  NAND2X1 U407 ( .A(logic_result[24]), .B(n417), .Y(n762) );
  NAND4X1 U408 ( .A(n1806), .B(n1807), .C(n1808), .D(n1809), .Y(n1800) );
  NAND2X1 U409 ( .A(n759), .B(n758), .Y(N2155) );
  OAI21XL U410 ( .A0(n1823), .A1(n1822), .B0(n778), .Y(n759) );
  NAND2X1 U411 ( .A(logic_result[22]), .B(n417), .Y(n758) );
  NAND4X1 U412 ( .A(n1824), .B(n1825), .C(n1826), .D(n1827), .Y(n1823) );
  NAND2X1 U413 ( .A(n761), .B(n760), .Y(N2156) );
  OAI21XL U414 ( .A0(n1812), .A1(n1811), .B0(n778), .Y(n761) );
  NAND2X1 U415 ( .A(logic_result[23]), .B(n417), .Y(n760) );
  NAND4X1 U416 ( .A(n1813), .B(n1814), .C(n1815), .D(n1816), .Y(n1812) );
  INVX1 U417 ( .A(n674), .Y(n670) );
  INVX1 U418 ( .A(n678), .Y(n676) );
  INVX1 U419 ( .A(n698), .Y(n695) );
  INVX1 U420 ( .A(n1157), .Y(n698) );
  INVX1 U421 ( .A(n2067), .Y(n2208) );
  OAI22XL U422 ( .A0(n747), .A1(n543), .B0(n751), .B1(n746), .Y(N2150) );
  NOR2X1 U423 ( .A(n1877), .B(n1878), .Y(n747) );
  INVX1 U424 ( .A(logic_result[17]), .Y(n746) );
  NAND4X1 U425 ( .A(n1883), .B(n1884), .C(n1885), .D(n1886), .Y(n1877) );
  OAI22XL U426 ( .A0(n749), .A1(n543), .B0(n751), .B1(n748), .Y(N2151) );
  NOR2X1 U427 ( .A(n1866), .B(n1867), .Y(n749) );
  INVX1 U428 ( .A(logic_result[18]), .Y(n748) );
  NAND4X1 U429 ( .A(n1872), .B(n1873), .C(n1874), .D(n1875), .Y(n1866) );
  INVX1 U430 ( .A(n2067), .Y(n710) );
  AND2X2 U431 ( .A(n711), .B(n710), .Y(n417) );
  BUFX3 U432 ( .A(n750), .Y(n543) );
  NAND2X1 U433 ( .A(n709), .B(n710), .Y(n750) );
  INVX1 U434 ( .A(n711), .Y(n709) );
  NAND2X1 U435 ( .A(n753), .B(n752), .Y(N2152) );
  OAI21XL U436 ( .A0(n1856), .A1(n1855), .B0(n778), .Y(n753) );
  NAND2X1 U437 ( .A(logic_result[19]), .B(n417), .Y(n752) );
  NAND4X1 U438 ( .A(n1857), .B(n1858), .C(n1859), .D(n1860), .Y(n1856) );
  NAND2X1 U439 ( .A(n755), .B(n754), .Y(N2153) );
  OAI21XL U440 ( .A0(n1845), .A1(n1844), .B0(n778), .Y(n755) );
  NAND2X1 U441 ( .A(logic_result[20]), .B(n417), .Y(n754) );
  NAND4X1 U442 ( .A(n1846), .B(n1847), .C(n1848), .D(n1849), .Y(n1845) );
  NAND2X1 U443 ( .A(n757), .B(n756), .Y(N2154) );
  OAI21XL U444 ( .A0(n1834), .A1(n1833), .B0(n778), .Y(n757) );
  NAND2X1 U445 ( .A(logic_result[21]), .B(n417), .Y(n756) );
  NAND4X1 U446 ( .A(n1835), .B(n1836), .C(n1837), .D(n1838), .Y(n1834) );
  NOR2X1 U447 ( .A(n2031), .B(n2032), .Y(n719) );
  INVX1 U448 ( .A(logic_result[3]), .Y(n718) );
  NAND4X1 U449 ( .A(n2037), .B(n2038), .C(n2039), .D(n2040), .Y(n2031) );
  NOR2X1 U450 ( .A(n2064), .B(n2065), .Y(n713) );
  INVX1 U451 ( .A(logic_result[0]), .Y(n712) );
  NAND4X1 U452 ( .A(n2078), .B(n2079), .C(n2080), .D(n2081), .Y(n2064) );
  NOR2X1 U453 ( .A(n2053), .B(n2054), .Y(n715) );
  INVX1 U454 ( .A(logic_result[1]), .Y(n714) );
  NAND4X1 U455 ( .A(n2059), .B(n2060), .C(n2061), .D(n2062), .Y(n2053) );
  NOR2X1 U456 ( .A(n2042), .B(n2043), .Y(n717) );
  INVX1 U457 ( .A(logic_result[2]), .Y(n716) );
  NAND4X1 U458 ( .A(n2048), .B(n2049), .C(n2050), .D(n2051), .Y(n2042) );
  NOR2X1 U459 ( .A(n2020), .B(n2021), .Y(n721) );
  INVX1 U460 ( .A(logic_result[4]), .Y(n720) );
  NAND4X1 U461 ( .A(n2026), .B(n2027), .C(n2028), .D(n2029), .Y(n2020) );
  NOR2X1 U462 ( .A(n2009), .B(n2010), .Y(n723) );
  INVX1 U463 ( .A(logic_result[5]), .Y(n722) );
  NAND4X1 U464 ( .A(n2015), .B(n2016), .C(n2017), .D(n2018), .Y(n2009) );
  NOR2X1 U465 ( .A(n1998), .B(n1999), .Y(n725) );
  INVX1 U466 ( .A(logic_result[6]), .Y(n724) );
  NAND4X1 U467 ( .A(n2004), .B(n2005), .C(n2006), .D(n2007), .Y(n1998) );
  NOR2X1 U468 ( .A(n1987), .B(n1988), .Y(n727) );
  INVX1 U469 ( .A(logic_result[7]), .Y(n726) );
  NAND4X1 U470 ( .A(n1993), .B(n1994), .C(n1995), .D(n1996), .Y(n1987) );
  NOR2X1 U471 ( .A(n1976), .B(n1977), .Y(n729) );
  INVX1 U472 ( .A(logic_result[8]), .Y(n728) );
  NAND4X1 U473 ( .A(n1982), .B(n1983), .C(n1984), .D(n1985), .Y(n1976) );
  NOR2X1 U474 ( .A(n1965), .B(n1966), .Y(n731) );
  INVX1 U475 ( .A(logic_result[9]), .Y(n730) );
  NAND4X1 U476 ( .A(n1971), .B(n1972), .C(n1973), .D(n1974), .Y(n1965) );
  NOR2X1 U477 ( .A(n1954), .B(n1955), .Y(n733) );
  INVX1 U478 ( .A(logic_result[10]), .Y(n732) );
  NAND4X1 U479 ( .A(n1960), .B(n1961), .C(n1962), .D(n1963), .Y(n1954) );
  NOR2X1 U480 ( .A(n1943), .B(n1944), .Y(n735) );
  INVX1 U481 ( .A(logic_result[11]), .Y(n734) );
  NAND4X1 U482 ( .A(n1949), .B(n1950), .C(n1951), .D(n1952), .Y(n1943) );
  NOR2X1 U483 ( .A(n1932), .B(n1933), .Y(n737) );
  INVX1 U484 ( .A(logic_result[12]), .Y(n736) );
  NAND4X1 U485 ( .A(n1938), .B(n1939), .C(n1940), .D(n1941), .Y(n1932) );
  NOR2X1 U486 ( .A(n1921), .B(n1922), .Y(n739) );
  INVX1 U487 ( .A(logic_result[13]), .Y(n738) );
  NAND4X1 U488 ( .A(n1927), .B(n1928), .C(n1929), .D(n1930), .Y(n1921) );
  OAI22X1 U489 ( .A0(n741), .A1(n543), .B0(n751), .B1(n740), .Y(N2147) );
  NOR2X1 U490 ( .A(n1910), .B(n1911), .Y(n741) );
  INVX1 U491 ( .A(logic_result[14]), .Y(n740) );
  NAND4X1 U492 ( .A(n1916), .B(n1917), .C(n1918), .D(n1919), .Y(n1910) );
  OAI22X1 U493 ( .A0(n743), .A1(n543), .B0(n751), .B1(n742), .Y(N2148) );
  NOR2X1 U494 ( .A(n1899), .B(n1900), .Y(n743) );
  NAND4X1 U495 ( .A(n1905), .B(n1906), .C(n1907), .D(n1908), .Y(n1899) );
  NOR2X1 U496 ( .A(n1888), .B(n1889), .Y(n745) );
  INVX1 U497 ( .A(logic_result[16]), .Y(n744) );
  NAND4X1 U498 ( .A(n1894), .B(n1895), .C(n1896), .D(n1897), .Y(n1888) );
  NAND2X1 U499 ( .A(n1692), .B(n1702), .Y(n1261) );
  NAND2X1 U500 ( .A(n1692), .B(n1693), .Y(n1153) );
  NAND2X1 U501 ( .A(n1692), .B(n1699), .Y(n1691) );
  NAND2X1 U502 ( .A(n1692), .B(n1700), .Y(n1694) );
  NAND2X1 U503 ( .A(n1698), .B(n1699), .Y(n1262) );
  NAND2X1 U504 ( .A(n1701), .B(n1693), .Y(n1155) );
  NAND2X1 U505 ( .A(n1699), .B(n1701), .Y(n1154) );
  NAND2X1 U506 ( .A(n1703), .B(n1693), .Y(n1582) );
  NAND2X1 U507 ( .A(n1699), .B(n1703), .Y(n1618) );
  NAND2X1 U509 ( .A(n1698), .B(n1693), .Y(n1695) );
  AOI31X1 U510 ( .A0(n1332), .A1(n29), .A2(n1333), .B0(reset), .Y(n1299) );
  AOI31X1 U511 ( .A0(n1259), .A1(n29), .A2(n1260), .B0(reset), .Y(n1226) );
  AND3X1 U512 ( .A(n1261), .B(n1262), .C(n1224), .Y(n1259) );
  AOI2BB1X1 U513 ( .A0N(n1368), .A1N(n1369), .B0(reset), .Y(n1335) );
  INVX1 U514 ( .A(n1665), .Y(n2192) );
  INVX1 U515 ( .A(n1666), .Y(n2193) );
  AOI22XL U516 ( .A0(n613), .A1(N944), .B0(N936), .B1(n611), .Y(n1666) );
  INVX1 U517 ( .A(n1667), .Y(n2194) );
  AOI22XL U518 ( .A0(n613), .A1(N943), .B0(N935), .B1(n611), .Y(n1667) );
  INVX1 U519 ( .A(n1668), .Y(n2195) );
  AOI22XL U520 ( .A0(n613), .A1(N942), .B0(N934), .B1(n611), .Y(n1668) );
  INVX1 U521 ( .A(n1669), .Y(n2196) );
  AOI22XL U522 ( .A0(n614), .A1(N941), .B0(N933), .B1(n611), .Y(n1669) );
  INVX1 U523 ( .A(n1670), .Y(n2197) );
  AOI22XL U524 ( .A0(n614), .A1(N940), .B0(N932), .B1(n611), .Y(n1670) );
  INVX1 U525 ( .A(n1671), .Y(n2198) );
  AOI22XL U526 ( .A0(n614), .A1(N939), .B0(N931), .B1(n611), .Y(n1671) );
  INVX1 U527 ( .A(n1672), .Y(n2199) );
  AOI22XL U528 ( .A0(n614), .A1(N938), .B0(N930), .B1(n611), .Y(n1672) );
  INVX1 U529 ( .A(n1673), .Y(n2200) );
  AOI22XL U530 ( .A0(n614), .A1(N937), .B0(N929), .B1(n611), .Y(n1673) );
  INVX1 U531 ( .A(n1674), .Y(n2201) );
  AOI22XL U532 ( .A0(n614), .A1(N936), .B0(N928), .B1(n611), .Y(n1674) );
  INVX1 U533 ( .A(n1675), .Y(n2202) );
  AOI22XL U534 ( .A0(n614), .A1(N935), .B0(N927), .B1(n611), .Y(n1675) );
  INVX1 U535 ( .A(n1676), .Y(n2203) );
  AOI22XL U536 ( .A0(n614), .A1(N934), .B0(N926), .B1(n611), .Y(n1676) );
  INVX1 U537 ( .A(n1677), .Y(n2204) );
  INVX1 U538 ( .A(n1678), .Y(n2205) );
  AOI22XL U539 ( .A0(n614), .A1(N932), .B0(N924), .B1(n611), .Y(n1678) );
  INVX1 U540 ( .A(n1679), .Y(n2206) );
  AOI22XL U541 ( .A0(n614), .A1(N931), .B0(N923), .B1(n611), .Y(n1679) );
  INVX1 U542 ( .A(n1680), .Y(n2207) );
  AOI22XL U543 ( .A0(n614), .A1(N930), .B0(N922), .B1(n611), .Y(n1680) );
  INVX1 U544 ( .A(n1681), .Y(n2177) );
  AOI22XL U545 ( .A0(n615), .A1(N929), .B0(data[7]), .B1(n611), .Y(n1681) );
  INVX1 U546 ( .A(n1682), .Y(n2178) );
  AOI22XL U547 ( .A0(n615), .A1(N928), .B0(data[6]), .B1(n611), .Y(n1682) );
  INVX1 U548 ( .A(n1683), .Y(n2179) );
  AOI22XL U549 ( .A0(n615), .A1(N927), .B0(data[5]), .B1(n611), .Y(n1683) );
  INVX1 U550 ( .A(n1684), .Y(n2180) );
  AOI22XL U551 ( .A0(n615), .A1(N926), .B0(data[4]), .B1(n611), .Y(n1684) );
  INVX1 U552 ( .A(n1685), .Y(n2181) );
  AOI22XL U553 ( .A0(n615), .A1(N925), .B0(data[3]), .B1(n611), .Y(n1685) );
  INVX1 U554 ( .A(n1686), .Y(n2182) );
  AOI22XL U555 ( .A0(n615), .A1(N924), .B0(data[2]), .B1(n611), .Y(n1686) );
  INVX1 U556 ( .A(n1687), .Y(n2183) );
  AOI22XL U557 ( .A0(n615), .A1(N923), .B0(data[1]), .B1(n611), .Y(n1687) );
  INVX1 U558 ( .A(n1688), .Y(n2219) );
  AOI22XL U559 ( .A0(n615), .A1(N922), .B0(data[0]), .B1(n611), .Y(n1688) );
  INVX1 U560 ( .A(n1594), .Y(n2130) );
  INVX1 U561 ( .A(n1595), .Y(n2131) );
  AOI22XL U562 ( .A0(n628), .A1(N880), .B0(N872), .B1(n1586), .Y(n1595) );
  INVX1 U563 ( .A(n1596), .Y(n2132) );
  AOI22XL U564 ( .A0(n42), .A1(N879), .B0(N871), .B1(n624), .Y(n1596) );
  INVX1 U565 ( .A(n1597), .Y(n2133) );
  AOI22XL U566 ( .A0(n43), .A1(N878), .B0(N870), .B1(n1586), .Y(n1597) );
  INVX1 U567 ( .A(n1598), .Y(n2134) );
  AOI22XL U568 ( .A0(n43), .A1(N877), .B0(N869), .B1(n624), .Y(n1598) );
  INVX1 U569 ( .A(n1599), .Y(n2135) );
  AOI22XL U570 ( .A0(n629), .A1(N876), .B0(N868), .B1(n1586), .Y(n1599) );
  INVX1 U571 ( .A(n1600), .Y(n2136) );
  AOI22XL U572 ( .A0(n43), .A1(N875), .B0(N867), .B1(n624), .Y(n1600) );
  INVX1 U573 ( .A(n1601), .Y(n2137) );
  AOI22XL U574 ( .A0(n628), .A1(N874), .B0(N866), .B1(n1586), .Y(n1601) );
  INVX1 U575 ( .A(n1602), .Y(n2138) );
  AOI22XL U576 ( .A0(n42), .A1(N873), .B0(N865), .B1(n624), .Y(n1602) );
  INVX1 U578 ( .A(n1603), .Y(n2139) );
  AOI22XL U579 ( .A0(n43), .A1(N872), .B0(N864), .B1(n1586), .Y(n1603) );
  INVX1 U580 ( .A(n1604), .Y(n2140) );
  AOI22XL U581 ( .A0(n629), .A1(N871), .B0(N863), .B1(n624), .Y(n1604) );
  INVX1 U582 ( .A(n1605), .Y(n2141) );
  AOI22XL U583 ( .A0(n629), .A1(N870), .B0(N862), .B1(n1586), .Y(n1605) );
  INVX1 U584 ( .A(n1606), .Y(n2142) );
  INVX1 U585 ( .A(n1607), .Y(n2143) );
  AOI22XL U586 ( .A0(n628), .A1(N868), .B0(N860), .B1(n624), .Y(n1607) );
  INVX1 U587 ( .A(n1608), .Y(n2144) );
  AOI22XL U588 ( .A0(n42), .A1(N867), .B0(N859), .B1(n624), .Y(n1608) );
  INVX1 U589 ( .A(n1609), .Y(n2145) );
  AOI22XL U590 ( .A0(n43), .A1(N866), .B0(N858), .B1(n624), .Y(n1609) );
  INVX1 U591 ( .A(n1610), .Y(n2115) );
  AOI22XL U592 ( .A0(n628), .A1(N865), .B0(data[7]), .B1(n624), .Y(n1610) );
  INVX1 U593 ( .A(n1611), .Y(n2116) );
  AOI22XL U594 ( .A0(n42), .A1(N864), .B0(data[6]), .B1(n624), .Y(n1611) );
  INVX1 U595 ( .A(n1612), .Y(n2117) );
  AOI22XL U596 ( .A0(n43), .A1(N863), .B0(data[5]), .B1(n624), .Y(n1612) );
  INVX1 U597 ( .A(n1613), .Y(n2118) );
  AOI22XL U598 ( .A0(n629), .A1(N862), .B0(data[4]), .B1(n624), .Y(n1613) );
  INVX1 U599 ( .A(n1614), .Y(n2119) );
  AOI22XL U600 ( .A0(n628), .A1(N861), .B0(data[3]), .B1(n624), .Y(n1614) );
  INVX1 U601 ( .A(n1615), .Y(n2120) );
  AOI22XL U602 ( .A0(n628), .A1(N860), .B0(data[2]), .B1(n624), .Y(n1615) );
  INVX1 U603 ( .A(n1616), .Y(n2121) );
  AOI22XL U604 ( .A0(n628), .A1(N859), .B0(data[1]), .B1(n624), .Y(n1616) );
  INVX1 U605 ( .A(n1617), .Y(n2221) );
  AOI22XL U606 ( .A0(n42), .A1(N858), .B0(data[0]), .B1(n624), .Y(n1617) );
  INVX1 U607 ( .A(n1521), .Y(n1887) );
  INVX1 U608 ( .A(n1522), .Y(n1898) );
  AOI22XL U609 ( .A0(n36), .A1(N816), .B0(N808), .B1(n639), .Y(n1522) );
  INVX1 U610 ( .A(n1523), .Y(n1909) );
  AOI22XL U612 ( .A0(n40), .A1(N815), .B0(N807), .B1(n639), .Y(n1523) );
  INVX1 U613 ( .A(n1524), .Y(n1920) );
  AOI22XL U614 ( .A0(n37), .A1(N814), .B0(N806), .B1(n639), .Y(n1524) );
  INVX1 U615 ( .A(n1525), .Y(n1931) );
  AOI22XL U616 ( .A0(n41), .A1(N813), .B0(N805), .B1(n639), .Y(n1525) );
  INVX1 U617 ( .A(n1526), .Y(n1942) );
  AOI22XL U618 ( .A0(n37), .A1(N812), .B0(N804), .B1(n1513), .Y(n1526) );
  INVX1 U619 ( .A(n1527), .Y(n1953) );
  AOI22XL U620 ( .A0(n41), .A1(N811), .B0(N803), .B1(n1513), .Y(n1527) );
  INVX1 U621 ( .A(n1528), .Y(n1964) );
  AOI22XL U622 ( .A0(n41), .A1(N810), .B0(N802), .B1(n1513), .Y(n1528) );
  INVX1 U623 ( .A(n1529), .Y(n1975) );
  AOI22XL U624 ( .A0(n36), .A1(N809), .B0(N801), .B1(n1513), .Y(n1529) );
  INVX1 U625 ( .A(n1530), .Y(n1986) );
  AOI22XL U626 ( .A0(n38), .A1(N808), .B0(N800), .B1(n1513), .Y(n1530) );
  INVX1 U627 ( .A(n1531), .Y(n1997) );
  AOI22XL U628 ( .A0(n41), .A1(N807), .B0(N799), .B1(n1513), .Y(n1531) );
  INVX1 U629 ( .A(n1532), .Y(n2008) );
  AOI22XL U630 ( .A0(n38), .A1(N806), .B0(N798), .B1(n1513), .Y(n1532) );
  INVX1 U631 ( .A(n1533), .Y(n2019) );
  INVX1 U632 ( .A(n1534), .Y(n2030) );
  AOI22XL U633 ( .A0(n37), .A1(N804), .B0(N796), .B1(n639), .Y(n1534) );
  INVX1 U634 ( .A(n1535), .Y(n2041) );
  AOI22XL U635 ( .A0(n40), .A1(N803), .B0(N795), .B1(n639), .Y(n1535) );
  INVX1 U636 ( .A(n1536), .Y(n2052) );
  AOI22XL U637 ( .A0(n36), .A1(N802), .B0(N794), .B1(n639), .Y(n1536) );
  INVX1 U638 ( .A(n1537), .Y(n1734) );
  AOI22XL U639 ( .A0(n40), .A1(N801), .B0(data[7]), .B1(n639), .Y(n1537) );
  INVX1 U640 ( .A(n1538), .Y(n1735) );
  AOI22XL U641 ( .A0(n41), .A1(N800), .B0(data[6]), .B1(n639), .Y(n1538) );
  INVX1 U642 ( .A(n1539), .Y(n1744) );
  AOI22XL U643 ( .A0(n41), .A1(N799), .B0(data[5]), .B1(n639), .Y(n1539) );
  INVX1 U644 ( .A(n1540), .Y(n1755) );
  AOI22XL U646 ( .A0(n37), .A1(N798), .B0(data[4]), .B1(n639), .Y(n1540) );
  INVX1 U647 ( .A(n1541), .Y(n1766) );
  AOI22XL U648 ( .A0(n38), .A1(N797), .B0(data[3]), .B1(n639), .Y(n1541) );
  INVX1 U649 ( .A(n1542), .Y(n1777) );
  AOI22XL U650 ( .A0(n36), .A1(N796), .B0(data[2]), .B1(n639), .Y(n1542) );
  INVX1 U651 ( .A(n1543), .Y(n1788) );
  AOI22XL U652 ( .A0(n37), .A1(N795), .B0(data[1]), .B1(n639), .Y(n1543) );
  INVX1 U653 ( .A(n1544), .Y(n2224) );
  AOI22XL U654 ( .A0(n37), .A1(N794), .B0(data[0]), .B1(n639), .Y(n1544) );
  INVX1 U655 ( .A(n1451), .Y(n1081) );
  INVX1 U656 ( .A(n1452), .Y(n1082) );
  AOI22XL U657 ( .A0(n651), .A1(N752), .B0(N744), .B1(n649), .Y(n1452) );
  INVX1 U658 ( .A(n1453), .Y(n1083) );
  AOI22XL U659 ( .A0(n651), .A1(N751), .B0(N743), .B1(n649), .Y(n1453) );
  INVX1 U660 ( .A(n1454), .Y(n1084) );
  AOI22XL U661 ( .A0(n651), .A1(N750), .B0(N742), .B1(n649), .Y(n1454) );
  INVX1 U662 ( .A(n1455), .Y(n1085) );
  AOI22XL U663 ( .A0(n651), .A1(N749), .B0(N741), .B1(n649), .Y(n1455) );
  INVX1 U664 ( .A(n1456), .Y(n1086) );
  AOI22XL U665 ( .A0(n651), .A1(N748), .B0(N740), .B1(n649), .Y(n1456) );
  INVX1 U666 ( .A(n1457), .Y(n1087) );
  AOI22XL U667 ( .A0(n651), .A1(N747), .B0(N739), .B1(n649), .Y(n1457) );
  INVX1 U668 ( .A(n1458), .Y(n1088) );
  AOI22XL U669 ( .A0(n651), .A1(N746), .B0(N738), .B1(n649), .Y(n1458) );
  INVX1 U670 ( .A(n1459), .Y(n1089) );
  AOI22XL U671 ( .A0(n651), .A1(N745), .B0(N737), .B1(n649), .Y(n1459) );
  INVX1 U672 ( .A(n1460), .Y(n1090) );
  AOI22XL U673 ( .A0(n651), .A1(N744), .B0(N736), .B1(n649), .Y(n1460) );
  INVX1 U674 ( .A(n1461), .Y(n1091) );
  AOI22XL U675 ( .A0(n651), .A1(N743), .B0(N735), .B1(n649), .Y(n1461) );
  INVX1 U676 ( .A(n1462), .Y(n1092) );
  AOI22XL U677 ( .A0(n651), .A1(N742), .B0(N734), .B1(n649), .Y(n1462) );
  INVX1 U678 ( .A(n1463), .Y(n1093) );
  INVX1 U681 ( .A(n1464), .Y(n1094) );
  AOI22XL U683 ( .A0(n651), .A1(N740), .B0(N732), .B1(n648), .Y(n1464) );
  INVX1 U684 ( .A(n1465), .Y(n1095) );
  AOI22XL U685 ( .A0(n651), .A1(N739), .B0(N731), .B1(n648), .Y(n1465) );
  INVX1 U687 ( .A(n1466), .Y(n1096) );
  AOI22XL U690 ( .A0(n651), .A1(N738), .B0(N730), .B1(n648), .Y(n1466) );
  INVX1 U691 ( .A(n1467), .Y(n1066) );
  AOI22XL U692 ( .A0(n652), .A1(N737), .B0(data[7]), .B1(n648), .Y(n1467) );
  INVX1 U693 ( .A(n1468), .Y(n1067) );
  AOI22XL U694 ( .A0(n652), .A1(N736), .B0(data[6]), .B1(n648), .Y(n1468) );
  INVX1 U695 ( .A(n1469), .Y(n1068) );
  AOI22XL U696 ( .A0(n652), .A1(N735), .B0(data[5]), .B1(n648), .Y(n1469) );
  INVX1 U698 ( .A(n1470), .Y(n1069) );
  AOI22XL U699 ( .A0(n652), .A1(N734), .B0(data[4]), .B1(n648), .Y(n1470) );
  INVX1 U700 ( .A(n1471), .Y(n1070) );
  AOI22XL U701 ( .A0(n652), .A1(N733), .B0(data[3]), .B1(n648), .Y(n1471) );
  INVX1 U704 ( .A(n1472), .Y(n1071) );
  AOI22XL U705 ( .A0(n652), .A1(N732), .B0(data[2]), .B1(n648), .Y(n1472) );
  INVX1 U706 ( .A(n1473), .Y(n1072) );
  AOI22XL U710 ( .A0(n652), .A1(N731), .B0(data[1]), .B1(n648), .Y(n1473) );
  INVX1 U711 ( .A(n1474), .Y(n2210) );
  AOI22XL U712 ( .A0(n652), .A1(N730), .B0(data[0]), .B1(n648), .Y(n1474) );
  INVX1 U713 ( .A(n1380), .Y(n1014) );
  AOI22X1 U714 ( .A0(n662), .A1(N689), .B0(N681), .B1(n51), .Y(n1380) );
  INVX1 U717 ( .A(n1381), .Y(n1015) );
  AOI22X1 U718 ( .A0(n662), .A1(N688), .B0(N680), .B1(n53), .Y(n1381) );
  INVX1 U719 ( .A(n1382), .Y(n1016) );
  AOI22X1 U720 ( .A0(n662), .A1(N687), .B0(N679), .B1(n54), .Y(n1382) );
  INVX1 U721 ( .A(n1383), .Y(n1017) );
  AOI22X1 U722 ( .A0(n662), .A1(N686), .B0(N678), .B1(n51), .Y(n1383) );
  INVX1 U723 ( .A(n1384), .Y(n1018) );
  AOI22X1 U724 ( .A0(n663), .A1(N685), .B0(N677), .B1(n53), .Y(n1384) );
  INVX1 U725 ( .A(n1385), .Y(n1019) );
  AOI22X1 U726 ( .A0(n663), .A1(N684), .B0(N676), .B1(n53), .Y(n1385) );
  INVX1 U727 ( .A(n1386), .Y(n1020) );
  AOI22X1 U728 ( .A0(n663), .A1(N683), .B0(N675), .B1(n53), .Y(n1386) );
  INVX1 U729 ( .A(n1387), .Y(n1021) );
  AOI22X1 U730 ( .A0(n663), .A1(N682), .B0(N674), .B1(n54), .Y(n1387) );
  INVX1 U731 ( .A(n1388), .Y(n1022) );
  AOI22X1 U732 ( .A0(n663), .A1(N681), .B0(N673), .B1(n54), .Y(n1388) );
  INVX1 U733 ( .A(n1389), .Y(n1023) );
  AOI22X1 U734 ( .A0(n663), .A1(N680), .B0(N672), .B1(n53), .Y(n1389) );
  INVX1 U735 ( .A(n1390), .Y(n1024) );
  AOI22X1 U736 ( .A0(n663), .A1(N679), .B0(N671), .B1(n54), .Y(n1390) );
  INVX1 U737 ( .A(n1391), .Y(n1025) );
  AOI22X1 U738 ( .A0(n663), .A1(N678), .B0(N670), .B1(n54), .Y(n1391) );
  INVX1 U739 ( .A(n1392), .Y(n1026) );
  AOI22X1 U740 ( .A0(n663), .A1(N677), .B0(N669), .B1(n54), .Y(n1392) );
  INVX1 U741 ( .A(n1393), .Y(n1027) );
  AOI22X1 U742 ( .A0(n663), .A1(N676), .B0(N668), .B1(n54), .Y(n1393) );
  INVX1 U743 ( .A(n1394), .Y(n1028) );
  AOI22X1 U744 ( .A0(n663), .A1(N675), .B0(N667), .B1(n53), .Y(n1394) );
  INVX1 U745 ( .A(n1395), .Y(n1029) );
  AOI22X1 U746 ( .A0(n663), .A1(N674), .B0(N666), .B1(n54), .Y(n1395) );
  INVX1 U747 ( .A(n1396), .Y(n999) );
  INVX1 U748 ( .A(n1397), .Y(n1000) );
  INVX1 U749 ( .A(n1398), .Y(n1001) );
  INVX1 U750 ( .A(n1399), .Y(n1002) );
  INVX1 U751 ( .A(n1400), .Y(n1003) );
  INVX1 U752 ( .A(n1401), .Y(n1004) );
  INVX1 U753 ( .A(n1402), .Y(n1005) );
  INVX1 U754 ( .A(n1403), .Y(n2212) );
  INVX1 U755 ( .A(n1308), .Y(n952) );
  AOI22X1 U756 ( .A0(n670), .A1(N625), .B0(N617), .B1(n46), .Y(n1308) );
  INVX1 U757 ( .A(n1309), .Y(n953) );
  AOI22X1 U758 ( .A0(n670), .A1(N624), .B0(N616), .B1(n44), .Y(n1309) );
  INVX1 U759 ( .A(n1310), .Y(n954) );
  AOI22X1 U760 ( .A0(n670), .A1(N623), .B0(N615), .B1(n45), .Y(n1310) );
  INVX1 U761 ( .A(n1311), .Y(n955) );
  AOI22X1 U762 ( .A0(n670), .A1(N622), .B0(N614), .B1(n45), .Y(n1311) );
  INVX1 U763 ( .A(n1312), .Y(n956) );
  AOI22X1 U764 ( .A0(n671), .A1(N621), .B0(N613), .B1(n44), .Y(n1312) );
  INVX1 U765 ( .A(n1313), .Y(n957) );
  AOI22X1 U766 ( .A0(n671), .A1(N620), .B0(N612), .B1(n46), .Y(n1313) );
  INVX1 U767 ( .A(n1314), .Y(n958) );
  AOI22X1 U768 ( .A0(n671), .A1(N619), .B0(N611), .B1(n44), .Y(n1314) );
  INVX1 U769 ( .A(n1315), .Y(n959) );
  AOI22X1 U770 ( .A0(n671), .A1(N618), .B0(N610), .B1(n45), .Y(n1315) );
  INVX1 U771 ( .A(n1316), .Y(n960) );
  AOI22X1 U772 ( .A0(n671), .A1(N617), .B0(N609), .B1(n46), .Y(n1316) );
  INVX1 U773 ( .A(n1317), .Y(n961) );
  AOI22X1 U774 ( .A0(n671), .A1(N616), .B0(N608), .B1(n45), .Y(n1317) );
  INVX1 U775 ( .A(n1318), .Y(n962) );
  AOI22X1 U776 ( .A0(n671), .A1(N615), .B0(N607), .B1(n45), .Y(n1318) );
  INVX1 U777 ( .A(n1319), .Y(n963) );
  AOI22X1 U778 ( .A0(n671), .A1(N614), .B0(N606), .B1(n46), .Y(n1319) );
  INVX1 U779 ( .A(n1320), .Y(n964) );
  AOI22X1 U780 ( .A0(n671), .A1(N613), .B0(N605), .B1(n45), .Y(n1320) );
  INVX1 U781 ( .A(n1321), .Y(n965) );
  AOI22X1 U782 ( .A0(n671), .A1(N612), .B0(N604), .B1(n46), .Y(n1321) );
  INVX1 U783 ( .A(n1322), .Y(n966) );
  AOI22X1 U784 ( .A0(n671), .A1(N611), .B0(N603), .B1(n44), .Y(n1322) );
  INVX1 U785 ( .A(n1323), .Y(n967) );
  AOI22X1 U786 ( .A0(n671), .A1(N610), .B0(N602), .B1(n45), .Y(n1323) );
  INVX1 U787 ( .A(n1324), .Y(n937) );
  INVX1 U788 ( .A(n1325), .Y(n938) );
  INVX1 U789 ( .A(n1326), .Y(n939) );
  INVX1 U790 ( .A(n1327), .Y(n940) );
  INVX1 U791 ( .A(n1328), .Y(n941) );
  INVX1 U792 ( .A(n1329), .Y(n942) );
  INVX1 U793 ( .A(n1330), .Y(n943) );
  INVX1 U794 ( .A(n1331), .Y(n2214) );
  INVX1 U795 ( .A(n1235), .Y(n891) );
  AOI22X1 U796 ( .A0(n683), .A1(N561), .B0(N553), .B1(n680), .Y(n1235) );
  INVX1 U797 ( .A(n1236), .Y(n892) );
  AOI22X1 U798 ( .A0(n683), .A1(N560), .B0(N552), .B1(n680), .Y(n1236) );
  INVX1 U799 ( .A(n1237), .Y(n893) );
  AOI22X1 U800 ( .A0(n683), .A1(N559), .B0(N551), .B1(n680), .Y(n1237) );
  INVX1 U801 ( .A(n1238), .Y(n894) );
  AOI22X1 U802 ( .A0(n683), .A1(N558), .B0(N550), .B1(n680), .Y(n1238) );
  INVX1 U803 ( .A(n1239), .Y(n895) );
  AOI22X1 U804 ( .A0(n683), .A1(N557), .B0(N549), .B1(n680), .Y(n1239) );
  INVX1 U805 ( .A(n1240), .Y(n896) );
  AOI22X1 U806 ( .A0(n683), .A1(N556), .B0(N548), .B1(n680), .Y(n1240) );
  INVX1 U807 ( .A(n1241), .Y(n897) );
  AOI22X1 U808 ( .A0(n683), .A1(N555), .B0(N547), .B1(n680), .Y(n1241) );
  INVX1 U809 ( .A(n1242), .Y(n898) );
  AOI22X1 U810 ( .A0(n683), .A1(N554), .B0(N546), .B1(n680), .Y(n1242) );
  INVX1 U811 ( .A(n1243), .Y(n899) );
  AOI22X1 U812 ( .A0(n683), .A1(N553), .B0(N545), .B1(n680), .Y(n1243) );
  INVX1 U813 ( .A(n1244), .Y(n900) );
  AOI22X1 U814 ( .A0(n683), .A1(N552), .B0(N544), .B1(n680), .Y(n1244) );
  INVX1 U815 ( .A(n1245), .Y(n901) );
  AOI22X1 U816 ( .A0(n683), .A1(N551), .B0(N543), .B1(n680), .Y(n1245) );
  INVX1 U817 ( .A(n1246), .Y(n902) );
  AOI22X1 U818 ( .A0(n683), .A1(N550), .B0(N542), .B1(n680), .Y(n1246) );
  INVX1 U819 ( .A(n1247), .Y(n903) );
  AOI22X1 U820 ( .A0(n683), .A1(N549), .B0(N541), .B1(n679), .Y(n1247) );
  INVX1 U821 ( .A(n1248), .Y(n904) );
  AOI22X1 U822 ( .A0(n683), .A1(N548), .B0(N540), .B1(n679), .Y(n1248) );
  INVX1 U823 ( .A(n1249), .Y(n905) );
  AOI22X1 U824 ( .A0(n683), .A1(N547), .B0(N539), .B1(n679), .Y(n1249) );
  INVX1 U825 ( .A(n1250), .Y(n906) );
  AOI22X1 U826 ( .A0(n683), .A1(N546), .B0(N538), .B1(n679), .Y(n1250) );
  INVX1 U827 ( .A(n1251), .Y(n876) );
  INVX1 U828 ( .A(n1252), .Y(n877) );
  INVX1 U829 ( .A(n1253), .Y(n878) );
  INVX1 U830 ( .A(n1254), .Y(n879) );
  INVX1 U831 ( .A(n1255), .Y(n880) );
  INVX1 U832 ( .A(n1256), .Y(n881) );
  INVX1 U833 ( .A(n1257), .Y(n882) );
  INVX1 U834 ( .A(n1258), .Y(n2216) );
  INVX1 U835 ( .A(n1629), .Y(n2161) );
  INVX1 U836 ( .A(n1630), .Y(n2162) );
  AOI22XL U837 ( .A0(n621), .A1(N912), .B0(N904), .B1(n10), .Y(n1630) );
  INVX1 U838 ( .A(n1631), .Y(n2163) );
  AOI22XL U839 ( .A0(n620), .A1(N911), .B0(N903), .B1(n9), .Y(n1631) );
  INVX1 U840 ( .A(n1632), .Y(n2164) );
  AOI22XL U841 ( .A0(n621), .A1(N910), .B0(N902), .B1(n10), .Y(n1632) );
  INVX1 U842 ( .A(n1633), .Y(n2165) );
  AOI22XL U843 ( .A0(n621), .A1(N909), .B0(N901), .B1(n6), .Y(n1633) );
  INVX1 U844 ( .A(n1634), .Y(n2166) );
  AOI22XL U845 ( .A0(n620), .A1(N908), .B0(N900), .B1(n4), .Y(n1634) );
  INVX1 U846 ( .A(n1635), .Y(n2167) );
  AOI22XL U847 ( .A0(n621), .A1(N907), .B0(N899), .B1(n11), .Y(n1635) );
  INVX1 U848 ( .A(n1636), .Y(n2168) );
  AOI22XL U849 ( .A0(n620), .A1(N906), .B0(N898), .B1(n12), .Y(n1636) );
  INVX1 U850 ( .A(n1637), .Y(n2169) );
  AOI22XL U851 ( .A0(n621), .A1(N905), .B0(N897), .B1(n10), .Y(n1637) );
  INVX1 U852 ( .A(n1638), .Y(n2170) );
  AOI22XL U853 ( .A0(n620), .A1(N904), .B0(N896), .B1(n11), .Y(n1638) );
  INVX1 U854 ( .A(n1639), .Y(n2171) );
  AOI22XL U855 ( .A0(n621), .A1(N903), .B0(N895), .B1(n9), .Y(n1639) );
  INVX1 U856 ( .A(n1640), .Y(n2172) );
  AOI22XL U857 ( .A0(n621), .A1(N902), .B0(N894), .B1(n10), .Y(n1640) );
  INVX1 U858 ( .A(n1641), .Y(n2173) );
  INVX1 U859 ( .A(n1642), .Y(n2174) );
  AOI22XL U860 ( .A0(n620), .A1(N900), .B0(N892), .B1(n4), .Y(n1642) );
  INVX1 U861 ( .A(n1643), .Y(n2175) );
  AOI22XL U862 ( .A0(n621), .A1(N899), .B0(N891), .B1(n11), .Y(n1643) );
  INVX1 U863 ( .A(n1644), .Y(n2176) );
  AOI22XL U864 ( .A0(n620), .A1(N898), .B0(N890), .B1(n12), .Y(n1644) );
  INVX1 U865 ( .A(n1645), .Y(n2146) );
  AOI22XL U866 ( .A0(n621), .A1(N897), .B0(data[7]), .B1(n11), .Y(n1645) );
  INVX1 U867 ( .A(n1646), .Y(n2147) );
  AOI22XL U868 ( .A0(n621), .A1(N896), .B0(data[6]), .B1(n12), .Y(n1646) );
  INVX1 U869 ( .A(n1647), .Y(n2148) );
  AOI22XL U870 ( .A0(n621), .A1(N895), .B0(data[5]), .B1(n9), .Y(n1647) );
  INVX1 U871 ( .A(n1648), .Y(n2149) );
  AOI22XL U872 ( .A0(n621), .A1(N894), .B0(data[4]), .B1(n10), .Y(n1648) );
  INVX1 U873 ( .A(n1649), .Y(n2150) );
  AOI22XL U874 ( .A0(n621), .A1(N893), .B0(data[3]), .B1(n12), .Y(n1649) );
  INVX1 U875 ( .A(n1650), .Y(n2151) );
  AOI22XL U876 ( .A0(n621), .A1(N892), .B0(data[2]), .B1(n6), .Y(n1650) );
  INVX1 U877 ( .A(n1651), .Y(n2152) );
  AOI22XL U878 ( .A0(n620), .A1(N891), .B0(data[1]), .B1(n6), .Y(n1651) );
  INVX1 U879 ( .A(n1652), .Y(n2220) );
  AOI22XL U880 ( .A0(n1620), .A1(N890), .B0(data[0]), .B1(n4), .Y(n1652) );
  INVX1 U881 ( .A(n1558), .Y(n2099) );
  INVX1 U882 ( .A(n1559), .Y(n2100) );
  AOI22XL U883 ( .A0(n637), .A1(N848), .B0(N840), .B1(n1550), .Y(n1559) );
  INVX1 U884 ( .A(n1560), .Y(n2101) );
  AOI22XL U885 ( .A0(n636), .A1(N847), .B0(N839), .B1(n632), .Y(n1560) );
  INVX1 U886 ( .A(n1561), .Y(n2102) );
  AOI22XL U887 ( .A0(n47), .A1(N846), .B0(N838), .B1(n1550), .Y(n1561) );
  INVX1 U888 ( .A(n1562), .Y(n2103) );
  AOI22XL U889 ( .A0(n636), .A1(N845), .B0(N837), .B1(n632), .Y(n1562) );
  INVX1 U890 ( .A(n1563), .Y(n2104) );
  AOI22XL U891 ( .A0(n636), .A1(N844), .B0(N836), .B1(n1550), .Y(n1563) );
  INVX1 U892 ( .A(n1564), .Y(n2105) );
  AOI22XL U893 ( .A0(n637), .A1(N843), .B0(N835), .B1(n632), .Y(n1564) );
  INVX1 U894 ( .A(n1565), .Y(n2106) );
  AOI22XL U895 ( .A0(n47), .A1(N842), .B0(N834), .B1(n1550), .Y(n1565) );
  INVX1 U896 ( .A(n1566), .Y(n2107) );
  AOI22XL U897 ( .A0(n48), .A1(N841), .B0(N833), .B1(n632), .Y(n1566) );
  INVX1 U898 ( .A(n1567), .Y(n2108) );
  AOI22XL U899 ( .A0(n637), .A1(N840), .B0(N832), .B1(n1550), .Y(n1567) );
  INVX1 U900 ( .A(n1568), .Y(n2109) );
  AOI22XL U901 ( .A0(n48), .A1(N839), .B0(N831), .B1(n632), .Y(n1568) );
  INVX1 U902 ( .A(n1569), .Y(n2110) );
  AOI22XL U903 ( .A0(n636), .A1(N838), .B0(N830), .B1(n1550), .Y(n1569) );
  INVX1 U904 ( .A(n1570), .Y(n2111) );
  INVX1 U905 ( .A(n1571), .Y(n2112) );
  AOI22XL U906 ( .A0(n48), .A1(N836), .B0(N828), .B1(n632), .Y(n1571) );
  INVX1 U907 ( .A(n1572), .Y(n2113) );
  AOI22XL U908 ( .A0(n47), .A1(N835), .B0(N827), .B1(n632), .Y(n1572) );
  INVX1 U909 ( .A(n1573), .Y(n2114) );
  AOI22XL U910 ( .A0(n637), .A1(N834), .B0(N826), .B1(n632), .Y(n1573) );
  INVX1 U911 ( .A(n1574), .Y(n2063) );
  AOI22XL U912 ( .A0(n47), .A1(N833), .B0(data[7]), .B1(n632), .Y(n1574) );
  INVX1 U913 ( .A(n1575), .Y(n2066) );
  AOI22XL U914 ( .A0(n637), .A1(N832), .B0(data[6]), .B1(n632), .Y(n1575) );
  INVX1 U915 ( .A(n1576), .Y(n2086) );
  AOI22XL U916 ( .A0(n48), .A1(N831), .B0(data[5]), .B1(n632), .Y(n1576) );
  INVX1 U917 ( .A(n1577), .Y(n2087) );
  AOI22XL U918 ( .A0(n47), .A1(N830), .B0(data[4]), .B1(n632), .Y(n1577) );
  INVX1 U919 ( .A(n1578), .Y(n2088) );
  AOI22XL U920 ( .A0(n47), .A1(N829), .B0(data[3]), .B1(n632), .Y(n1578) );
  INVX1 U921 ( .A(n1579), .Y(n2089) );
  AOI22XL U922 ( .A0(n48), .A1(N828), .B0(data[2]), .B1(n632), .Y(n1579) );
  INVX1 U923 ( .A(n1580), .Y(n2090) );
  AOI22XL U924 ( .A0(n636), .A1(N827), .B0(data[1]), .B1(n632), .Y(n1580) );
  INVX1 U925 ( .A(n1581), .Y(n2222) );
  AOI22XL U926 ( .A0(n636), .A1(N826), .B0(data[0]), .B1(n632), .Y(n1581) );
  INVX1 U927 ( .A(n1485), .Y(n1112) );
  INVX1 U928 ( .A(n1486), .Y(n1149) );
  AOI22XL U929 ( .A0(n645), .A1(N784), .B0(N776), .B1(n642), .Y(n1486) );
  INVX1 U930 ( .A(n1487), .Y(n1265) );
  AOI22XL U931 ( .A0(n644), .A1(N783), .B0(N775), .B1(n642), .Y(n1487) );
  INVX1 U932 ( .A(n1488), .Y(n1272) );
  AOI22XL U933 ( .A0(n49), .A1(N782), .B0(N774), .B1(n642), .Y(n1488) );
  INVX1 U934 ( .A(n1489), .Y(n1300) );
  AOI22XL U935 ( .A0(n646), .A1(N781), .B0(N773), .B1(n642), .Y(n1489) );
  INVX1 U936 ( .A(n1490), .Y(n1704) );
  AOI22XL U937 ( .A0(n645), .A1(N780), .B0(N772), .B1(n641), .Y(n1490) );
  INVX1 U938 ( .A(n1491), .Y(n1705) );
  AOI22XL U939 ( .A0(n644), .A1(N779), .B0(N771), .B1(n1477), .Y(n1491) );
  INVX1 U940 ( .A(n1492), .Y(n1706) );
  AOI22XL U941 ( .A0(n49), .A1(N778), .B0(N770), .B1(n1477), .Y(n1492) );
  INVX1 U942 ( .A(n1493), .Y(n1707) );
  AOI22XL U943 ( .A0(n646), .A1(N777), .B0(N769), .B1(n1477), .Y(n1493) );
  INVX1 U944 ( .A(n1494), .Y(n1708) );
  AOI22XL U945 ( .A0(n645), .A1(N776), .B0(N768), .B1(n1477), .Y(n1494) );
  INVX1 U946 ( .A(n1495), .Y(n1717) );
  AOI22XL U947 ( .A0(n644), .A1(N775), .B0(N767), .B1(n1477), .Y(n1495) );
  INVX1 U948 ( .A(n1496), .Y(n1718) );
  AOI22XL U949 ( .A0(n49), .A1(N774), .B0(N766), .B1(n1477), .Y(n1496) );
  INVX1 U950 ( .A(n1497), .Y(n1719) );
  INVX1 U951 ( .A(n1498), .Y(n1730) );
  AOI22XL U952 ( .A0(n646), .A1(N772), .B0(N764), .B1(n641), .Y(n1498) );
  INVX1 U953 ( .A(n1499), .Y(n1732) );
  AOI22XL U954 ( .A0(n645), .A1(N771), .B0(N763), .B1(n641), .Y(n1499) );
  INVX1 U955 ( .A(n1500), .Y(n1733) );
  AOI22XL U956 ( .A0(n644), .A1(N770), .B0(N762), .B1(n641), .Y(n1500) );
  INVX1 U957 ( .A(n1501), .Y(n1097) );
  AOI22XL U958 ( .A0(n49), .A1(N769), .B0(data[7]), .B1(n641), .Y(n1501) );
  INVX1 U959 ( .A(n1502), .Y(n1098) );
  AOI22XL U960 ( .A0(n646), .A1(N768), .B0(data[6]), .B1(n641), .Y(n1502) );
  INVX1 U961 ( .A(n1503), .Y(n1099) );
  AOI22XL U962 ( .A0(n645), .A1(N767), .B0(data[5]), .B1(n641), .Y(n1503) );
  INVX1 U963 ( .A(n1504), .Y(n1100) );
  AOI22XL U964 ( .A0(n644), .A1(N766), .B0(data[4]), .B1(n641), .Y(n1504) );
  INVX1 U965 ( .A(n1505), .Y(n1101) );
  AOI22XL U966 ( .A0(n49), .A1(N765), .B0(data[3]), .B1(n641), .Y(n1505) );
  INVX1 U967 ( .A(n1506), .Y(n1102) );
  AOI22XL U968 ( .A0(n646), .A1(N764), .B0(data[2]), .B1(n641), .Y(n1506) );
  INVX1 U969 ( .A(n1507), .Y(n1103) );
  AOI22XL U970 ( .A0(n645), .A1(N763), .B0(data[1]), .B1(n641), .Y(n1507) );
  INVX1 U971 ( .A(n1508), .Y(n2223) );
  AOI22XL U972 ( .A0(n644), .A1(N762), .B0(data[0]), .B1(n641), .Y(n1508) );
  AOI22XL U973 ( .A0(n659), .A1(N720), .B0(N712), .B1(n655), .Y(n1417) );
  AOI22XL U974 ( .A0(n659), .A1(N719), .B0(N711), .B1(n655), .Y(n1418) );
  AOI22XL U975 ( .A0(n659), .A1(N718), .B0(N710), .B1(n655), .Y(n1419) );
  AOI22XL U976 ( .A0(n659), .A1(N717), .B0(N709), .B1(n655), .Y(n1420) );
  AOI22XL U977 ( .A0(n659), .A1(N716), .B0(N708), .B1(n655), .Y(n1421) );
  AOI22XL U978 ( .A0(n659), .A1(N715), .B0(N707), .B1(n655), .Y(n1422) );
  AOI22XL U979 ( .A0(n659), .A1(N714), .B0(N706), .B1(n655), .Y(n1423) );
  AOI22XL U980 ( .A0(n659), .A1(N713), .B0(N705), .B1(n655), .Y(n1424) );
  AOI22XL U981 ( .A0(n659), .A1(N712), .B0(N704), .B1(n655), .Y(n1425) );
  AOI22XL U982 ( .A0(n659), .A1(N711), .B0(N703), .B1(n655), .Y(n1426) );
  AOI22XL U983 ( .A0(n659), .A1(N710), .B0(N702), .B1(n655), .Y(n1427) );
  INVX1 U984 ( .A(n1428), .Y(n1062) );
  INVX1 U985 ( .A(n1429), .Y(n1063) );
  AOI22XL U986 ( .A0(n659), .A1(N708), .B0(N700), .B1(n654), .Y(n1429) );
  INVX1 U987 ( .A(n1430), .Y(n1064) );
  AOI22XL U988 ( .A0(n659), .A1(N707), .B0(N699), .B1(n654), .Y(n1430) );
  AOI22XL U989 ( .A0(n659), .A1(N706), .B0(N698), .B1(n654), .Y(n1431) );
  INVX1 U990 ( .A(n1432), .Y(n1030) );
  AOI22XL U991 ( .A0(n660), .A1(N705), .B0(data[7]), .B1(n654), .Y(n1432) );
  INVX1 U992 ( .A(n1433), .Y(n1031) );
  AOI22XL U993 ( .A0(n660), .A1(N704), .B0(data[6]), .B1(n654), .Y(n1433) );
  INVX1 U994 ( .A(n1434), .Y(n1032) );
  AOI22XL U995 ( .A0(n660), .A1(N703), .B0(data[5]), .B1(n654), .Y(n1434) );
  INVX1 U996 ( .A(n1435), .Y(n1033) );
  AOI22XL U997 ( .A0(n660), .A1(N702), .B0(data[4]), .B1(n654), .Y(n1435) );
  INVX1 U998 ( .A(n1436), .Y(n1034) );
  AOI22XL U999 ( .A0(n660), .A1(N701), .B0(data[3]), .B1(n654), .Y(n1436) );
  INVX1 U1000 ( .A(n1437), .Y(n1035) );
  AOI22XL U1001 ( .A0(n660), .A1(N700), .B0(data[2]), .B1(n654), .Y(n1437) );
  INVX1 U1002 ( .A(n1438), .Y(n1036) );
  AOI22XL U1003 ( .A0(n660), .A1(N699), .B0(data[1]), .B1(n654), .Y(n1438) );
  INVX1 U1004 ( .A(n1439), .Y(n2211) );
  AOI22XL U1005 ( .A0(n660), .A1(N698), .B0(data[0]), .B1(n654), .Y(n1439) );
  INVX1 U1006 ( .A(n1344), .Y(n983) );
  AOI22X1 U1007 ( .A0(n666), .A1(N657), .B0(N649), .B1(n55), .Y(n1344) );
  INVX1 U1008 ( .A(n1345), .Y(n984) );
  AOI22X1 U1009 ( .A0(n666), .A1(N656), .B0(N648), .B1(n60), .Y(n1345) );
  INVX1 U1010 ( .A(n1346), .Y(n985) );
  AOI22X1 U1011 ( .A0(n666), .A1(N655), .B0(N647), .B1(n61), .Y(n1346) );
  INVX1 U1012 ( .A(n1347), .Y(n986) );
  AOI22X1 U1013 ( .A0(n666), .A1(N654), .B0(N646), .B1(n55), .Y(n1347) );
  INVX1 U1014 ( .A(n1348), .Y(n987) );
  AOI22X1 U1015 ( .A0(n667), .A1(N653), .B0(N645), .B1(n59), .Y(n1348) );
  INVX1 U1016 ( .A(n1349), .Y(n988) );
  AOI22X1 U1017 ( .A0(n667), .A1(N652), .B0(N644), .B1(n60), .Y(n1349) );
  INVX1 U1018 ( .A(n1350), .Y(n989) );
  AOI22X1 U1019 ( .A0(n667), .A1(N651), .B0(N643), .B1(n59), .Y(n1350) );
  INVX1 U1020 ( .A(n1351), .Y(n990) );
  AOI22X1 U1021 ( .A0(n667), .A1(N650), .B0(N642), .B1(n60), .Y(n1351) );
  INVX1 U1022 ( .A(n1352), .Y(n991) );
  AOI22X1 U1023 ( .A0(n667), .A1(N649), .B0(N641), .B1(n61), .Y(n1352) );
  INVX1 U1024 ( .A(n1353), .Y(n992) );
  AOI22X1 U1025 ( .A0(n667), .A1(N648), .B0(N640), .B1(n59), .Y(n1353) );
  INVX1 U1026 ( .A(n1354), .Y(n993) );
  AOI22X1 U1027 ( .A0(n667), .A1(N647), .B0(N639), .B1(n61), .Y(n1354) );
  INVX1 U1028 ( .A(n1355), .Y(n994) );
  AOI22X1 U1029 ( .A0(n667), .A1(N646), .B0(N638), .B1(n61), .Y(n1355) );
  INVX1 U1030 ( .A(n1356), .Y(n995) );
  AOI22X1 U1031 ( .A0(n667), .A1(N645), .B0(N637), .B1(n61), .Y(n1356) );
  INVX1 U1032 ( .A(n1357), .Y(n996) );
  AOI22X1 U1033 ( .A0(n667), .A1(N644), .B0(N636), .B1(n61), .Y(n1357) );
  INVX1 U1034 ( .A(n1358), .Y(n997) );
  AOI22X1 U1035 ( .A0(n667), .A1(N643), .B0(N635), .B1(n59), .Y(n1358) );
  INVX1 U1036 ( .A(n1359), .Y(n998) );
  AOI22X1 U1037 ( .A0(n667), .A1(N642), .B0(N634), .B1(n60), .Y(n1359) );
  INVX1 U1038 ( .A(n1360), .Y(n968) );
  INVX1 U1039 ( .A(n1361), .Y(n969) );
  INVX1 U1040 ( .A(n1362), .Y(n970) );
  INVX1 U1041 ( .A(n1363), .Y(n971) );
  INVX1 U1042 ( .A(n1364), .Y(n972) );
  INVX1 U1043 ( .A(n1365), .Y(n973) );
  INVX1 U1044 ( .A(n1366), .Y(n974) );
  INVX1 U1045 ( .A(n1367), .Y(n2213) );
  INVX1 U1046 ( .A(n1273), .Y(n921) );
  AOI22X1 U1047 ( .A0(n676), .A1(N593), .B0(N585), .B1(n675), .Y(n1273) );
  INVX1 U1048 ( .A(n1274), .Y(n922) );
  AOI22X1 U1049 ( .A0(n676), .A1(N592), .B0(N584), .B1(n675), .Y(n1274) );
  INVX1 U1050 ( .A(n1275), .Y(n923) );
  AOI22X1 U1051 ( .A0(n676), .A1(N591), .B0(N583), .B1(n675), .Y(n1275) );
  INVX1 U1052 ( .A(n1276), .Y(n924) );
  AOI22X1 U1053 ( .A0(n676), .A1(N590), .B0(N582), .B1(n675), .Y(n1276) );
  INVX1 U1054 ( .A(n1277), .Y(n925) );
  AOI22X1 U1055 ( .A0(n677), .A1(N589), .B0(N581), .B1(n675), .Y(n1277) );
  INVX1 U1056 ( .A(n1278), .Y(n926) );
  AOI22X1 U1057 ( .A0(n677), .A1(N588), .B0(N580), .B1(n675), .Y(n1278) );
  INVX1 U1058 ( .A(n1279), .Y(n927) );
  AOI22X1 U1059 ( .A0(n677), .A1(N587), .B0(N579), .B1(n675), .Y(n1279) );
  INVX1 U1060 ( .A(n1280), .Y(n928) );
  AOI22X1 U1061 ( .A0(n677), .A1(N586), .B0(N578), .B1(n675), .Y(n1280) );
  INVX1 U1062 ( .A(n1281), .Y(n929) );
  AOI22X1 U1063 ( .A0(n677), .A1(N585), .B0(N577), .B1(n675), .Y(n1281) );
  INVX1 U1064 ( .A(n1282), .Y(n930) );
  AOI22X1 U1065 ( .A0(n677), .A1(N584), .B0(N576), .B1(n675), .Y(n1282) );
  INVX1 U1066 ( .A(n1283), .Y(n931) );
  AOI22X1 U1067 ( .A0(n677), .A1(N583), .B0(N575), .B1(n675), .Y(n1283) );
  INVX1 U1068 ( .A(n1284), .Y(n932) );
  AOI22X1 U1069 ( .A0(n677), .A1(N582), .B0(N574), .B1(n675), .Y(n1284) );
  INVX1 U1070 ( .A(n1285), .Y(n933) );
  AOI22X1 U1071 ( .A0(n677), .A1(N581), .B0(N573), .B1(n675), .Y(n1285) );
  INVX1 U1072 ( .A(n1286), .Y(n934) );
  AOI22X1 U1073 ( .A0(n677), .A1(N580), .B0(N572), .B1(n675), .Y(n1286) );
  INVX1 U1074 ( .A(n1287), .Y(n935) );
  AOI22X1 U1075 ( .A0(n677), .A1(N579), .B0(N571), .B1(n675), .Y(n1287) );
  INVX1 U1076 ( .A(n1288), .Y(n936) );
  AOI22X1 U1077 ( .A0(n677), .A1(N578), .B0(N570), .B1(n675), .Y(n1288) );
  INVX1 U1078 ( .A(n1289), .Y(n907) );
  INVX1 U1079 ( .A(n1290), .Y(n908) );
  INVX1 U1080 ( .A(n1291), .Y(n909) );
  INVX1 U1081 ( .A(n1292), .Y(n910) );
  INVX1 U1082 ( .A(n1293), .Y(n911) );
  INVX1 U1083 ( .A(n1294), .Y(n912) );
  INVX1 U1084 ( .A(n1295), .Y(n913) );
  INVX1 U1085 ( .A(n1296), .Y(n2215) );
  INVX1 U1086 ( .A(n1199), .Y(n860) );
  AOI22X1 U1087 ( .A0(n1190), .A1(N529), .B0(N521), .B1(n687), .Y(n1199) );
  INVX1 U1088 ( .A(n1200), .Y(n861) );
  AOI22X1 U1089 ( .A0(n1190), .A1(N528), .B0(N520), .B1(n687), .Y(n1200) );
  INVX1 U1090 ( .A(n1201), .Y(n862) );
  AOI22X1 U1091 ( .A0(n1190), .A1(N527), .B0(N519), .B1(n687), .Y(n1201) );
  INVX1 U1092 ( .A(n1202), .Y(n863) );
  AOI22X1 U1093 ( .A0(n1190), .A1(N526), .B0(N518), .B1(n687), .Y(n1202) );
  INVX1 U1094 ( .A(n1203), .Y(n864) );
  AOI22X1 U1095 ( .A0(n1190), .A1(N525), .B0(N517), .B1(n687), .Y(n1203) );
  INVX1 U1096 ( .A(n1204), .Y(n865) );
  AOI22X1 U1097 ( .A0(n1190), .A1(N524), .B0(N516), .B1(n687), .Y(n1204) );
  INVX1 U1098 ( .A(n1205), .Y(n866) );
  AOI22X1 U1099 ( .A0(n1190), .A1(N523), .B0(N515), .B1(n687), .Y(n1205) );
  INVX1 U1100 ( .A(n1206), .Y(n867) );
  AOI22X1 U1101 ( .A0(n1190), .A1(N522), .B0(N514), .B1(n687), .Y(n1206) );
  INVX1 U1104 ( .A(n1207), .Y(n868) );
  AOI22X1 U1107 ( .A0(n1190), .A1(N521), .B0(N513), .B1(n687), .Y(n1207) );
  INVX1 U1108 ( .A(n1208), .Y(n869) );
  AOI22X1 U1109 ( .A0(n1190), .A1(N520), .B0(N512), .B1(n687), .Y(n1208) );
  INVX1 U1110 ( .A(n1209), .Y(n870) );
  AOI22X1 U1111 ( .A0(n1190), .A1(N519), .B0(N511), .B1(n687), .Y(n1209) );
  INVX1 U1112 ( .A(n1210), .Y(n871) );
  AOI22X1 U1113 ( .A0(n1190), .A1(N518), .B0(N510), .B1(n687), .Y(n1210) );
  INVX1 U1114 ( .A(n1211), .Y(n872) );
  AOI22X1 U1117 ( .A0(n1190), .A1(N517), .B0(N509), .B1(n686), .Y(n1211) );
  INVX1 U1118 ( .A(n1212), .Y(n873) );
  AOI22X1 U1121 ( .A0(n1190), .A1(N516), .B0(N508), .B1(n686), .Y(n1212) );
  INVX1 U1122 ( .A(n1213), .Y(n874) );
  AOI22X1 U1123 ( .A0(n1190), .A1(N515), .B0(N507), .B1(n686), .Y(n1213) );
  INVX1 U1125 ( .A(n1214), .Y(n875) );
  AOI22X1 U1126 ( .A0(n1190), .A1(N514), .B0(N506), .B1(n686), .Y(n1214) );
  INVX1 U1127 ( .A(n1215), .Y(n845) );
  INVX1 U1128 ( .A(n1216), .Y(n846) );
  INVX1 U1130 ( .A(n1217), .Y(n847) );
  INVX1 U1131 ( .A(n1218), .Y(n848) );
  INVX1 U1132 ( .A(n1219), .Y(n849) );
  INVX1 U1133 ( .A(n1220), .Y(n850) );
  INVX1 U1134 ( .A(n1221), .Y(n851) );
  INVX1 U1136 ( .A(n1222), .Y(n2217) );
  INVX1 U1137 ( .A(n1655), .Y(n2184) );
  INVX1 U1138 ( .A(n1658), .Y(n2185) );
  AOI22XL U1139 ( .A0(n613), .A1(buffer[6]), .B0(N944), .B1(n1657), .Y(n1658)
         );
  INVX1 U1140 ( .A(n1659), .Y(n2186) );
  AOI22XL U1141 ( .A0(n613), .A1(buffer[5]), .B0(N943), .B1(n1657), .Y(n1659)
         );
  INVX1 U1142 ( .A(n1660), .Y(n2187) );
  AOI22XL U1143 ( .A0(n613), .A1(buffer[4]), .B0(N942), .B1(n1657), .Y(n1660)
         );
  INVX1 U1144 ( .A(n1661), .Y(n2188) );
  AOI22XL U1145 ( .A0(n613), .A1(buffer[3]), .B0(N941), .B1(n1657), .Y(n1661)
         );
  INVX1 U1146 ( .A(n1662), .Y(n2189) );
  AOI22XL U1147 ( .A0(n613), .A1(buffer[2]), .B0(N940), .B1(n1657), .Y(n1662)
         );
  INVX1 U1148 ( .A(n1663), .Y(n2190) );
  AOI22XL U1149 ( .A0(n613), .A1(buffer[1]), .B0(N939), .B1(n1657), .Y(n1663)
         );
  INVX1 U1150 ( .A(n1664), .Y(n2191) );
  AOI22XL U1151 ( .A0(n613), .A1(buffer[0]), .B0(N938), .B1(n1657), .Y(n1664)
         );
  INVX1 U1152 ( .A(n1619), .Y(n2153) );
  INVX1 U1153 ( .A(n1622), .Y(n2154) );
  AOI22XL U1154 ( .A0(n620), .A1(buffer[14]), .B0(N912), .B1(n4), .Y(n1622) );
  INVX1 U1155 ( .A(n1623), .Y(n2155) );
  AOI22XL U1156 ( .A0(n621), .A1(buffer[13]), .B0(N911), .B1(n11), .Y(n1623)
         );
  INVX1 U1157 ( .A(n1624), .Y(n2156) );
  AOI22XL U1158 ( .A0(n620), .A1(buffer[12]), .B0(N910), .B1(n12), .Y(n1624)
         );
  INVX1 U1159 ( .A(n1625), .Y(n2157) );
  AOI22XL U1160 ( .A0(n621), .A1(buffer[11]), .B0(N909), .B1(n4), .Y(n1625) );
  INVX1 U1161 ( .A(n1626), .Y(n2158) );
  AOI22XL U1162 ( .A0(n620), .A1(buffer[10]), .B0(N908), .B1(n9), .Y(n1626) );
  INVX1 U1163 ( .A(n1627), .Y(n2159) );
  AOI22XL U1164 ( .A0(n621), .A1(buffer[9]), .B0(N907), .B1(n9), .Y(n1627) );
  INVX1 U1165 ( .A(n1628), .Y(n2160) );
  AOI22XL U1166 ( .A0(n620), .A1(buffer[8]), .B0(N906), .B1(n10), .Y(n1628) );
  INVX1 U1167 ( .A(n1584), .Y(n2122) );
  INVX1 U1168 ( .A(n1587), .Y(n2123) );
  AOI22XL U1169 ( .A0(n629), .A1(buffer[22]), .B0(N880), .B1(n625), .Y(n1587)
         );
  INVX1 U1170 ( .A(n1588), .Y(n2124) );
  AOI22XL U1171 ( .A0(n628), .A1(buffer[21]), .B0(N879), .B1(n625), .Y(n1588)
         );
  INVX1 U1172 ( .A(n1589), .Y(n2125) );
  AOI22XL U1173 ( .A0(n628), .A1(buffer[20]), .B0(N878), .B1(n625), .Y(n1589)
         );
  INVX1 U1174 ( .A(n1590), .Y(n2126) );
  AOI22XL U1175 ( .A0(n42), .A1(buffer[19]), .B0(N877), .B1(n625), .Y(n1590)
         );
  INVX1 U1176 ( .A(n1591), .Y(n2127) );
  AOI22XL U1177 ( .A0(n43), .A1(buffer[18]), .B0(N876), .B1(n625), .Y(n1591)
         );
  INVX1 U1178 ( .A(n1592), .Y(n2128) );
  AOI22XL U1179 ( .A0(n629), .A1(buffer[17]), .B0(N875), .B1(n625), .Y(n1592)
         );
  INVX1 U1180 ( .A(n1593), .Y(n2129) );
  AOI22XL U1181 ( .A0(n43), .A1(buffer[16]), .B0(N874), .B1(n625), .Y(n1593)
         );
  INVX1 U1182 ( .A(n1548), .Y(n2091) );
  INVX1 U1183 ( .A(n1551), .Y(n2092) );
  AOI22XL U1184 ( .A0(n636), .A1(buffer[30]), .B0(N848), .B1(n633), .Y(n1551)
         );
  INVX1 U1185 ( .A(n1552), .Y(n2093) );
  AOI22XL U1186 ( .A0(n47), .A1(buffer[29]), .B0(N847), .B1(n633), .Y(n1552)
         );
  INVX1 U1187 ( .A(n1553), .Y(n2094) );
  AOI22XL U1188 ( .A0(n47), .A1(buffer[28]), .B0(N846), .B1(n633), .Y(n1553)
         );
  INVX1 U1189 ( .A(n1554), .Y(n2095) );
  AOI22XL U1190 ( .A0(n48), .A1(buffer[27]), .B0(N845), .B1(n633), .Y(n1554)
         );
  INVX1 U1191 ( .A(n1555), .Y(n2096) );
  AOI22XL U1192 ( .A0(n637), .A1(buffer[26]), .B0(N844), .B1(n633), .Y(n1555)
         );
  INVX1 U1193 ( .A(n1556), .Y(n2097) );
  AOI22XL U1194 ( .A0(n637), .A1(buffer[25]), .B0(N843), .B1(n633), .Y(n1556)
         );
  INVX1 U1195 ( .A(n1557), .Y(n2098) );
  AOI22XL U1196 ( .A0(n48), .A1(buffer[24]), .B0(N842), .B1(n633), .Y(n1557)
         );
  INVX1 U1197 ( .A(n1511), .Y(n1799) );
  INVX1 U1198 ( .A(n1514), .Y(n1810) );
  AOI22XL U1199 ( .A0(n38), .A1(buffer[38]), .B0(N816), .B1(n639), .Y(n1514)
         );
  INVX1 U1200 ( .A(n1515), .Y(n1821) );
  AOI22XL U1201 ( .A0(n40), .A1(buffer[37]), .B0(N815), .B1(n639), .Y(n1515)
         );
  INVX1 U1202 ( .A(n1516), .Y(n1832) );
  AOI22XL U1203 ( .A0(n38), .A1(buffer[36]), .B0(N814), .B1(n639), .Y(n1516)
         );
  INVX1 U1204 ( .A(n1517), .Y(n1843) );
  AOI22XL U1205 ( .A0(n41), .A1(buffer[35]), .B0(N813), .B1(n639), .Y(n1517)
         );
  INVX1 U1206 ( .A(n1518), .Y(n1854) );
  AOI22XL U1207 ( .A0(n36), .A1(buffer[34]), .B0(N812), .B1(n639), .Y(n1518)
         );
  INVX1 U1208 ( .A(n1519), .Y(n1865) );
  AOI22XL U1209 ( .A0(n38), .A1(buffer[33]), .B0(N811), .B1(n639), .Y(n1519)
         );
  INVX1 U1210 ( .A(n1520), .Y(n1876) );
  AOI22XL U1211 ( .A0(n40), .A1(buffer[32]), .B0(N810), .B1(n639), .Y(n1520)
         );
  INVX1 U1212 ( .A(n1475), .Y(n1104) );
  INVX1 U1213 ( .A(n1478), .Y(n1105) );
  AOI22XL U1214 ( .A0(n646), .A1(buffer[46]), .B0(N784), .B1(n642), .Y(n1478)
         );
  INVX1 U1215 ( .A(n1479), .Y(n1106) );
  AOI22XL U1216 ( .A0(n645), .A1(buffer[45]), .B0(N783), .B1(n642), .Y(n1479)
         );
  INVX1 U1217 ( .A(n1480), .Y(n1107) );
  AOI22XL U1218 ( .A0(n644), .A1(buffer[44]), .B0(N782), .B1(n642), .Y(n1480)
         );
  INVX1 U1219 ( .A(n1481), .Y(n1108) );
  AOI22XL U1220 ( .A0(n49), .A1(buffer[43]), .B0(N781), .B1(n642), .Y(n1481)
         );
  INVX1 U1221 ( .A(n1482), .Y(n1109) );
  AOI22XL U1222 ( .A0(n646), .A1(buffer[42]), .B0(N780), .B1(n642), .Y(n1482)
         );
  INVX1 U1223 ( .A(n1483), .Y(n1110) );
  AOI22XL U1224 ( .A0(n645), .A1(buffer[41]), .B0(N779), .B1(n642), .Y(n1483)
         );
  INVX1 U1225 ( .A(n1484), .Y(n1111) );
  AOI22XL U1226 ( .A0(n644), .A1(buffer[40]), .B0(N778), .B1(n642), .Y(n1484)
         );
  INVX1 U1227 ( .A(n1441), .Y(n1073) );
  INVX1 U1228 ( .A(n1444), .Y(n1074) );
  AOI22XL U1229 ( .A0(n651), .A1(buffer[54]), .B0(N752), .B1(n649), .Y(n1444)
         );
  INVX1 U1230 ( .A(n1445), .Y(n1075) );
  AOI22XL U1231 ( .A0(n651), .A1(buffer[53]), .B0(N751), .B1(n649), .Y(n1445)
         );
  INVX1 U1232 ( .A(n1446), .Y(n1076) );
  AOI22XL U1233 ( .A0(n651), .A1(buffer[52]), .B0(N750), .B1(n649), .Y(n1446)
         );
  INVX1 U1234 ( .A(n1447), .Y(n1077) );
  AOI22XL U1235 ( .A0(n651), .A1(buffer[51]), .B0(N749), .B1(n649), .Y(n1447)
         );
  INVX1 U1236 ( .A(n1448), .Y(n1078) );
  AOI22XL U1237 ( .A0(n651), .A1(buffer[50]), .B0(N748), .B1(n649), .Y(n1448)
         );
  INVX1 U1238 ( .A(n1449), .Y(n1079) );
  AOI22XL U1239 ( .A0(n651), .A1(buffer[49]), .B0(N747), .B1(n649), .Y(n1449)
         );
  INVX1 U1240 ( .A(n1450), .Y(n1080) );
  AOI22XL U1241 ( .A0(n651), .A1(buffer[48]), .B0(N746), .B1(n649), .Y(n1450)
         );
  INVX1 U1242 ( .A(n1406), .Y(n1037) );
  INVX1 U1243 ( .A(n1409), .Y(n1038) );
  AOI22XL U1244 ( .A0(n659), .A1(buffer[62]), .B0(N720), .B1(n656), .Y(n1409)
         );
  INVX1 U1245 ( .A(n1410), .Y(n1039) );
  AOI22XL U1246 ( .A0(n659), .A1(buffer[61]), .B0(N719), .B1(n656), .Y(n1410)
         );
  INVX1 U1247 ( .A(n1411), .Y(n1040) );
  AOI22XL U1248 ( .A0(n659), .A1(buffer[60]), .B0(N718), .B1(n656), .Y(n1411)
         );
  INVX1 U1249 ( .A(n1412), .Y(n1041) );
  AOI22XL U1250 ( .A0(n659), .A1(buffer[59]), .B0(N717), .B1(n656), .Y(n1412)
         );
  INVX1 U1251 ( .A(n1413), .Y(n1042) );
  AOI22XL U1252 ( .A0(n659), .A1(buffer[58]), .B0(N716), .B1(n656), .Y(n1413)
         );
  INVX1 U1253 ( .A(n1414), .Y(n1043) );
  AOI22XL U1254 ( .A0(n659), .A1(buffer[57]), .B0(N715), .B1(n656), .Y(n1414)
         );
  INVX1 U1255 ( .A(n1415), .Y(n1044) );
  AOI22XL U1256 ( .A0(n659), .A1(buffer[56]), .B0(N714), .B1(n656), .Y(n1415)
         );
  INVX1 U1257 ( .A(n1370), .Y(n1006) );
  AOI22X1 U1258 ( .A0(n662), .A1(buffer[71]), .B0(N689), .B1(n51), .Y(n1370)
         );
  INVX1 U1259 ( .A(n1373), .Y(n1007) );
  AOI22X1 U1260 ( .A0(n662), .A1(buffer[70]), .B0(N688), .B1(n54), .Y(n1373)
         );
  INVX1 U1261 ( .A(n1374), .Y(n1008) );
  AOI22X1 U1262 ( .A0(n662), .A1(buffer[69]), .B0(N687), .B1(n51), .Y(n1374)
         );
  INVX1 U1263 ( .A(n1375), .Y(n1009) );
  AOI22X1 U1264 ( .A0(n662), .A1(buffer[68]), .B0(N686), .B1(n53), .Y(n1375)
         );
  INVX1 U1265 ( .A(n1376), .Y(n1010) );
  AOI22X1 U1266 ( .A0(n662), .A1(buffer[67]), .B0(N685), .B1(n53), .Y(n1376)
         );
  INVX1 U1267 ( .A(n1377), .Y(n1011) );
  AOI22X1 U1268 ( .A0(n662), .A1(buffer[66]), .B0(N684), .B1(n54), .Y(n1377)
         );
  INVX1 U1269 ( .A(n1378), .Y(n1012) );
  AOI22X1 U1270 ( .A0(n662), .A1(buffer[65]), .B0(N683), .B1(n53), .Y(n1378)
         );
  INVX1 U1271 ( .A(n1379), .Y(n1013) );
  AOI22X1 U1272 ( .A0(n662), .A1(buffer[64]), .B0(N682), .B1(n51), .Y(n1379)
         );
  INVX1 U1273 ( .A(n1334), .Y(n975) );
  AOI22X1 U1274 ( .A0(n666), .A1(buffer[79]), .B0(N657), .B1(n55), .Y(n1334)
         );
  INVX1 U1275 ( .A(n1337), .Y(n976) );
  AOI22X1 U1276 ( .A0(n666), .A1(buffer[78]), .B0(N656), .B1(n59), .Y(n1337)
         );
  INVX1 U1277 ( .A(n1338), .Y(n977) );
  AOI22X1 U1278 ( .A0(n666), .A1(buffer[77]), .B0(N655), .B1(n55), .Y(n1338)
         );
  INVX1 U1279 ( .A(n1339), .Y(n978) );
  AOI22X1 U1280 ( .A0(n666), .A1(buffer[76]), .B0(N654), .B1(n59), .Y(n1339)
         );
  INVX1 U1281 ( .A(n1340), .Y(n979) );
  AOI22X1 U1282 ( .A0(n666), .A1(buffer[75]), .B0(N653), .B1(n60), .Y(n1340)
         );
  INVX1 U1283 ( .A(n1341), .Y(n980) );
  AOI22X1 U1284 ( .A0(n666), .A1(buffer[74]), .B0(N652), .B1(n61), .Y(n1341)
         );
  INVX1 U1285 ( .A(n1342), .Y(n981) );
  AOI22X1 U1286 ( .A0(n666), .A1(buffer[73]), .B0(N651), .B1(n59), .Y(n1342)
         );
  INVX1 U1287 ( .A(n1343), .Y(n982) );
  AOI22X1 U1288 ( .A0(n666), .A1(buffer[72]), .B0(N650), .B1(n60), .Y(n1343)
         );
  INVX1 U1289 ( .A(n1298), .Y(n944) );
  AOI22X1 U1290 ( .A0(n670), .A1(buffer[87]), .B0(N625), .B1(n45), .Y(n1298)
         );
  INVX1 U1291 ( .A(n1301), .Y(n945) );
  AOI22X1 U1292 ( .A0(n670), .A1(buffer[86]), .B0(N624), .B1(n44), .Y(n1301)
         );
  INVX1 U1293 ( .A(n1302), .Y(n946) );
  AOI22X1 U1294 ( .A0(n670), .A1(buffer[85]), .B0(N623), .B1(n44), .Y(n1302)
         );
  INVX1 U1295 ( .A(n1303), .Y(n947) );
  AOI22X1 U1296 ( .A0(n670), .A1(buffer[84]), .B0(N622), .B1(n45), .Y(n1303)
         );
  INVX1 U1297 ( .A(n1304), .Y(n948) );
  AOI22X1 U1298 ( .A0(n670), .A1(buffer[83]), .B0(N621), .B1(n44), .Y(n1304)
         );
  INVX1 U1299 ( .A(n1305), .Y(n949) );
  AOI22X1 U1300 ( .A0(n670), .A1(buffer[82]), .B0(N620), .B1(n45), .Y(n1305)
         );
  INVX1 U1301 ( .A(n1306), .Y(n950) );
  AOI22X1 U1302 ( .A0(n670), .A1(buffer[81]), .B0(N619), .B1(n44), .Y(n1306)
         );
  INVX1 U1303 ( .A(n1307), .Y(n951) );
  AOI22X1 U1304 ( .A0(n670), .A1(buffer[80]), .B0(N618), .B1(n46), .Y(n1307)
         );
  INVX1 U1305 ( .A(n1263), .Y(n914) );
  AOI22X1 U1306 ( .A0(n676), .A1(buffer[95]), .B0(N593), .B1(n675), .Y(n1263)
         );
  INVX1 U1307 ( .A(n1266), .Y(n915) );
  AOI22X1 U1308 ( .A0(n676), .A1(buffer[94]), .B0(N592), .B1(n675), .Y(n1266)
         );
  INVX1 U1309 ( .A(n1267), .Y(n916) );
  AOI22X1 U1310 ( .A0(n676), .A1(buffer[93]), .B0(N591), .B1(n675), .Y(n1267)
         );
  INVX1 U1311 ( .A(n1268), .Y(n917) );
  AOI22X1 U1312 ( .A0(n676), .A1(buffer[92]), .B0(N590), .B1(n675), .Y(n1268)
         );
  INVX1 U1313 ( .A(n1269), .Y(n918) );
  AOI22X1 U1314 ( .A0(n676), .A1(buffer[91]), .B0(N589), .B1(n675), .Y(n1269)
         );
  INVX1 U1315 ( .A(n1270), .Y(n919) );
  AOI22X1 U1316 ( .A0(n676), .A1(buffer[90]), .B0(N588), .B1(n675), .Y(n1270)
         );
  INVX1 U1317 ( .A(n1271), .Y(n920) );
  AOI22X1 U1318 ( .A0(n676), .A1(buffer[89]), .B0(N587), .B1(n675), .Y(n1271)
         );
  INVX1 U1319 ( .A(n1225), .Y(n883) );
  AOI22X1 U1320 ( .A0(n684), .A1(buffer[103]), .B0(N561), .B1(n680), .Y(n1225)
         );
  INVX1 U1321 ( .A(n1228), .Y(n884) );
  AOI22X1 U1322 ( .A0(n684), .A1(buffer[102]), .B0(N560), .B1(n680), .Y(n1228)
         );
  INVX1 U1323 ( .A(n1229), .Y(n885) );
  AOI22X1 U1324 ( .A0(n684), .A1(buffer[101]), .B0(N559), .B1(n680), .Y(n1229)
         );
  INVX1 U1325 ( .A(n1230), .Y(n886) );
  AOI22X1 U1326 ( .A0(n684), .A1(buffer[100]), .B0(N558), .B1(n680), .Y(n1230)
         );
  INVX1 U1327 ( .A(n1231), .Y(n887) );
  AOI22X1 U1328 ( .A0(n684), .A1(buffer[99]), .B0(N557), .B1(n680), .Y(n1231)
         );
  INVX1 U1329 ( .A(n1232), .Y(n888) );
  AOI22X1 U1330 ( .A0(n684), .A1(buffer[98]), .B0(N556), .B1(n680), .Y(n1232)
         );
  INVX1 U1331 ( .A(n1233), .Y(n889) );
  AOI22X1 U1332 ( .A0(n684), .A1(buffer[97]), .B0(N555), .B1(n680), .Y(n1233)
         );
  INVX1 U1333 ( .A(n1234), .Y(n890) );
  AOI22X1 U1334 ( .A0(n684), .A1(buffer[96]), .B0(N554), .B1(n680), .Y(n1234)
         );
  INVX1 U1335 ( .A(n1189), .Y(n852) );
  AOI22X1 U1336 ( .A0(n1190), .A1(buffer[111]), .B0(N529), .B1(n687), .Y(n1189) );
  INVX1 U1337 ( .A(n1192), .Y(n853) );
  AOI22X1 U1338 ( .A0(n1190), .A1(buffer[110]), .B0(N528), .B1(n687), .Y(n1192) );
  INVX1 U1339 ( .A(n1193), .Y(n854) );
  AOI22X1 U1340 ( .A0(n1190), .A1(buffer[109]), .B0(N527), .B1(n687), .Y(n1193) );
  INVX1 U1341 ( .A(n1194), .Y(n855) );
  AOI22X1 U1342 ( .A0(n1190), .A1(buffer[108]), .B0(N526), .B1(n687), .Y(n1194) );
  INVX1 U1343 ( .A(n1195), .Y(n856) );
  AOI22X1 U1344 ( .A0(n1190), .A1(buffer[107]), .B0(N525), .B1(n687), .Y(n1195) );
  INVX1 U1345 ( .A(n1196), .Y(n857) );
  AOI22X1 U1346 ( .A0(n1190), .A1(buffer[106]), .B0(N524), .B1(n687), .Y(n1196) );
  INVX1 U1347 ( .A(n1197), .Y(n858) );
  AOI22X1 U1348 ( .A0(n1190), .A1(buffer[105]), .B0(N523), .B1(n687), .Y(n1197) );
  INVX1 U1349 ( .A(n1198), .Y(n859) );
  AOI22X1 U1350 ( .A0(n1190), .A1(buffer[104]), .B0(N522), .B1(n687), .Y(n1198) );
  AND3X1 U1351 ( .A(n1691), .B(n1261), .C(write_enable), .Y(n1697) );
  AOI2BB1X1 U1352 ( .A0N(n1147), .A1N(n1148), .B0(reset), .Y(n1114) );
  NAND4X1 U1353 ( .A(n29), .B(n1150), .C(n1151), .D(n1152), .Y(n1148) );
  NAND4XL U1354 ( .A(write_enable), .B(n1153), .C(n1154), .D(n1155), .Y(n1147)
         );
  INVX1 U1355 ( .A(n1166), .Y(n829) );
  AOI22X1 U1356 ( .A0(n695), .A1(N497), .B0(N489), .B1(n691), .Y(n1166) );
  INVX1 U1357 ( .A(n1167), .Y(n830) );
  AOI22X1 U1358 ( .A0(n695), .A1(N496), .B0(N488), .B1(n691), .Y(n1167) );
  INVX1 U1359 ( .A(n1168), .Y(n831) );
  AOI22X1 U1360 ( .A0(n695), .A1(N495), .B0(N487), .B1(n691), .Y(n1168) );
  INVX1 U1361 ( .A(n1169), .Y(n832) );
  AOI22X1 U1362 ( .A0(n695), .A1(N494), .B0(N486), .B1(n691), .Y(n1169) );
  INVX1 U1363 ( .A(n1170), .Y(n833) );
  AOI22X1 U1364 ( .A0(n696), .A1(N493), .B0(N485), .B1(n691), .Y(n1170) );
  INVX1 U1365 ( .A(n1171), .Y(n834) );
  AOI22X1 U1366 ( .A0(n696), .A1(N492), .B0(N484), .B1(n691), .Y(n1171) );
  INVX1 U1367 ( .A(n1172), .Y(n835) );
  AOI22X1 U1368 ( .A0(n696), .A1(N491), .B0(N483), .B1(n691), .Y(n1172) );
  INVX1 U1369 ( .A(n1173), .Y(n836) );
  AOI22X1 U1370 ( .A0(n696), .A1(N490), .B0(N482), .B1(n691), .Y(n1173) );
  INVX1 U1371 ( .A(n1174), .Y(n837) );
  AOI22X1 U1372 ( .A0(n696), .A1(N489), .B0(N481), .B1(n691), .Y(n1174) );
  INVX1 U1373 ( .A(n1175), .Y(n838) );
  AOI22X1 U1374 ( .A0(n696), .A1(N488), .B0(N480), .B1(n691), .Y(n1175) );
  INVX1 U1375 ( .A(n1176), .Y(n839) );
  AOI22X1 U1376 ( .A0(n696), .A1(N487), .B0(N479), .B1(n691), .Y(n1176) );
  AOI22X1 U1377 ( .A0(n696), .A1(N486), .B0(N478), .B1(n691), .Y(n1177) );
  INVX1 U1378 ( .A(n1178), .Y(n841) );
  AOI22X1 U1379 ( .A0(n696), .A1(N485), .B0(N477), .B1(n690), .Y(n1178) );
  INVX1 U1380 ( .A(n1179), .Y(n842) );
  AOI22X1 U1381 ( .A0(n696), .A1(N484), .B0(N476), .B1(n690), .Y(n1179) );
  INVX1 U1382 ( .A(n1180), .Y(n843) );
  AOI22X1 U1383 ( .A0(n696), .A1(N483), .B0(N475), .B1(n690), .Y(n1180) );
  INVX1 U1384 ( .A(n1181), .Y(n844) );
  AOI22X1 U1385 ( .A0(n696), .A1(N482), .B0(N474), .B1(n690), .Y(n1181) );
  INVX1 U1386 ( .A(n1182), .Y(n814) );
  INVX1 U1387 ( .A(n1183), .Y(n815) );
  INVX1 U1388 ( .A(n1184), .Y(n816) );
  INVX1 U1389 ( .A(n1185), .Y(n817) );
  INVX1 U1390 ( .A(n1186), .Y(n818) );
  INVX1 U1391 ( .A(n1187), .Y(n819) );
  INVX1 U1392 ( .A(n1188), .Y(n820) );
  INVX1 U1393 ( .A(n1123), .Y(n798) );
  AOI22X1 U1394 ( .A0(n704), .A1(N465), .B0(N457), .B1(n700), .Y(n1123) );
  INVX1 U1395 ( .A(n1124), .Y(n799) );
  AOI22X1 U1396 ( .A0(n704), .A1(N464), .B0(N456), .B1(n700), .Y(n1124) );
  INVX1 U1397 ( .A(n1125), .Y(n800) );
  AOI22X1 U1398 ( .A0(n704), .A1(N463), .B0(N455), .B1(n700), .Y(n1125) );
  INVX1 U1399 ( .A(n1126), .Y(n801) );
  AOI22X1 U1400 ( .A0(n704), .A1(N462), .B0(N454), .B1(n700), .Y(n1126) );
  INVX1 U1401 ( .A(n1127), .Y(n802) );
  AOI22X1 U1402 ( .A0(n705), .A1(N461), .B0(N453), .B1(n700), .Y(n1127) );
  INVX1 U1403 ( .A(n1128), .Y(n803) );
  AOI22X1 U1404 ( .A0(n705), .A1(N460), .B0(N452), .B1(n700), .Y(n1128) );
  INVX1 U1405 ( .A(n1129), .Y(n804) );
  AOI22X1 U1406 ( .A0(n705), .A1(N459), .B0(N451), .B1(n700), .Y(n1129) );
  INVX1 U1407 ( .A(n1130), .Y(n805) );
  AOI22X1 U1408 ( .A0(n705), .A1(N458), .B0(N450), .B1(n700), .Y(n1130) );
  INVX1 U1409 ( .A(n1131), .Y(n806) );
  AOI22X1 U1410 ( .A0(n705), .A1(N457), .B0(N449), .B1(n700), .Y(n1131) );
  INVX1 U1411 ( .A(n1132), .Y(n807) );
  AOI22X1 U1412 ( .A0(n705), .A1(N456), .B0(N448), .B1(n700), .Y(n1132) );
  INVX1 U1413 ( .A(n1133), .Y(n808) );
  AOI22X1 U1414 ( .A0(n705), .A1(N455), .B0(N447), .B1(n700), .Y(n1133) );
  INVX1 U1415 ( .A(n1134), .Y(n809) );
  AOI22X1 U1416 ( .A0(n705), .A1(N454), .B0(N446), .B1(n700), .Y(n1134) );
  INVX1 U1417 ( .A(n1135), .Y(n810) );
  INVX1 U1418 ( .A(n1136), .Y(n811) );
  AOI22X1 U1419 ( .A0(n705), .A1(N452), .B0(N444), .B1(n699), .Y(n1136) );
  INVX1 U1420 ( .A(n1137), .Y(n812) );
  AOI22X1 U1421 ( .A0(n705), .A1(N451), .B0(N443), .B1(n699), .Y(n1137) );
  INVX1 U1422 ( .A(n1138), .Y(n813) );
  AOI22X1 U1423 ( .A0(n705), .A1(N450), .B0(N442), .B1(n699), .Y(n1138) );
  INVX1 U1424 ( .A(n1139), .Y(n783) );
  INVX1 U1425 ( .A(n1140), .Y(n784) );
  INVX1 U1426 ( .A(n1141), .Y(n785) );
  INVX1 U1427 ( .A(n1142), .Y(n786) );
  INVX1 U1428 ( .A(n1143), .Y(n787) );
  INVX1 U1429 ( .A(n1144), .Y(n788) );
  INVX1 U1430 ( .A(n1145), .Y(n789) );
  INVX1 U1431 ( .A(n1146), .Y(n2218) );
  INVX1 U1432 ( .A(n1156), .Y(n821) );
  AOI22X1 U1433 ( .A0(n695), .A1(buffer[119]), .B0(N497), .B1(n692), .Y(n1156)
         );
  INVX1 U1434 ( .A(n1159), .Y(n822) );
  AOI22X1 U1435 ( .A0(n695), .A1(buffer[118]), .B0(N496), .B1(n692), .Y(n1159)
         );
  INVX1 U1436 ( .A(n1160), .Y(n823) );
  AOI22X1 U1437 ( .A0(n695), .A1(buffer[117]), .B0(N495), .B1(n692), .Y(n1160)
         );
  INVX1 U1438 ( .A(n1161), .Y(n824) );
  AOI22X1 U1439 ( .A0(n695), .A1(buffer[116]), .B0(N494), .B1(n692), .Y(n1161)
         );
  INVX1 U1440 ( .A(n1162), .Y(n825) );
  AOI22X1 U1441 ( .A0(n695), .A1(buffer[115]), .B0(N493), .B1(n692), .Y(n1162)
         );
  INVX1 U1442 ( .A(n1163), .Y(n826) );
  AOI22X1 U1443 ( .A0(n695), .A1(buffer[114]), .B0(N492), .B1(n692), .Y(n1163)
         );
  INVX1 U1444 ( .A(n1164), .Y(n827) );
  AOI22X1 U1445 ( .A0(n695), .A1(buffer[113]), .B0(N491), .B1(n692), .Y(n1164)
         );
  INVX1 U1446 ( .A(n1165), .Y(n828) );
  AOI22X1 U1447 ( .A0(n695), .A1(buffer[112]), .B0(N490), .B1(n692), .Y(n1165)
         );
  INVX1 U1448 ( .A(n1113), .Y(n790) );
  AOI22X1 U1449 ( .A0(n704), .A1(buffer[127]), .B0(N465), .B1(n701), .Y(n1113)
         );
  INVX1 U1450 ( .A(n1116), .Y(n791) );
  AOI22X1 U1451 ( .A0(n704), .A1(buffer[126]), .B0(N464), .B1(n701), .Y(n1116)
         );
  INVX1 U1452 ( .A(n1117), .Y(n792) );
  AOI22X1 U1453 ( .A0(n704), .A1(buffer[125]), .B0(N463), .B1(n701), .Y(n1117)
         );
  INVX1 U1454 ( .A(n1118), .Y(n793) );
  AOI22X1 U1455 ( .A0(n704), .A1(buffer[124]), .B0(N462), .B1(n701), .Y(n1118)
         );
  INVX1 U1456 ( .A(n1119), .Y(n794) );
  AOI22X1 U1457 ( .A0(n704), .A1(buffer[123]), .B0(N461), .B1(n701), .Y(n1119)
         );
  INVX1 U1458 ( .A(n1120), .Y(n795) );
  AOI22X1 U1459 ( .A0(n704), .A1(buffer[122]), .B0(N460), .B1(n701), .Y(n1120)
         );
  INVX1 U1460 ( .A(n1121), .Y(n796) );
  AOI22X1 U1461 ( .A0(n704), .A1(buffer[121]), .B0(N459), .B1(n701), .Y(n1121)
         );
  INVX1 U1462 ( .A(n1122), .Y(n797) );
  AOI22X1 U1463 ( .A0(n704), .A1(buffer[120]), .B0(N458), .B1(n701), .Y(n1122)
         );
  NOR2BX1 U1464 ( .AN(write_enable), .B(reset), .Y(n2085) );
  NAND4BBX1 U1465 ( .AN(counter2[4]), .BN(counter2[5]), .C(counter2[6]), .D(
        n1720), .Y(n2084) );
  XOR3X2 U1466 ( .A(R14[18]), .B(R14[7]), .C(R14[3]), .Y(sigma0[0]) );
  XOR3X2 U1467 ( .A(R1[19]), .B(R1[17]), .C(R1[10]), .Y(sigma1[0]) );
  XOR3X2 U1468 ( .A(R14[27]), .B(R14[16]), .C(R14[12]), .Y(sigma0[9]) );
  XOR3X2 U1469 ( .A(R14[20]), .B(R14[9]), .C(R14[5]), .Y(sigma0[2]) );
  XOR3X2 U1470 ( .A(R14[19]), .B(R14[8]), .C(R14[4]), .Y(sigma0[1]) );
  XOR3X2 U1471 ( .A(R14[23]), .B(R14[12]), .C(R14[8]), .Y(sigma0[5]) );
  XOR3X2 U1472 ( .A(R14[25]), .B(R14[14]), .C(R14[10]), .Y(sigma0[7]) );
  XOR3X2 U1473 ( .A(R14[24]), .B(R14[13]), .C(R14[9]), .Y(sigma0[6]) );
  XOR3X2 U1474 ( .A(R14[22]), .B(R14[11]), .C(R14[7]), .Y(sigma0[4]) );
  XOR3X2 U1475 ( .A(R1[20]), .B(R1[18]), .C(R1[11]), .Y(sigma1[1]) );
  XOR3X2 U1476 ( .A(R1[22]), .B(R1[24]), .C(R1[15]), .Y(sigma1[5]) );
  XOR3X2 U1477 ( .A(R1[24]), .B(R1[26]), .C(R1[17]), .Y(sigma1[7]) );
  XOR3X2 U1478 ( .A(R1[26]), .B(R1[28]), .C(R1[19]), .Y(sigma1[9]) );
  XOR3X2 U1479 ( .A(R1[23]), .B(R1[25]), .C(R1[16]), .Y(sigma1[6]) );
  XOR3X2 U1480 ( .A(R1[21]), .B(R1[23]), .C(R1[14]), .Y(sigma1[4]) );
  XOR3X2 U1481 ( .A(R14[18]), .B(R14[29]), .C(R14[14]), .Y(sigma0[11]) );
  XOR3X2 U1482 ( .A(R14[19]), .B(R14[30]), .C(R14[15]), .Y(sigma0[12]) );
  XOR3X2 U1483 ( .A(R14[20]), .B(R14[31]), .C(R14[16]), .Y(sigma0[13]) );
  XOR3X2 U1484 ( .A(R14[21]), .B(R14[17]), .C(R14[0]), .Y(sigma0[14]) );
  XOR3X2 U1485 ( .A(R14[28]), .B(R14[17]), .C(R14[13]), .Y(sigma0[10]) );
  XOR3X2 U1486 ( .A(R14[26]), .B(R14[15]), .C(R14[11]), .Y(sigma0[8]) );
  XOR3X2 U1487 ( .A(R1[25]), .B(R1[2]), .C(R1[0]), .Y(sigma1[15]) );
  XOR3X2 U1488 ( .A(R1[26]), .B(R1[3]), .C(R1[1]), .Y(sigma1[16]) );
  XOR3X2 U1489 ( .A(R14[18]), .B(R14[22]), .C(R14[1]), .Y(sigma0[15]) );
  XOR3X2 U1490 ( .A(R14[20]), .B(R14[24]), .C(R14[3]), .Y(sigma0[17]) );
  XOR3X2 U1491 ( .A(R14[21]), .B(R14[25]), .C(R14[4]), .Y(sigma0[18]) );
  XOR3X2 U1492 ( .A(R14[22]), .B(R14[26]), .C(R14[5]), .Y(sigma0[19]) );
  XOR3X2 U1493 ( .A(R1[28]), .B(R1[30]), .C(R1[21]), .Y(sigma1[11]) );
  XOR3X2 U1494 ( .A(R1[24]), .B(R1[31]), .C(R1[1]), .Y(sigma1[14]) );
  XOR3X2 U1495 ( .A(R1[29]), .B(R1[31]), .C(R1[22]), .Y(sigma1[12]) );
  XOR3X2 U1496 ( .A(R1[23]), .B(R1[30]), .C(R1[0]), .Y(sigma1[13]) );
  XOR3X2 U1497 ( .A(R1[25]), .B(R1[27]), .C(R1[18]), .Y(sigma1[8]) );
  XOR3X2 U1498 ( .A(R1[27]), .B(R1[29]), .C(R1[20]), .Y(sigma1[10]) );
  XOR3X2 U1499 ( .A(R1[27]), .B(R1[4]), .C(R1[2]), .Y(sigma1[17]) );
  XOR3X2 U1500 ( .A(R1[28]), .B(R1[5]), .C(R1[3]), .Y(sigma1[18]) );
  XOR3X2 U1501 ( .A(R1[29]), .B(R1[6]), .C(R1[4]), .Y(sigma1[19]) );
  NOR2X1 U1502 ( .A(counter1[4]), .B(counter1[5]), .Y(n1692) );
  NOR2X1 U1503 ( .A(counter1[2]), .B(counter1[3]), .Y(n1699) );
  NOR2X1 U1504 ( .A(n1057), .B(counter1[3]), .Y(n1693) );
  NOR2BX1 U1505 ( .AN(counter1[3]), .B(counter1[2]), .Y(n1702) );
  NOR2BX1 U1506 ( .AN(counter1[3]), .B(n1057), .Y(n1700) );
  XOR3X2 U1507 ( .A(R14[25]), .B(R14[29]), .C(R14[8]), .Y(sigma0[22]) );
  XOR3X2 U1508 ( .A(R14[26]), .B(R14[30]), .C(R14[9]), .Y(sigma0[23]) );
  XOR3X2 U1509 ( .A(R14[24]), .B(R14[28]), .C(R14[7]), .Y(sigma0[21]) );
  XOR3X2 U1510 ( .A(R14[19]), .B(R14[23]), .C(R14[2]), .Y(sigma0[16]) );
  XOR3X2 U1511 ( .A(R14[23]), .B(R14[27]), .C(R14[6]), .Y(sigma0[20]) );
  XOR3X2 U1512 ( .A(R1[30]), .B(R1[7]), .C(R1[5]), .Y(sigma1[20]) );
  XOR3X2 U1513 ( .A(R1[31]), .B(R1[8]), .C(R1[6]), .Y(sigma1[21]) );
  XOR2X1 U1514 ( .A(R1[7]), .B(R1[9]), .Y(sigma1[22]) );
  NOR3X1 U1515 ( .A(n1653), .B(counter1[6]), .C(n1689), .Y(n1546) );
  NOR2X1 U1516 ( .A(n1056), .B(counter1[4]), .Y(n1701) );
  NOR2BX1 U1517 ( .AN(counter1[4]), .B(counter1[5]), .Y(n1698) );
  NOR2BX1 U1518 ( .AN(counter1[4]), .B(n1056), .Y(n1703) );
  NOR2X1 U1519 ( .A(counter2[2]), .B(counter2[1]), .Y(n2077) );
  XOR3X2 U1520 ( .A(R14[27]), .B(R14[31]), .C(R14[10]), .Y(sigma0[24]) );
  XOR3X2 U1521 ( .A(R14[13]), .B(R14[30]), .C(R14[2]), .Y(sigma0[27]) );
  XOR3X2 U1522 ( .A(R14[12]), .B(R14[29]), .C(R14[1]), .Y(sigma0[26]) );
  XOR3X2 U1523 ( .A(R14[11]), .B(R14[28]), .C(R14[0]), .Y(sigma0[25]) );
  XOR2X1 U1524 ( .A(R1[12]), .B(R1[14]), .Y(sigma1[27]) );
  NOR2X1 U1525 ( .A(counter2[3]), .B(counter2[0]), .Y(n2073) );
  NOR2BX1 U1526 ( .AN(counter2[2]), .B(n1060), .Y(n2072) );
  NAND4X1 U1527 ( .A(n2033), .B(n2034), .C(n2035), .D(n2036), .Y(n2032) );
  AOI22X1 U1528 ( .A0(n1715), .A1(N605), .B0(n1716), .B1(N573), .Y(n2035) );
  AOI22X1 U1529 ( .A0(n605), .A1(N477), .B0(n1720), .B1(N445), .Y(n2033) );
  AOI22X1 U1530 ( .A0(n609), .A1(N541), .B0(n607), .B1(N509), .Y(n2034) );
  AOI22X1 U1531 ( .A0(n1713), .A1(N669), .B0(n1714), .B1(N637), .Y(n2036) );
  XOR3X2 U1532 ( .A(R14[14]), .B(R14[31]), .C(R14[3]), .Y(sigma0[28]) );
  XOR2X1 U1533 ( .A(R14[4]), .B(R14[15]), .Y(sigma0[29]) );
  XOR2X1 U1534 ( .A(R14[5]), .B(R14[16]), .Y(sigma0[30]) );
  XOR2X1 U1535 ( .A(R1[14]), .B(R1[16]), .Y(sigma1[29]) );
  XOR2X1 U1536 ( .A(R1[15]), .B(R1[17]), .Y(sigma1[30]) );
  NOR2X1 U1537 ( .A(n1060), .B(counter2[2]), .Y(n2076) );
  NAND4X1 U1538 ( .A(n1802), .B(n1803), .C(n1804), .D(n1805), .Y(n1801) );
  AOI22X1 U1539 ( .A0(n1715), .A1(buffer[80]), .B0(n1716), .B1(buffer[88]), 
        .Y(n1804) );
  AOI22X1 U1540 ( .A0(n1713), .A1(buffer[64]), .B0(n1714), .B1(buffer[72]), 
        .Y(n1805) );
  AOI22X1 U1541 ( .A0(n610), .A1(buffer[96]), .B0(n607), .B1(buffer[104]), .Y(
        n1803) );
  NAND4X1 U1542 ( .A(n1791), .B(n1792), .C(n1793), .D(n1794), .Y(n1790) );
  AOI22X1 U1543 ( .A0(n1715), .A1(buffer[81]), .B0(n1716), .B1(buffer[89]), 
        .Y(n1793) );
  AOI22X1 U1544 ( .A0(n1713), .A1(buffer[65]), .B0(n1714), .B1(buffer[73]), 
        .Y(n1794) );
  AOI22X1 U1545 ( .A0(n610), .A1(buffer[97]), .B0(n608), .B1(buffer[105]), .Y(
        n1792) );
  NAND4X1 U1546 ( .A(n1780), .B(n1781), .C(n1782), .D(n1783), .Y(n1779) );
  AOI22X1 U1547 ( .A0(n1715), .A1(buffer[82]), .B0(n1716), .B1(buffer[90]), 
        .Y(n1782) );
  AOI22X1 U1548 ( .A0(n1713), .A1(buffer[66]), .B0(n1714), .B1(buffer[74]), 
        .Y(n1783) );
  AOI22X1 U1549 ( .A0(n610), .A1(buffer[98]), .B0(n607), .B1(buffer[106]), .Y(
        n1781) );
  NOR2BX1 U1550 ( .AN(counter2[2]), .B(counter2[1]), .Y(n2075) );
  NOR2X1 U1551 ( .A(n1059), .B(counter2[0]), .Y(n2082) );
  NOR2X1 U1552 ( .A(n1061), .B(counter2[3]), .Y(n2074) );
  NAND4X1 U1553 ( .A(n1861), .B(n1862), .C(n1863), .D(n1864), .Y(n1855) );
  AOI22X1 U1554 ( .A0(n1727), .A1(N877), .B0(n1728), .B1(N845), .Y(n1863) );
  AOI22X1 U1555 ( .A0(n1731), .A1(N749), .B0(n602), .B1(N717), .Y(n1861) );
  AOI22X1 U1556 ( .A0(n1725), .A1(N941), .B0(n1726), .B1(N909), .Y(n1864) );
  NAND4X1 U1557 ( .A(n1850), .B(n1851), .C(n1852), .D(n1853), .Y(n1844) );
  AOI22X1 U1558 ( .A0(n1727), .A1(N878), .B0(n1728), .B1(N846), .Y(n1852) );
  AOI22X1 U1559 ( .A0(n1731), .A1(N750), .B0(n602), .B1(N718), .Y(n1850) );
  AOI22X1 U1560 ( .A0(n1725), .A1(N942), .B0(n1726), .B1(N910), .Y(n1853) );
  NAND4X1 U1561 ( .A(n1839), .B(n1840), .C(n1841), .D(n1842), .Y(n1833) );
  AOI22X1 U1562 ( .A0(n1727), .A1(N879), .B0(n1728), .B1(N847), .Y(n1841) );
  AOI22X1 U1563 ( .A0(n1731), .A1(N751), .B0(n602), .B1(N719), .Y(n1839) );
  AOI22X1 U1564 ( .A0(n1725), .A1(N943), .B0(n1726), .B1(N911), .Y(n1842) );
  NAND4X1 U1565 ( .A(n1828), .B(n1829), .C(n1830), .D(n1831), .Y(n1822) );
  AOI22X1 U1566 ( .A0(n1727), .A1(N880), .B0(n1728), .B1(N848), .Y(n1830) );
  AOI22X1 U1567 ( .A0(n1731), .A1(N752), .B0(n602), .B1(N720), .Y(n1828) );
  AOI22X1 U1568 ( .A0(n1725), .A1(N944), .B0(n1726), .B1(N912), .Y(n1831) );
  NAND4X1 U1569 ( .A(n1817), .B(n1818), .C(n1819), .D(n1820), .Y(n1811) );
  AOI22X1 U1570 ( .A0(n1727), .A1(N881), .B0(n1728), .B1(N849), .Y(n1819) );
  AOI22X1 U1571 ( .A0(n1731), .A1(N753), .B0(n602), .B1(N721), .Y(n1817) );
  AOI22X1 U1572 ( .A0(n1725), .A1(N945), .B0(n1726), .B1(N913), .Y(n1820) );
  NAND4X1 U1573 ( .A(n1773), .B(n1774), .C(n1775), .D(n1776), .Y(n1767) );
  AOI22X1 U1574 ( .A0(n1727), .A1(buffer[19]), .B0(n1728), .B1(buffer[27]), 
        .Y(n1775) );
  AOI22X1 U1575 ( .A0(n1731), .A1(buffer[51]), .B0(n602), .B1(buffer[59]), .Y(
        n1773) );
  AOI22X1 U1576 ( .A0(n1725), .A1(buffer[3]), .B0(n1726), .B1(buffer[11]), .Y(
        n1776) );
  NAND4X1 U1577 ( .A(n1762), .B(n1763), .C(n1764), .D(n1765), .Y(n1756) );
  AOI22X1 U1578 ( .A0(n1727), .A1(buffer[20]), .B0(n1728), .B1(buffer[28]), 
        .Y(n1764) );
  AOI22X1 U1579 ( .A0(n1731), .A1(buffer[52]), .B0(n601), .B1(buffer[60]), .Y(
        n1762) );
  AOI22X1 U1580 ( .A0(n1725), .A1(buffer[4]), .B0(n1726), .B1(buffer[12]), .Y(
        n1765) );
  NAND4X1 U1581 ( .A(n1751), .B(n1752), .C(n1753), .D(n1754), .Y(n1745) );
  AOI22X1 U1582 ( .A0(n1727), .A1(buffer[21]), .B0(n1728), .B1(buffer[29]), 
        .Y(n1753) );
  AOI22X1 U1583 ( .A0(n1731), .A1(buffer[53]), .B0(n602), .B1(buffer[61]), .Y(
        n1751) );
  AOI22X1 U1584 ( .A0(n1725), .A1(buffer[5]), .B0(n1726), .B1(buffer[13]), .Y(
        n1754) );
  NAND4X1 U1585 ( .A(n1742), .B(n1743), .C(n1740), .D(n1741), .Y(n774) );
  AOI22X1 U1586 ( .A0(n1727), .A1(buffer[22]), .B0(n1728), .B1(buffer[30]), 
        .Y(n1742) );
  AOI22X1 U1587 ( .A0(n1725), .A1(buffer[6]), .B0(n1726), .B1(buffer[14]), .Y(
        n1743) );
  AOI22X1 U1588 ( .A0(n1731), .A1(buffer[54]), .B0(n602), .B1(buffer[62]), .Y(
        n1740) );
  NAND4X1 U1589 ( .A(n1723), .B(n1724), .C(n1721), .D(n1722), .Y(n779) );
  AOI22X1 U1590 ( .A0(n1727), .A1(buffer[23]), .B0(n1728), .B1(buffer[31]), 
        .Y(n1723) );
  AOI22X1 U1591 ( .A0(n1725), .A1(buffer[7]), .B0(n1726), .B1(buffer[15]), .Y(
        n1724) );
  AOI22X1 U1592 ( .A0(n1731), .A1(buffer[55]), .B0(n601), .B1(buffer[63]), .Y(
        n1721) );
  NOR2X1 U1593 ( .A(n1059), .B(n1061), .Y(n2083) );
  NAND4X1 U1594 ( .A(n2068), .B(n2069), .C(n2070), .D(n2071), .Y(n2065) );
  AOI22X1 U1595 ( .A0(n1715), .A1(N602), .B0(n1716), .B1(N570), .Y(n2070) );
  AOI22X1 U1596 ( .A0(n1713), .A1(N666), .B0(n1714), .B1(N634), .Y(n2071) );
  AOI22X1 U1597 ( .A0(n605), .A1(N474), .B0(n1720), .B1(N442), .Y(n2068) );
  NAND4X1 U1598 ( .A(n2055), .B(n2056), .C(n2057), .D(n2058), .Y(n2054) );
  AOI22X1 U1599 ( .A0(n1715), .A1(N603), .B0(n1716), .B1(N571), .Y(n2057) );
  AOI22X1 U1600 ( .A0(n1713), .A1(N667), .B0(n1714), .B1(N635), .Y(n2058) );
  AOI22X1 U1601 ( .A0(n605), .A1(N475), .B0(n1720), .B1(N443), .Y(n2055) );
  NAND4X1 U1602 ( .A(n2044), .B(n2045), .C(n2046), .D(n2047), .Y(n2043) );
  AOI22X1 U1603 ( .A0(n1715), .A1(N604), .B0(n1716), .B1(N572), .Y(n2046) );
  AOI22X1 U1604 ( .A0(n1713), .A1(N668), .B0(n1714), .B1(N636), .Y(n2047) );
  AOI22X1 U1605 ( .A0(n605), .A1(N476), .B0(n1720), .B1(N444), .Y(n2044) );
  NAND4X1 U1606 ( .A(n2022), .B(n2023), .C(n2024), .D(n2025), .Y(n2021) );
  AOI22X1 U1607 ( .A0(n1715), .A1(N606), .B0(n1716), .B1(N574), .Y(n2024) );
  AOI22X1 U1608 ( .A0(n1713), .A1(N670), .B0(n1714), .B1(N638), .Y(n2025) );
  AOI22X1 U1609 ( .A0(n605), .A1(N478), .B0(n1720), .B1(N446), .Y(n2022) );
  NAND4X1 U1610 ( .A(n2011), .B(n2012), .C(n2013), .D(n2014), .Y(n2010) );
  AOI22X1 U1611 ( .A0(n1715), .A1(N607), .B0(n1716), .B1(N575), .Y(n2013) );
  AOI22X1 U1612 ( .A0(n1713), .A1(N671), .B0(n1714), .B1(N639), .Y(n2014) );
  AOI22X1 U1613 ( .A0(n605), .A1(N479), .B0(n1720), .B1(N447), .Y(n2011) );
  NAND4X1 U1614 ( .A(n2000), .B(n2001), .C(n2002), .D(n2003), .Y(n1999) );
  AOI22X1 U1615 ( .A0(n1715), .A1(N608), .B0(n1716), .B1(N576), .Y(n2002) );
  AOI22X1 U1616 ( .A0(n1713), .A1(N672), .B0(n1714), .B1(N640), .Y(n2003) );
  AOI22X1 U1617 ( .A0(n605), .A1(N480), .B0(n1720), .B1(N448), .Y(n2000) );
  NAND4X1 U1618 ( .A(n1989), .B(n1990), .C(n1991), .D(n1992), .Y(n1988) );
  AOI22X1 U1619 ( .A0(n1715), .A1(N609), .B0(n1716), .B1(N577), .Y(n1991) );
  AOI22X1 U1620 ( .A0(n1713), .A1(N673), .B0(n1714), .B1(N641), .Y(n1992) );
  AOI22X1 U1621 ( .A0(n605), .A1(N481), .B0(n1720), .B1(N449), .Y(n1989) );
  NAND4X1 U1622 ( .A(n1978), .B(n1979), .C(n1980), .D(n1981), .Y(n1977) );
  AOI22X1 U1623 ( .A0(n1715), .A1(N610), .B0(n1716), .B1(N578), .Y(n1980) );
  AOI22X1 U1624 ( .A0(n1713), .A1(N674), .B0(n1714), .B1(N642), .Y(n1981) );
  AOI22X1 U1625 ( .A0(n605), .A1(N482), .B0(n1720), .B1(N450), .Y(n1978) );
  NAND4X1 U1626 ( .A(n1967), .B(n1968), .C(n1969), .D(n1970), .Y(n1966) );
  AOI22X1 U1627 ( .A0(n1715), .A1(N611), .B0(n1716), .B1(N579), .Y(n1969) );
  AOI22X1 U1628 ( .A0(n1713), .A1(N675), .B0(n1714), .B1(N643), .Y(n1970) );
  AOI22X1 U1629 ( .A0(n605), .A1(N483), .B0(n1720), .B1(N451), .Y(n1967) );
  NAND4X1 U1630 ( .A(n1956), .B(n1957), .C(n1958), .D(n1959), .Y(n1955) );
  AOI22X1 U1631 ( .A0(n1715), .A1(N612), .B0(n1716), .B1(N580), .Y(n1958) );
  AOI22X1 U1632 ( .A0(n1713), .A1(N676), .B0(n1714), .B1(N644), .Y(n1959) );
  AOI22X1 U1633 ( .A0(n605), .A1(N484), .B0(n1720), .B1(N452), .Y(n1956) );
  NAND4X1 U1634 ( .A(n1945), .B(n1946), .C(n1947), .D(n1948), .Y(n1944) );
  AOI22X1 U1635 ( .A0(n1715), .A1(N613), .B0(n1716), .B1(N581), .Y(n1947) );
  AOI22X1 U1636 ( .A0(n1713), .A1(N677), .B0(n1714), .B1(N645), .Y(n1948) );
  AOI22X1 U1637 ( .A0(n605), .A1(N485), .B0(n1720), .B1(N453), .Y(n1945) );
  NAND4X1 U1638 ( .A(n1934), .B(n1935), .C(n1936), .D(n1937), .Y(n1933) );
  AOI22X1 U1639 ( .A0(n1715), .A1(N614), .B0(n1716), .B1(N582), .Y(n1936) );
  AOI22X1 U1640 ( .A0(n1713), .A1(N678), .B0(n1714), .B1(N646), .Y(n1937) );
  AOI22X1 U1641 ( .A0(n606), .A1(N486), .B0(n1720), .B1(N454), .Y(n1934) );
  NAND4X1 U1642 ( .A(n1923), .B(n1924), .C(n1925), .D(n1926), .Y(n1922) );
  AOI22X1 U1643 ( .A0(n1715), .A1(N615), .B0(n1716), .B1(N583), .Y(n1925) );
  AOI22X1 U1644 ( .A0(n1713), .A1(N679), .B0(n1714), .B1(N647), .Y(n1926) );
  AOI22X1 U1645 ( .A0(n606), .A1(N487), .B0(n1720), .B1(N455), .Y(n1923) );
  NAND4X1 U1646 ( .A(n1912), .B(n1913), .C(n1914), .D(n1915), .Y(n1911) );
  AOI22X1 U1647 ( .A0(n1715), .A1(N616), .B0(n1716), .B1(N584), .Y(n1914) );
  AOI22X1 U1648 ( .A0(n1713), .A1(N680), .B0(n1714), .B1(N648), .Y(n1915) );
  AOI22X1 U1649 ( .A0(n606), .A1(N488), .B0(n1720), .B1(N456), .Y(n1912) );
  NAND4X1 U1650 ( .A(n1901), .B(n1902), .C(n1903), .D(n1904), .Y(n1900) );
  AOI22X1 U1651 ( .A0(n1715), .A1(N617), .B0(n1716), .B1(N585), .Y(n1903) );
  AOI22X1 U1652 ( .A0(n1713), .A1(N681), .B0(n1714), .B1(N649), .Y(n1904) );
  AOI22X1 U1653 ( .A0(n606), .A1(N489), .B0(n1720), .B1(N457), .Y(n1901) );
  NAND4X1 U1654 ( .A(n1890), .B(n1891), .C(n1892), .D(n1893), .Y(n1889) );
  AOI22X1 U1655 ( .A0(n1715), .A1(N618), .B0(n1716), .B1(N586), .Y(n1892) );
  AOI22X1 U1656 ( .A0(n1713), .A1(N682), .B0(n1714), .B1(N650), .Y(n1893) );
  AOI22X1 U1657 ( .A0(n606), .A1(N490), .B0(n1720), .B1(N458), .Y(n1890) );
  NAND4X1 U1658 ( .A(n1879), .B(n1880), .C(n1881), .D(n1882), .Y(n1878) );
  AOI22X1 U1659 ( .A0(n1715), .A1(N619), .B0(n1716), .B1(N587), .Y(n1881) );
  AOI22X1 U1660 ( .A0(n1713), .A1(N683), .B0(n1714), .B1(N651), .Y(n1882) );
  AOI22X1 U1661 ( .A0(n606), .A1(N491), .B0(n1720), .B1(N459), .Y(n1879) );
  NAND4X1 U1662 ( .A(n1868), .B(n1869), .C(n1870), .D(n1871), .Y(n1867) );
  AOI22X1 U1663 ( .A0(n1715), .A1(N620), .B0(n1716), .B1(N588), .Y(n1870) );
  AOI22X1 U1664 ( .A0(n1713), .A1(N684), .B0(n1714), .B1(N652), .Y(n1871) );
  AOI22X1 U1665 ( .A0(n606), .A1(N492), .B0(n1720), .B1(N460), .Y(n1868) );
  AOI22X1 U1666 ( .A0(n1725), .A1(N922), .B0(n1726), .B1(N890), .Y(n2081) );
  AOI22X1 U1667 ( .A0(n1725), .A1(N923), .B0(n1726), .B1(N891), .Y(n2062) );
  AOI22X1 U1668 ( .A0(n1725), .A1(N924), .B0(n1726), .B1(N892), .Y(n2051) );
  AOI22X1 U1669 ( .A0(n1725), .A1(N925), .B0(n1726), .B1(N893), .Y(n2040) );
  AOI22X1 U1670 ( .A0(n1725), .A1(N926), .B0(n1726), .B1(N894), .Y(n2029) );
  AOI22X1 U1671 ( .A0(n1725), .A1(N927), .B0(n1726), .B1(N895), .Y(n2018) );
  AOI22X1 U1672 ( .A0(n1725), .A1(N928), .B0(n1726), .B1(N896), .Y(n2007) );
  AOI22X1 U1673 ( .A0(n1725), .A1(N929), .B0(n1726), .B1(N897), .Y(n1996) );
  AOI22X1 U1674 ( .A0(n1725), .A1(N930), .B0(n1726), .B1(N898), .Y(n1985) );
  AOI22X1 U1675 ( .A0(n1725), .A1(N931), .B0(n1726), .B1(N899), .Y(n1974) );
  AOI22X1 U1676 ( .A0(n1725), .A1(N932), .B0(n1726), .B1(N900), .Y(n1963) );
  AOI22X1 U1677 ( .A0(n1725), .A1(N933), .B0(n1726), .B1(N901), .Y(n1952) );
  AOI22X1 U1678 ( .A0(n1725), .A1(N934), .B0(n1726), .B1(N902), .Y(n1941) );
  AOI22X1 U1679 ( .A0(n1725), .A1(N935), .B0(n1726), .B1(N903), .Y(n1930) );
  AOI22X1 U1680 ( .A0(n1725), .A1(N936), .B0(n1726), .B1(N904), .Y(n1919) );
  AOI22X1 U1681 ( .A0(n1725), .A1(N937), .B0(n1726), .B1(N905), .Y(n1908) );
  AOI22X1 U1682 ( .A0(n1725), .A1(N938), .B0(n1726), .B1(N906), .Y(n1897) );
  AOI22X1 U1683 ( .A0(n1725), .A1(N939), .B0(n1726), .B1(N907), .Y(n1886) );
  AOI22X1 U1684 ( .A0(n1725), .A1(N940), .B0(n1726), .B1(N908), .Y(n1875) );
  AOI22X1 U1685 ( .A0(n1713), .A1(N685), .B0(n1714), .B1(N653), .Y(n1860) );
  AOI22X1 U1686 ( .A0(n1713), .A1(N686), .B0(n1714), .B1(N654), .Y(n1849) );
  AOI22X1 U1687 ( .A0(n1713), .A1(N687), .B0(n1714), .B1(N655), .Y(n1838) );
  AOI22X1 U1688 ( .A0(n1713), .A1(N688), .B0(n1714), .B1(N656), .Y(n1827) );
  AOI22X1 U1689 ( .A0(n1713), .A1(N689), .B0(n1714), .B1(N657), .Y(n1816) );
  AOI22X1 U1690 ( .A0(n1727), .A1(N858), .B0(n1728), .B1(N826), .Y(n2080) );
  AOI22X1 U1691 ( .A0(n1727), .A1(N859), .B0(n1728), .B1(N827), .Y(n2061) );
  AOI22X1 U1692 ( .A0(n1727), .A1(N860), .B0(n1728), .B1(N828), .Y(n2050) );
  AOI22X1 U1693 ( .A0(n1727), .A1(N861), .B0(n1728), .B1(N829), .Y(n2039) );
  AOI22X1 U1694 ( .A0(n1727), .A1(N862), .B0(n1728), .B1(N830), .Y(n2028) );
  AOI22X1 U1695 ( .A0(n1727), .A1(N863), .B0(n1728), .B1(N831), .Y(n2017) );
  AOI22X1 U1696 ( .A0(n1727), .A1(N864), .B0(n1728), .B1(N832), .Y(n2006) );
  AOI22X1 U1697 ( .A0(n1727), .A1(N865), .B0(n1728), .B1(N833), .Y(n1995) );
  AOI22X1 U1698 ( .A0(n1727), .A1(N866), .B0(n1728), .B1(N834), .Y(n1984) );
  AOI22X1 U1699 ( .A0(n1727), .A1(N867), .B0(n1728), .B1(N835), .Y(n1973) );
  AOI22X1 U1700 ( .A0(n1727), .A1(N868), .B0(n1728), .B1(N836), .Y(n1962) );
  AOI22X1 U1701 ( .A0(n1727), .A1(N869), .B0(n1728), .B1(N837), .Y(n1951) );
  AOI22X1 U1702 ( .A0(n1727), .A1(N870), .B0(n1728), .B1(N838), .Y(n1940) );
  AOI22X1 U1703 ( .A0(n1727), .A1(N871), .B0(n1728), .B1(N839), .Y(n1929) );
  AOI22X1 U1704 ( .A0(n1727), .A1(N872), .B0(n1728), .B1(N840), .Y(n1918) );
  AOI22X1 U1705 ( .A0(n1727), .A1(N873), .B0(n1728), .B1(N841), .Y(n1907) );
  AOI22X1 U1706 ( .A0(n1727), .A1(N874), .B0(n1728), .B1(N842), .Y(n1896) );
  AOI22X1 U1707 ( .A0(n1727), .A1(N875), .B0(n1728), .B1(N843), .Y(n1885) );
  AOI22X1 U1708 ( .A0(n1727), .A1(N876), .B0(n1728), .B1(N844), .Y(n1874) );
  AOI22X1 U1709 ( .A0(n1715), .A1(N621), .B0(n1716), .B1(N589), .Y(n1859) );
  AOI22X1 U1710 ( .A0(n1715), .A1(N622), .B0(n1716), .B1(N590), .Y(n1848) );
  AOI22X1 U1711 ( .A0(n1715), .A1(N623), .B0(n1716), .B1(N591), .Y(n1837) );
  AOI22X1 U1712 ( .A0(n1715), .A1(N624), .B0(n1716), .B1(N592), .Y(n1826) );
  AOI22X1 U1713 ( .A0(n1715), .A1(N625), .B0(n1716), .B1(N593), .Y(n1815) );
  AOI22X1 U1714 ( .A0(n1725), .A1(buffer[0]), .B0(n1726), .B1(buffer[8]), .Y(
        n1809) );
  AOI22X1 U1715 ( .A0(n1725), .A1(buffer[1]), .B0(n1726), .B1(buffer[9]), .Y(
        n1798) );
  AOI22X1 U1716 ( .A0(n1725), .A1(buffer[2]), .B0(n1726), .B1(buffer[10]), .Y(
        n1787) );
  AOI22X1 U1717 ( .A0(n1713), .A1(buffer[67]), .B0(n1714), .B1(buffer[75]), 
        .Y(n1772) );
  AOI22X1 U1718 ( .A0(n1713), .A1(buffer[68]), .B0(n1714), .B1(buffer[76]), 
        .Y(n1761) );
  AOI22X1 U1719 ( .A0(n1713), .A1(buffer[69]), .B0(n1714), .B1(buffer[77]), 
        .Y(n1750) );
  AOI22X1 U1720 ( .A0(n1729), .A1(buffer[38]), .B0(n604), .B1(buffer[46]), .Y(
        n1741) );
  AOI22X1 U1721 ( .A0(n610), .A1(buffer[102]), .B0(n608), .B1(buffer[110]), 
        .Y(n1737) );
  AOI22X1 U1722 ( .A0(n1729), .A1(buffer[39]), .B0(n603), .B1(buffer[47]), .Y(
        n1722) );
  AOI22X1 U1723 ( .A0(n610), .A1(buffer[103]), .B0(n607), .B1(buffer[111]), 
        .Y(n1710) );
  AOI22X1 U1724 ( .A0(n609), .A1(N538), .B0(n607), .B1(N506), .Y(n2069) );
  AOI22X1 U1725 ( .A0(n1729), .A1(N794), .B0(n603), .B1(N762), .Y(n2079) );
  AOI22X1 U1726 ( .A0(n609), .A1(N539), .B0(n607), .B1(N507), .Y(n2056) );
  AOI22X1 U1727 ( .A0(n1729), .A1(N795), .B0(n603), .B1(N763), .Y(n2060) );
  AOI22X1 U1728 ( .A0(n609), .A1(N540), .B0(n607), .B1(N508), .Y(n2045) );
  AOI22X1 U1729 ( .A0(n1729), .A1(N796), .B0(n603), .B1(N764), .Y(n2049) );
  AOI22X1 U1730 ( .A0(n1729), .A1(N797), .B0(n603), .B1(N765), .Y(n2038) );
  AOI22X1 U1731 ( .A0(n609), .A1(N542), .B0(n607), .B1(N510), .Y(n2023) );
  AOI22X1 U1732 ( .A0(n1729), .A1(N798), .B0(n603), .B1(N766), .Y(n2027) );
  AOI22X1 U1733 ( .A0(n609), .A1(N543), .B0(n607), .B1(N511), .Y(n2012) );
  AOI22X1 U1734 ( .A0(n1729), .A1(N799), .B0(n603), .B1(N767), .Y(n2016) );
  AOI22X1 U1735 ( .A0(n609), .A1(N544), .B0(n607), .B1(N512), .Y(n2001) );
  AOI22X1 U1736 ( .A0(n1729), .A1(N800), .B0(n603), .B1(N768), .Y(n2005) );
  AOI22X1 U1737 ( .A0(n609), .A1(N545), .B0(n607), .B1(N513), .Y(n1990) );
  AOI22X1 U1738 ( .A0(n1729), .A1(N801), .B0(n603), .B1(N769), .Y(n1994) );
  AOI22X1 U1739 ( .A0(n609), .A1(N546), .B0(n607), .B1(N514), .Y(n1979) );
  AOI22X1 U1740 ( .A0(n1729), .A1(N802), .B0(n603), .B1(N770), .Y(n1983) );
  AOI22X1 U1741 ( .A0(n609), .A1(N547), .B0(n607), .B1(N515), .Y(n1968) );
  AOI22X1 U1742 ( .A0(n1729), .A1(N803), .B0(n603), .B1(N771), .Y(n1972) );
  AOI22X1 U1743 ( .A0(n609), .A1(N548), .B0(n607), .B1(N516), .Y(n1957) );
  AOI22X1 U1744 ( .A0(n1729), .A1(N804), .B0(n603), .B1(N772), .Y(n1961) );
  AOI22X1 U1745 ( .A0(n609), .A1(N549), .B0(n607), .B1(N517), .Y(n1946) );
  AOI22X1 U1746 ( .A0(n1729), .A1(N805), .B0(n603), .B1(N773), .Y(n1950) );
  AOI22X1 U1747 ( .A0(n609), .A1(N550), .B0(n608), .B1(N518), .Y(n1935) );
  AOI22X1 U1748 ( .A0(n1729), .A1(N806), .B0(n604), .B1(N774), .Y(n1939) );
  AOI22X1 U1749 ( .A0(n610), .A1(N551), .B0(n608), .B1(N519), .Y(n1924) );
  AOI22X1 U1750 ( .A0(n1729), .A1(N807), .B0(n604), .B1(N775), .Y(n1928) );
  AOI22X1 U1751 ( .A0(n610), .A1(N552), .B0(n608), .B1(N520), .Y(n1913) );
  AOI22X1 U1752 ( .A0(n1729), .A1(N808), .B0(n604), .B1(N776), .Y(n1917) );
  AOI22X1 U1753 ( .A0(n609), .A1(N553), .B0(n608), .B1(N521), .Y(n1902) );
  AOI22X1 U1754 ( .A0(n1729), .A1(N809), .B0(n604), .B1(N777), .Y(n1906) );
  AOI22X1 U1755 ( .A0(n610), .A1(N554), .B0(n608), .B1(N522), .Y(n1891) );
  AOI22X1 U1756 ( .A0(n1729), .A1(N810), .B0(n604), .B1(N778), .Y(n1895) );
  AOI22X1 U1757 ( .A0(n609), .A1(N555), .B0(n608), .B1(N523), .Y(n1880) );
  AOI22X1 U1758 ( .A0(n1729), .A1(N811), .B0(n604), .B1(N779), .Y(n1884) );
  AOI22X1 U1759 ( .A0(n609), .A1(N556), .B0(n608), .B1(N524), .Y(n1869) );
  AOI22X1 U1760 ( .A0(n1729), .A1(N812), .B0(n604), .B1(N780), .Y(n1873) );
  AOI22X1 U1761 ( .A0(n1729), .A1(N813), .B0(n604), .B1(N781), .Y(n1862) );
  AOI22X1 U1762 ( .A0(n610), .A1(N557), .B0(n608), .B1(N525), .Y(n1858) );
  AOI22X1 U1763 ( .A0(n1729), .A1(N814), .B0(n604), .B1(N782), .Y(n1851) );
  AOI22X1 U1764 ( .A0(n610), .A1(N558), .B0(n608), .B1(N526), .Y(n1847) );
  AOI22X1 U1765 ( .A0(n1729), .A1(N815), .B0(n604), .B1(N783), .Y(n1840) );
  AOI22X1 U1766 ( .A0(n610), .A1(N559), .B0(n608), .B1(N527), .Y(n1836) );
  AOI22X1 U1767 ( .A0(n1729), .A1(N816), .B0(n604), .B1(N784), .Y(n1829) );
  AOI22X1 U1768 ( .A0(n610), .A1(N560), .B0(n608), .B1(N528), .Y(n1825) );
  AOI22X1 U1769 ( .A0(n1729), .A1(N817), .B0(n604), .B1(N785), .Y(n1818) );
  AOI22X1 U1770 ( .A0(n610), .A1(N561), .B0(n608), .B1(N529), .Y(n1814) );
  AOI22X1 U1771 ( .A0(n1731), .A1(N730), .B0(n601), .B1(N698), .Y(n2078) );
  AOI22X1 U1772 ( .A0(n1731), .A1(N731), .B0(n601), .B1(N699), .Y(n2059) );
  AOI22X1 U1773 ( .A0(n1731), .A1(N732), .B0(n601), .B1(N700), .Y(n2048) );
  AOI22X1 U1774 ( .A0(n1731), .A1(N733), .B0(n601), .B1(N701), .Y(n2037) );
  AOI22X1 U1775 ( .A0(n1731), .A1(N734), .B0(n601), .B1(N702), .Y(n2026) );
  AOI22X1 U1776 ( .A0(n1731), .A1(N735), .B0(n601), .B1(N703), .Y(n2015) );
  AOI22X1 U1777 ( .A0(n1731), .A1(N736), .B0(n601), .B1(N704), .Y(n2004) );
  AOI22X1 U1778 ( .A0(n1731), .A1(N737), .B0(n601), .B1(N705), .Y(n1993) );
  AOI22X1 U1779 ( .A0(n1731), .A1(N738), .B0(n601), .B1(N706), .Y(n1982) );
  AOI22X1 U1780 ( .A0(n1731), .A1(N739), .B0(n601), .B1(N707), .Y(n1971) );
  AOI22X1 U1781 ( .A0(n1731), .A1(N740), .B0(n601), .B1(N708), .Y(n1960) );
  AOI22X1 U1782 ( .A0(n1731), .A1(N741), .B0(n601), .B1(N709), .Y(n1949) );
  AOI22X1 U1783 ( .A0(n1731), .A1(N742), .B0(n602), .B1(N710), .Y(n1938) );
  AOI22X1 U1784 ( .A0(n1731), .A1(N743), .B0(n602), .B1(N711), .Y(n1927) );
  AOI22X1 U1785 ( .A0(n1731), .A1(N744), .B0(n602), .B1(N712), .Y(n1916) );
  AOI22X1 U1786 ( .A0(n1731), .A1(N745), .B0(n602), .B1(N713), .Y(n1905) );
  AOI22X1 U1787 ( .A0(n1731), .A1(N746), .B0(n602), .B1(N714), .Y(n1894) );
  AOI22X1 U1788 ( .A0(n1731), .A1(N747), .B0(n602), .B1(N715), .Y(n1883) );
  AOI22X1 U1789 ( .A0(n1731), .A1(N748), .B0(n602), .B1(N716), .Y(n1872) );
  AOI22X1 U1790 ( .A0(n606), .A1(N493), .B0(n1720), .B1(N461), .Y(n1857) );
  AOI22X1 U1791 ( .A0(n606), .A1(N494), .B0(n1720), .B1(N462), .Y(n1846) );
  AOI22X1 U1792 ( .A0(n606), .A1(N495), .B0(n1720), .B1(N463), .Y(n1835) );
  AOI22X1 U1793 ( .A0(n606), .A1(N496), .B0(n1720), .B1(N464), .Y(n1824) );
  AOI22X1 U1794 ( .A0(n606), .A1(N497), .B0(n1720), .B1(N465), .Y(n1813) );
  AOI22X1 U1795 ( .A0(n1727), .A1(buffer[16]), .B0(n1728), .B1(buffer[24]), 
        .Y(n1808) );
  AOI22X1 U1796 ( .A0(n1727), .A1(buffer[17]), .B0(n1728), .B1(buffer[25]), 
        .Y(n1797) );
  AOI22X1 U1797 ( .A0(n1727), .A1(buffer[18]), .B0(n1728), .B1(buffer[26]), 
        .Y(n1786) );
  AOI22X1 U1798 ( .A0(n1715), .A1(buffer[83]), .B0(n1716), .B1(buffer[91]), 
        .Y(n1771) );
  AOI22X1 U1799 ( .A0(n1715), .A1(buffer[84]), .B0(n1716), .B1(buffer[92]), 
        .Y(n1760) );
  AOI22X1 U1800 ( .A0(n1715), .A1(buffer[85]), .B0(n1716), .B1(buffer[93]), 
        .Y(n1749) );
  AOI22X1 U1801 ( .A0(n606), .A1(buffer[118]), .B0(n1720), .B1(buffer[126]), 
        .Y(n1736) );
  AOI22X1 U1802 ( .A0(n605), .A1(buffer[119]), .B0(n1720), .B1(buffer[127]), 
        .Y(n1709) );
  AOI22X1 U1803 ( .A0(n1729), .A1(buffer[32]), .B0(n603), .B1(buffer[40]), .Y(
        n1807) );
  AOI22X1 U1804 ( .A0(n1729), .A1(buffer[33]), .B0(n604), .B1(buffer[41]), .Y(
        n1796) );
  AOI22X1 U1805 ( .A0(n1729), .A1(buffer[34]), .B0(n603), .B1(buffer[42]), .Y(
        n1785) );
  AOI22X1 U1806 ( .A0(n1729), .A1(buffer[35]), .B0(n604), .B1(buffer[43]), .Y(
        n1774) );
  AOI22X1 U1807 ( .A0(n610), .A1(buffer[99]), .B0(n608), .B1(buffer[107]), .Y(
        n1770) );
  AOI22X1 U1808 ( .A0(n1729), .A1(buffer[36]), .B0(n604), .B1(buffer[44]), .Y(
        n1763) );
  AOI22X1 U1809 ( .A0(n610), .A1(buffer[100]), .B0(n608), .B1(buffer[108]), 
        .Y(n1759) );
  AOI22X1 U1810 ( .A0(n1729), .A1(buffer[37]), .B0(n603), .B1(buffer[45]), .Y(
        n1752) );
  AOI22X1 U1811 ( .A0(n610), .A1(buffer[101]), .B0(n607), .B1(buffer[109]), 
        .Y(n1748) );
  AOI22X1 U1812 ( .A0(n1713), .A1(buffer[70]), .B0(n1714), .B1(buffer[78]), 
        .Y(n1739) );
  AOI22X1 U1813 ( .A0(n1713), .A1(buffer[71]), .B0(n1714), .B1(buffer[79]), 
        .Y(n1712) );
  AOI22X1 U1814 ( .A0(n605), .A1(buffer[112]), .B0(n1720), .B1(buffer[120]), 
        .Y(n1802) );
  AOI22X1 U1815 ( .A0(n1731), .A1(buffer[48]), .B0(n601), .B1(buffer[56]), .Y(
        n1806) );
  AOI22X1 U1816 ( .A0(n606), .A1(buffer[113]), .B0(n1720), .B1(buffer[121]), 
        .Y(n1791) );
  AOI22X1 U1817 ( .A0(n1731), .A1(buffer[49]), .B0(n601), .B1(buffer[57]), .Y(
        n1795) );
  AOI22X1 U1818 ( .A0(n605), .A1(buffer[114]), .B0(n1720), .B1(buffer[122]), 
        .Y(n1780) );
  AOI22X1 U1819 ( .A0(n1731), .A1(buffer[50]), .B0(n602), .B1(buffer[58]), .Y(
        n1784) );
  AOI22X1 U1820 ( .A0(n606), .A1(buffer[115]), .B0(n1720), .B1(buffer[123]), 
        .Y(n1769) );
  AOI22X1 U1821 ( .A0(n606), .A1(buffer[116]), .B0(n1720), .B1(buffer[124]), 
        .Y(n1758) );
  AOI22X1 U1822 ( .A0(n605), .A1(buffer[117]), .B0(n1720), .B1(buffer[125]), 
        .Y(n1747) );
  AOI22X1 U1823 ( .A0(n1715), .A1(buffer[86]), .B0(n1716), .B1(buffer[94]), 
        .Y(n1738) );
  AOI22X1 U1824 ( .A0(n1715), .A1(buffer[87]), .B0(n1716), .B1(buffer[95]), 
        .Y(n1711) );
  OR2X2 U1825 ( .A(n418), .B(counter2[4]), .Y(n711) );
  OR2X2 U1826 ( .A(counter2[5]), .B(counter2[6]), .Y(n418) );
  XOR2X1 U1827 ( .A(R14[6]), .B(R14[17]), .Y(sigma0[31]) );
  OAI22X1 U1828 ( .A0(n719), .A1(n543), .B0(n751), .B1(n718), .Y(N2136) );
endmodule


module hash_core_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [31:2] carry;

  ADDFHX4 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX4 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX4 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX4 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX4 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX4 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX4 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  NAND2X4 U1 ( .A(n1), .B(n19), .Y(carry[4]) );
  NAND2X4 U2 ( .A(A[23]), .B(carry[23]), .Y(n23) );
  NAND2X4 U3 ( .A(B[23]), .B(carry[23]), .Y(n22) );
  NAND3X4 U4 ( .A(n12), .B(n10), .C(n11), .Y(carry[20]) );
  NAND2X4 U5 ( .A(A[14]), .B(carry[14]), .Y(n5) );
  ADDFHX2 U6 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(n2) );
  NAND3X4 U7 ( .A(n24), .B(n22), .C(n23), .Y(carry[24]) );
  NAND3X4 U8 ( .A(n6), .B(n4), .C(n5), .Y(carry[15]) );
  NAND2X2 U9 ( .A(B[14]), .B(n2), .Y(n4) );
  NAND2X4 U10 ( .A(B[19]), .B(carry[19]), .Y(n11) );
  NAND2X4 U11 ( .A(A[19]), .B(n7), .Y(n10) );
  ADDFHX4 U12 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(n7) );
  AND2X2 U13 ( .A(B[1]), .B(A[1]), .Y(n13) );
  NAND2X2 U14 ( .A(A[3]), .B(B[3]), .Y(n20) );
  NAND2X1 U15 ( .A(B[19]), .B(A[19]), .Y(n12) );
  ADDFX2 U16 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(n8) );
  NAND2X1 U17 ( .A(A[14]), .B(B[14]), .Y(n6) );
  AND2X4 U18 ( .A(n20), .B(n18), .Y(n1) );
  XOR2XL U19 ( .A(B[14]), .B(A[14]), .Y(n3) );
  XOR2X1 U20 ( .A(carry[14]), .B(n3), .Y(SUM[14]) );
  NAND2X4 U21 ( .A(B[3]), .B(carry[3]), .Y(n18) );
  XOR2X1 U22 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U23 ( .A(A[19]), .B(B[19]), .Y(n9) );
  XOR2X1 U24 ( .A(n8), .B(n9), .Y(SUM[19]) );
  NAND3BX4 U25 ( .AN(n13), .B(n15), .C(n16), .Y(carry[2]) );
  NAND2X2 U26 ( .A(A[1]), .B(n25), .Y(n15) );
  NAND2X2 U27 ( .A(B[1]), .B(n25), .Y(n16) );
  AND2X4 U28 ( .A(B[0]), .B(A[0]), .Y(n25) );
  XOR2X1 U29 ( .A(A[1]), .B(B[1]), .Y(n14) );
  XOR2X1 U30 ( .A(n25), .B(n14), .Y(SUM[1]) );
  NAND2X1 U31 ( .A(A[3]), .B(carry[3]), .Y(n19) );
  XOR2X1 U32 ( .A(B[3]), .B(A[3]), .Y(n17) );
  NAND2X1 U33 ( .A(A[23]), .B(B[23]), .Y(n24) );
  XOR2X1 U34 ( .A(carry[3]), .B(n17), .Y(SUM[3]) );
  XOR2X1 U35 ( .A(B[23]), .B(A[23]), .Y(n21) );
  XOR2X1 U36 ( .A(carry[23]), .B(n21), .Y(SUM[23]) );
endmodule


module hash_core_DW01_add_1 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [31:2] carry;

  ADDFHX4 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX4 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_1 ( .A(B[1]), .B(A[1]), .CI(n26), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX4 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX4 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX4 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX4 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  NAND3X2 U1 ( .A(n11), .B(n9), .C(n10), .Y(carry[4]) );
  NAND2X4 U2 ( .A(A[3]), .B(carry[3]), .Y(n10) );
  ADDFHX4 U3 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(n4) );
  NAND2X4 U4 ( .A(n3), .B(B[3]), .Y(n9) );
  NAND2X4 U5 ( .A(B[19]), .B(carry[19]), .Y(n14) );
  NAND3X4 U6 ( .A(n15), .B(n13), .C(n14), .Y(carry[20]) );
  NAND2X4 U7 ( .A(A[19]), .B(n6), .Y(n13) );
  ADDFHX4 U8 ( .A(A[18]), .B(B[18]), .CI(n4), .CO(n6) );
  INVX1 U9 ( .A(A[27]), .Y(n5) );
  NAND2X1 U10 ( .A(B[27]), .B(A[27]), .Y(n19) );
  NAND2X1 U11 ( .A(A[3]), .B(B[3]), .Y(n11) );
  INVX1 U12 ( .A(B[31]), .Y(n2) );
  NAND2X1 U13 ( .A(B[19]), .B(A[19]), .Y(n15) );
  AND2X4 U14 ( .A(n19), .B(n17), .Y(n1) );
  XNOR3X4 U15 ( .A(A[31]), .B(n2), .C(carry[31]), .Y(SUM[31]) );
  XOR2X1 U16 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  ADDFHX4 U17 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(n3) );
  NAND2BX4 U18 ( .AN(n5), .B(carry[27]), .Y(n17) );
  NAND2X4 U19 ( .A(n20), .B(n21), .Y(carry[24]) );
  NAND2X1 U20 ( .A(carry[23]), .B(B[23]), .Y(n20) );
  ADDFHXL U21 ( .A(A[18]), .B(B[18]), .CI(n4), .CO(n7) );
  XOR2X1 U22 ( .A(B[3]), .B(A[3]), .Y(n8) );
  XOR2X1 U23 ( .A(n3), .B(n8), .Y(SUM[3]) );
  XOR2X1 U24 ( .A(A[19]), .B(B[19]), .Y(n12) );
  XOR2X1 U25 ( .A(n7), .B(n12), .Y(SUM[19]) );
  NAND2X4 U26 ( .A(n1), .B(n18), .Y(carry[28]) );
  NAND2X1 U27 ( .A(B[27]), .B(carry[27]), .Y(n18) );
  XOR2X1 U28 ( .A(A[27]), .B(B[27]), .Y(n16) );
  XOR2X1 U29 ( .A(carry[27]), .B(n16), .Y(SUM[27]) );
  AND2X4 U30 ( .A(n24), .B(n25), .Y(n21) );
  NAND2BX4 U31 ( .AN(n22), .B(carry[23]), .Y(n24) );
  NAND2X1 U32 ( .A(B[23]), .B(A[23]), .Y(n25) );
  INVX1 U33 ( .A(A[23]), .Y(n22) );
  AND2X4 U34 ( .A(B[0]), .B(A[0]), .Y(n26) );
  XOR2X1 U35 ( .A(A[23]), .B(B[23]), .Y(n23) );
  XOR2X1 U36 ( .A(carry[23]), .B(n23), .Y(SUM[23]) );
endmodule


module hash_core_DW01_add_2 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   [31:2] carry;

  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX4 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX4 U1_1 ( .A(A[1]), .B(B[1]), .CI(n12), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX4 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX4 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX4 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX4 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX4 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  NAND2X4 U1 ( .A(B[25]), .B(carry[25]), .Y(n9) );
  NAND2X4 U2 ( .A(A[25]), .B(carry[25]), .Y(n10) );
  NAND3X4 U3 ( .A(n10), .B(n9), .C(n11), .Y(carry[26]) );
  ADDFX2 U4 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(n7) );
  NAND2X1 U5 ( .A(A[2]), .B(B[2]), .Y(n6) );
  ADDFX2 U6 ( .A(A[1]), .B(B[1]), .CI(n12), .CO(n2) );
  ADDFHX4 U7 ( .A(A[1]), .B(B[1]), .CI(n12), .CO(n1) );
  XOR2XL U8 ( .A(B[2]), .B(A[2]), .Y(n3) );
  XOR2X1 U9 ( .A(n2), .B(n3), .Y(SUM[2]) );
  NAND2X4 U10 ( .A(B[2]), .B(n1), .Y(n4) );
  NAND2X4 U11 ( .A(A[2]), .B(carry[2]), .Y(n5) );
  NAND3X4 U12 ( .A(n6), .B(n4), .C(n5), .Y(carry[3]) );
  AND2X4 U13 ( .A(B[0]), .B(A[0]), .Y(n12) );
  NAND2XL U14 ( .A(A[25]), .B(B[25]), .Y(n11) );
  XOR2XL U15 ( .A(B[25]), .B(A[25]), .Y(n8) );
  XOR2X1 U16 ( .A(n7), .B(n8), .Y(SUM[25]) );
  XOR2XL U17 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module hash_core_DW01_add_4 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [31:2] carry;

  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n24), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX4 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX4 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX4 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX4 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX4 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX4 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX4 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  NAND2BX4 U1 ( .AN(n1), .B(carry[17]), .Y(n17) );
  CLKINVX20 U2 ( .A(A[17]), .Y(n1) );
  NAND2X4 U3 ( .A(n19), .B(n17), .Y(n2) );
  NAND2X4 U4 ( .A(n3), .B(n18), .Y(carry[18]) );
  CLKINVX8 U5 ( .A(n2), .Y(n3) );
  NAND2X4 U6 ( .A(B[17]), .B(A[17]), .Y(n19) );
  NAND2X4 U7 ( .A(A[19]), .B(carry[19]), .Y(n21) );
  NAND2X4 U8 ( .A(B[19]), .B(carry[19]), .Y(n22) );
  NAND3X4 U9 ( .A(n22), .B(n21), .C(n23), .Y(carry[20]) );
  ADDFHX2 U10 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(n4) );
  NAND2X1 U11 ( .A(B[15]), .B(A[15]), .Y(n15) );
  INVX1 U12 ( .A(A[15]), .Y(n11) );
  NAND2X1 U13 ( .A(B[25]), .B(A[25]), .Y(n8) );
  NAND2X2 U14 ( .A(A[25]), .B(n4), .Y(n6) );
  XOR2XL U15 ( .A(A[25]), .B(B[25]), .Y(n5) );
  XOR2X1 U16 ( .A(carry[25]), .B(n5), .Y(SUM[25]) );
  NAND2X4 U17 ( .A(B[25]), .B(carry[25]), .Y(n7) );
  NAND3X4 U18 ( .A(n8), .B(n6), .C(n7), .Y(carry[26]) );
  NAND2X4 U19 ( .A(n15), .B(n14), .Y(n9) );
  NAND2X4 U20 ( .A(n10), .B(n13), .Y(carry[16]) );
  CLKINVX8 U21 ( .A(n9), .Y(n10) );
  NAND2BX1 U22 ( .AN(n11), .B(carry[15]), .Y(n13) );
  NAND2X4 U23 ( .A(B[15]), .B(carry[15]), .Y(n14) );
  XOR2X1 U24 ( .A(A[15]), .B(B[15]), .Y(n12) );
  XOR2X1 U25 ( .A(carry[15]), .B(n12), .Y(SUM[15]) );
  NAND2X1 U26 ( .A(B[17]), .B(carry[17]), .Y(n18) );
  XOR2X1 U27 ( .A(A[17]), .B(B[17]), .Y(n16) );
  XOR2X1 U28 ( .A(carry[17]), .B(n16), .Y(SUM[17]) );
  XOR2XL U29 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X4 U30 ( .A(B[0]), .B(A[0]), .Y(n24) );
  NAND2X1 U31 ( .A(B[19]), .B(A[19]), .Y(n23) );
  XOR2X1 U32 ( .A(A[19]), .B(B[19]), .Y(n20) );
  XOR2X1 U33 ( .A(carry[19]), .B(n20), .Y(SUM[19]) );
endmodule


module hash_core_DW01_add_5 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [31:2] carry;

  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n10), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX4 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX4 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX4 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX4 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  AND2X4 U1 ( .A(A[0]), .B(B[0]), .Y(n10) );
  NAND3X4 U2 ( .A(n7), .B(n8), .C(n9), .Y(carry[19]) );
  ADDFHX2 U3 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(n1) );
  NAND2X2 U4 ( .A(A[18]), .B(carry[18]), .Y(n7) );
  NAND2X2 U5 ( .A(B[18]), .B(carry[18]), .Y(n8) );
  XOR2XL U6 ( .A(A[23]), .B(B[23]), .Y(n2) );
  XOR2X1 U7 ( .A(carry[23]), .B(n2), .Y(SUM[23]) );
  NAND2X4 U8 ( .A(A[23]), .B(n1), .Y(n3) );
  NAND2X4 U9 ( .A(B[23]), .B(carry[23]), .Y(n4) );
  NAND2X4 U10 ( .A(B[23]), .B(A[23]), .Y(n5) );
  NAND3X4 U11 ( .A(n5), .B(n3), .C(n4), .Y(carry[24]) );
  XOR2XL U12 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X1 U13 ( .A(B[18]), .B(A[18]), .Y(n9) );
  XOR2X1 U14 ( .A(A[18]), .B(B[18]), .Y(n6) );
  XOR2X1 U15 ( .A(carry[18]), .B(n6), .Y(SUM[18]) );
endmodule


module hash_core_DW01_add_6 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;
  wire   [31:2] carry;

  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX4 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX4 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX4 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX4 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX4 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX4 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  NAND2X2 U1 ( .A(B[17]), .B(carry[17]), .Y(n18) );
  NAND2X2 U2 ( .A(A[17]), .B(carry[17]), .Y(n17) );
  NAND2X4 U3 ( .A(B[10]), .B(carry[10]), .Y(n14) );
  NAND2X4 U4 ( .A(A[10]), .B(carry[10]), .Y(n13) );
  NAND2X4 U5 ( .A(n7), .B(n5), .Y(n1) );
  NAND2X4 U6 ( .A(n2), .B(n6), .Y(carry[22]) );
  CLKINVX8 U7 ( .A(n1), .Y(n2) );
  NAND2X4 U8 ( .A(B[21]), .B(A[21]), .Y(n7) );
  NAND2X4 U9 ( .A(A[21]), .B(carry[21]), .Y(n5) );
  NAND3X4 U10 ( .A(n11), .B(n9), .C(n10), .Y(carry[5]) );
  NAND3X4 U11 ( .A(n15), .B(n13), .C(n14), .Y(carry[11]) );
  NAND3X2 U12 ( .A(n19), .B(n17), .C(n18), .Y(carry[18]) );
  XOR2X1 U13 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X4 U14 ( .A(B[0]), .B(A[0]), .Y(n3) );
  NAND2X2 U15 ( .A(B[4]), .B(carry[4]), .Y(n10) );
  NAND2X1 U16 ( .A(B[21]), .B(carry[21]), .Y(n6) );
  NAND2X1 U17 ( .A(B[17]), .B(A[17]), .Y(n19) );
  NAND2X1 U18 ( .A(B[10]), .B(A[10]), .Y(n15) );
  NAND2X1 U19 ( .A(B[4]), .B(A[4]), .Y(n11) );
  NAND2X2 U20 ( .A(A[4]), .B(carry[4]), .Y(n9) );
  XOR2X1 U21 ( .A(A[21]), .B(B[21]), .Y(n4) );
  XOR2X1 U22 ( .A(carry[21]), .B(n4), .Y(SUM[21]) );
  XOR2X1 U23 ( .A(A[4]), .B(B[4]), .Y(n8) );
  XOR2X1 U24 ( .A(carry[4]), .B(n8), .Y(SUM[4]) );
  XOR2X1 U25 ( .A(A[10]), .B(B[10]), .Y(n12) );
  XOR2X1 U26 ( .A(carry[10]), .B(n12), .Y(SUM[10]) );
  XOR2X1 U27 ( .A(A[17]), .B(B[17]), .Y(n16) );
  XOR2X1 U28 ( .A(carry[17]), .B(n16), .Y(SUM[17]) );
endmodule


module hash_core_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module hash_core_DW01_add_15 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236;

  INVX8 U2 ( .A(n105), .Y(n102) );
  OAI21X2 U3 ( .A0(n209), .A1(n188), .B0(n191), .Y(n207) );
  OAI2BB1X4 U4 ( .A0N(n210), .A1N(n211), .B0(n212), .Y(n191) );
  AOI21X2 U5 ( .A0(n82), .A1(n90), .B0(n91), .Y(n89) );
  NAND2X4 U6 ( .A(B[11]), .B(A[11]), .Y(n217) );
  OR2X4 U7 ( .A(A[28]), .B(B[28]), .Y(n82) );
  OR2X4 U8 ( .A(n172), .B(n158), .Y(n1) );
  NAND2X4 U9 ( .A(n1), .B(n160), .Y(n169) );
  CLKINVX3 U10 ( .A(n173), .Y(n172) );
  NAND2X2 U11 ( .A(n110), .B(n3), .Y(n4) );
  NAND2X2 U12 ( .A(n2), .B(n111), .Y(n5) );
  NAND2X2 U13 ( .A(n4), .B(n5), .Y(SUM[26]) );
  INVX1 U14 ( .A(n110), .Y(n2) );
  INVX2 U15 ( .A(n111), .Y(n3) );
  NAND2X4 U16 ( .A(n112), .B(n101), .Y(n110) );
  NAND2X2 U17 ( .A(B[6]), .B(A[6]), .Y(n46) );
  NOR2X4 U18 ( .A(A[13]), .B(B[13]), .Y(n28) );
  NOR2BXL U19 ( .AN(n182), .B(n186), .Y(n200) );
  INVX4 U20 ( .A(n182), .Y(n181) );
  NAND2X1 U21 ( .A(B[15]), .B(A[15]), .Y(n182) );
  XOR2X2 U22 ( .A(A[30]), .B(B[30]), .Y(n30) );
  NOR2X1 U23 ( .A(n22), .B(n195), .Y(n27) );
  NOR2X1 U24 ( .A(n195), .B(n22), .Y(n23) );
  CLKINVX3 U25 ( .A(n192), .Y(n22) );
  INVX4 U26 ( .A(n35), .Y(n209) );
  OAI21X4 U27 ( .A0(n108), .A1(n103), .B0(n109), .Y(n106) );
  INVX4 U28 ( .A(n110), .Y(n108) );
  NAND2X1 U29 ( .A(A[24]), .B(B[24]), .Y(n100) );
  INVX1 U30 ( .A(B[27]), .Y(n7) );
  INVX1 U31 ( .A(B[25]), .Y(n10) );
  AOI21X2 U32 ( .A0(n168), .A1(n169), .B0(n170), .Y(n167) );
  INVX4 U33 ( .A(n168), .Y(n150) );
  NAND2BX1 U34 ( .AN(n27), .B(n194), .Y(n35) );
  NAND2X1 U35 ( .A(n175), .B(n159), .Y(n173) );
  INVX1 U36 ( .A(n82), .Y(n79) );
  INVX1 U37 ( .A(n194), .Y(n193) );
  OAI21X1 U38 ( .A0(n225), .A1(n34), .B0(n33), .Y(n221) );
  INVX1 U39 ( .A(n31), .Y(n225) );
  OR2X2 U40 ( .A(A[7]), .B(B[7]), .Y(n43) );
  NAND2X1 U41 ( .A(B[5]), .B(A[5]), .Y(n52) );
  NAND2X2 U42 ( .A(B[20]), .B(A[20]), .Y(n128) );
  NAND2X2 U43 ( .A(n18), .B(n107), .Y(n21) );
  INVX2 U44 ( .A(n106), .Y(n18) );
  NAND2X1 U45 ( .A(n106), .B(n19), .Y(n20) );
  INVX1 U46 ( .A(n107), .Y(n19) );
  INVX1 U47 ( .A(n11), .Y(n12) );
  OAI21X1 U48 ( .A0(n201), .A1(n187), .B0(n185), .Y(n199) );
  INVX1 U49 ( .A(n202), .Y(n201) );
  NAND2X2 U50 ( .A(n120), .B(n128), .Y(n140) );
  XOR2X1 U51 ( .A(n202), .B(n203), .Y(SUM[14]) );
  NAND2X2 U52 ( .A(n17), .B(n183), .Y(n204) );
  NAND2X1 U53 ( .A(n196), .B(n207), .Y(n17) );
  OAI21X1 U54 ( .A0(n233), .A1(n234), .B0(n59), .Y(n192) );
  NAND4BBX1 U55 ( .AN(n51), .BN(n29), .C(n49), .D(n43), .Y(n195) );
  INVX1 U56 ( .A(n196), .Y(n206) );
  CLKINVX3 U57 ( .A(n28), .Y(n9) );
  NAND2X2 U58 ( .A(B[23]), .B(A[23]), .Y(n126) );
  OR2X4 U59 ( .A(A[23]), .B(B[23]), .Y(n6) );
  OAI21X4 U60 ( .A0(n70), .A1(n71), .B0(n72), .Y(n69) );
  NAND2X2 U61 ( .A(B[29]), .B(A[29]), .Y(n78) );
  CLKINVX8 U62 ( .A(n104), .Y(n103) );
  NAND2BX4 U63 ( .AN(A[27]), .B(n7), .Y(n105) );
  AND4X4 U64 ( .A(n9), .B(n196), .C(n197), .D(n198), .Y(n8) );
  NOR2BX1 U65 ( .AN(n185), .B(n187), .Y(n203) );
  INVX3 U66 ( .A(n197), .Y(n187) );
  INVX3 U67 ( .A(n198), .Y(n186) );
  NAND2XL U68 ( .A(A[19]), .B(B[19]), .Y(n157) );
  NAND2X1 U69 ( .A(n152), .B(n153), .Y(n147) );
  OAI21X1 U70 ( .A0(n50), .A1(n51), .B0(n52), .Y(n47) );
  OAI21X1 U71 ( .A0(n44), .A1(n45), .B0(n46), .Y(n39) );
  AOI21X4 U72 ( .A0(n154), .A1(n155), .B0(n156), .Y(n145) );
  CLKINVX3 U73 ( .A(n157), .Y(n156) );
  NAND2X4 U74 ( .A(B[30]), .B(A[30]), .Y(n72) );
  NOR2X4 U75 ( .A(B[30]), .B(A[30]), .Y(n74) );
  NAND2BX4 U76 ( .AN(n10), .B(A[25]), .Y(n101) );
  INVXL U77 ( .A(n117), .Y(n11) );
  XOR2X4 U78 ( .A(n166), .B(n167), .Y(SUM[19]) );
  OAI211X2 U79 ( .A0(n28), .A1(n183), .B0(n184), .C0(n185), .Y(n180) );
  NAND2X2 U80 ( .A(n226), .B(n37), .Y(n31) );
  NAND2X4 U81 ( .A(B[26]), .B(A[26]), .Y(n109) );
  NAND2X4 U82 ( .A(n8), .B(n189), .Y(n177) );
  NOR2X4 U83 ( .A(n186), .B(n187), .Y(n179) );
  XOR2X2 U84 ( .A(n25), .B(n80), .Y(SUM[28]) );
  NAND2X4 U85 ( .A(n13), .B(n66), .Y(n16) );
  AOI21X4 U86 ( .A0(n179), .A1(n180), .B0(n181), .Y(n178) );
  XNOR2X4 U87 ( .A(A[31]), .B(B[31]), .Y(n65) );
  NOR2BX1 U88 ( .AN(n98), .B(n102), .Y(n107) );
  NAND2X4 U89 ( .A(n14), .B(n65), .Y(n15) );
  NAND2X4 U90 ( .A(n15), .B(n16), .Y(SUM[31]) );
  CLKINVX3 U91 ( .A(n65), .Y(n13) );
  INVX4 U92 ( .A(n66), .Y(n14) );
  OR2X4 U93 ( .A(A[11]), .B(B[11]), .Y(n212) );
  NAND2X4 U94 ( .A(B[12]), .B(A[12]), .Y(n183) );
  NAND2X4 U95 ( .A(n20), .B(n21), .Y(SUM[27]) );
  NOR2X2 U96 ( .A(n23), .B(n193), .Y(n190) );
  OAI21X4 U97 ( .A0(n190), .A1(n188), .B0(n191), .Y(n189) );
  XOR2X4 U98 ( .A(n134), .B(n135), .Y(SUM[23]) );
  OAI21X2 U99 ( .A0(n136), .A1(n131), .B0(n130), .Y(n134) );
  OAI2BB1X1 U100 ( .A0N(n139), .A1N(n140), .B0(n129), .Y(n137) );
  XOR2X2 U101 ( .A(n88), .B(n89), .Y(SUM[29]) );
  NAND2X4 U102 ( .A(n204), .B(n9), .Y(n24) );
  NAND2X2 U103 ( .A(n24), .B(n184), .Y(n202) );
  NAND2X2 U104 ( .A(B[13]), .B(A[13]), .Y(n184) );
  NAND2X2 U105 ( .A(B[2]), .B(A[2]), .Y(n63) );
  OR2XL U106 ( .A(A[2]), .B(B[2]), .Y(n84) );
  NAND2X1 U107 ( .A(B[24]), .B(A[24]), .Y(n116) );
  NOR2X1 U108 ( .A(A[4]), .B(B[4]), .Y(n29) );
  NAND2X1 U109 ( .A(B[7]), .B(A[7]), .Y(n41) );
  NAND2X2 U110 ( .A(A[27]), .B(B[27]), .Y(n98) );
  AOI21X4 U111 ( .A0(n95), .A1(n96), .B0(n97), .Y(n94) );
  AND2X1 U112 ( .A(n116), .B(n118), .Y(n119) );
  OAI21XL U113 ( .A0(n164), .A1(n165), .B0(n87), .Y(n236) );
  NOR2BX1 U114 ( .AN(n183), .B(n206), .Y(n208) );
  NOR2BX1 U115 ( .AN(n33), .B(n34), .Y(n32) );
  NAND3X1 U116 ( .A(n213), .B(n214), .C(n215), .Y(n211) );
  INVX2 U117 ( .A(n214), .Y(n34) );
  NOR2BX1 U118 ( .AN(n184), .B(n28), .Y(n205) );
  NAND2X1 U119 ( .A(A[21]), .B(B[21]), .Y(n129) );
  NAND2X2 U120 ( .A(B[10]), .B(A[10]), .Y(n216) );
  OR2X2 U121 ( .A(A[5]), .B(B[5]), .Y(n229) );
  NOR2X4 U122 ( .A(n151), .B(n150), .Y(n154) );
  NAND2X2 U123 ( .A(n113), .B(n114), .Y(n112) );
  NAND2X4 U124 ( .A(n116), .B(n92), .Y(n114) );
  OAI2BB1X2 U125 ( .A0N(n227), .A1N(n228), .B0(n43), .Y(n194) );
  NAND2XL U126 ( .A(n81), .B(n82), .Y(n25) );
  NOR2BXL U127 ( .AN(n161), .B(n150), .Y(n171) );
  AND2X2 U128 ( .A(n216), .B(n217), .Y(n210) );
  NAND2XL U129 ( .A(n35), .B(n218), .Y(n226) );
  AND2X1 U130 ( .A(n101), .B(n113), .Y(n115) );
  AND2X1 U131 ( .A(n126), .B(n6), .Y(n135) );
  INVXL U132 ( .A(n49), .Y(n45) );
  NAND2XL U133 ( .A(n212), .B(n217), .Y(n219) );
  AND2X1 U134 ( .A(n128), .B(n143), .Y(n144) );
  XOR2X1 U135 ( .A(n35), .B(n36), .Y(SUM[8]) );
  AND2X1 U136 ( .A(n159), .B(n152), .Y(n176) );
  NOR2BXL U137 ( .AN(n87), .B(n164), .Y(n163) );
  INVXL U138 ( .A(n232), .Y(n60) );
  INVXL U139 ( .A(n165), .Y(n86) );
  NAND2X2 U140 ( .A(B[18]), .B(A[18]), .Y(n161) );
  NAND2X2 U141 ( .A(A[14]), .B(B[14]), .Y(n185) );
  NAND2XL U142 ( .A(B[1]), .B(A[1]), .Y(n87) );
  NAND2XL U143 ( .A(B[3]), .B(A[3]), .Y(n59) );
  OR2X4 U144 ( .A(A[24]), .B(B[24]), .Y(n118) );
  NAND2X1 U145 ( .A(B[17]), .B(A[17]), .Y(n160) );
  NAND2X2 U146 ( .A(B[16]), .B(A[16]), .Y(n159) );
  OR2X1 U147 ( .A(A[12]), .B(B[12]), .Y(n196) );
  NOR2BX1 U148 ( .AN(n165), .B(n26), .Y(SUM[0]) );
  NOR2XL U149 ( .A(A[0]), .B(B[0]), .Y(n26) );
  INVX1 U150 ( .A(n81), .Y(n91) );
  INVXL U151 ( .A(n132), .Y(n131) );
  INVX1 U152 ( .A(n229), .Y(n51) );
  NAND4BBX2 U153 ( .AN(n38), .BN(n34), .C(n213), .D(n212), .Y(n188) );
  NOR2BXL U154 ( .AN(n129), .B(n127), .Y(n141) );
  NOR2BX1 U155 ( .AN(n130), .B(n131), .Y(n138) );
  INVX1 U156 ( .A(n137), .Y(n136) );
  INVX1 U157 ( .A(n98), .Y(n97) );
  INVX1 U158 ( .A(n218), .Y(n38) );
  NAND3X1 U159 ( .A(n229), .B(n49), .C(n230), .Y(n228) );
  NOR2BX1 U160 ( .AN(n46), .B(n231), .Y(n227) );
  NAND2X1 U161 ( .A(n52), .B(n55), .Y(n230) );
  NAND2XL U162 ( .A(n75), .B(n78), .Y(n88) );
  XOR2X1 U163 ( .A(n169), .B(n171), .Y(SUM[18]) );
  NAND2XL U164 ( .A(n157), .B(n162), .Y(n166) );
  INVX1 U165 ( .A(n161), .Y(n170) );
  XOR2X1 U166 ( .A(n173), .B(n174), .Y(SUM[17]) );
  NOR2BXL U167 ( .AN(n160), .B(n158), .Y(n174) );
  NAND2X1 U168 ( .A(n33), .B(n37), .Y(n215) );
  INVX1 U169 ( .A(n41), .Y(n231) );
  XOR2X1 U170 ( .A(n114), .B(n115), .Y(SUM[25]) );
  XOR2X1 U171 ( .A(n140), .B(n141), .Y(SUM[21]) );
  XOR2X1 U172 ( .A(n142), .B(n144), .Y(SUM[20]) );
  XOR2X1 U173 ( .A(n137), .B(n138), .Y(SUM[22]) );
  NOR2X1 U174 ( .A(n235), .B(n236), .Y(n233) );
  NAND2X1 U175 ( .A(n84), .B(n232), .Y(n234) );
  INVX1 U176 ( .A(n63), .Y(n235) );
  AOI21X1 U177 ( .A0(n213), .A1(n221), .B0(n222), .Y(n220) );
  INVX1 U178 ( .A(n216), .Y(n222) );
  INVX1 U179 ( .A(n85), .Y(n164) );
  XOR2X1 U180 ( .A(n207), .B(n208), .Y(SUM[12]) );
  XOR2X1 U181 ( .A(n221), .B(n223), .Y(SUM[10]) );
  NOR2BX1 U182 ( .AN(n216), .B(n224), .Y(n223) );
  INVX1 U183 ( .A(n213), .Y(n224) );
  XOR2X1 U184 ( .A(n31), .B(n32), .Y(SUM[9]) );
  OAI21XL U185 ( .A0(n29), .A1(n22), .B0(n55), .Y(n53) );
  INVX1 U186 ( .A(n53), .Y(n50) );
  NOR2BX1 U187 ( .AN(n37), .B(n38), .Y(n36) );
  XOR2X1 U188 ( .A(n53), .B(n54), .Y(SUM[5]) );
  NOR2BX1 U189 ( .AN(n52), .B(n51), .Y(n54) );
  XOR2X1 U190 ( .A(n47), .B(n48), .Y(SUM[6]) );
  NOR2BX1 U191 ( .AN(n46), .B(n45), .Y(n48) );
  INVX1 U192 ( .A(n43), .Y(n42) );
  XOR2X1 U193 ( .A(n39), .B(n40), .Y(SUM[7]) );
  NOR2BX1 U194 ( .AN(n41), .B(n42), .Y(n40) );
  INVX1 U195 ( .A(n47), .Y(n44) );
  INVX1 U196 ( .A(n84), .Y(n62) );
  XOR2X1 U197 ( .A(n64), .B(n83), .Y(SUM[2]) );
  NOR2BX1 U198 ( .AN(n63), .B(n62), .Y(n83) );
  OAI2BB1X1 U199 ( .A0N(n85), .A1N(n86), .B0(n87), .Y(n64) );
  XOR2X1 U200 ( .A(n192), .B(n56), .Y(SUM[4]) );
  NOR2BX1 U201 ( .AN(n55), .B(n29), .Y(n56) );
  XOR2X1 U202 ( .A(n57), .B(n58), .Y(SUM[3]) );
  OAI21XL U203 ( .A0(n61), .A1(n62), .B0(n63), .Y(n57) );
  NOR2BX1 U204 ( .AN(n59), .B(n60), .Y(n58) );
  INVX1 U205 ( .A(n64), .Y(n61) );
  XOR2X1 U206 ( .A(n86), .B(n163), .Y(SUM[1]) );
  NAND2X2 U207 ( .A(B[28]), .B(A[28]), .Y(n81) );
  NAND2X1 U208 ( .A(B[9]), .B(A[9]), .Y(n33) );
  NAND2X1 U209 ( .A(B[8]), .B(A[8]), .Y(n37) );
  XNOR2X4 U210 ( .A(n30), .B(n76), .Y(SUM[30]) );
  OR2X2 U211 ( .A(A[6]), .B(B[6]), .Y(n49) );
  OR2X2 U212 ( .A(A[16]), .B(B[16]), .Y(n152) );
  OR2X2 U213 ( .A(A[20]), .B(B[20]), .Y(n143) );
  OR2X2 U214 ( .A(A[8]), .B(B[8]), .Y(n218) );
  OR2X2 U215 ( .A(A[9]), .B(B[9]), .Y(n214) );
  NAND2X1 U216 ( .A(B[4]), .B(A[4]), .Y(n55) );
  OR2X2 U217 ( .A(A[3]), .B(B[3]), .Y(n232) );
  OR2X2 U218 ( .A(A[1]), .B(B[1]), .Y(n85) );
  XOR2X1 U219 ( .A(n219), .B(n220), .Y(SUM[11]) );
  XOR2X1 U220 ( .A(n204), .B(n205), .Y(SUM[13]) );
  NAND2X1 U221 ( .A(B[0]), .B(A[0]), .Y(n165) );
  NAND2X4 U222 ( .A(n177), .B(n178), .Y(n148) );
  OR2XL U223 ( .A(A[25]), .B(B[25]), .Y(n113) );
  NAND2XL U224 ( .A(A[29]), .B(B[29]), .Y(n71) );
  NAND2XL U225 ( .A(n148), .B(n152), .Y(n175) );
  XOR2X1 U226 ( .A(n148), .B(n176), .Y(SUM[16]) );
  XOR2X1 U227 ( .A(n199), .B(n200), .Y(SUM[15]) );
  INVX4 U228 ( .A(n162), .Y(n151) );
  NAND3BX2 U229 ( .AN(n99), .B(n104), .C(n105), .Y(n93) );
  AND2X4 U230 ( .A(n133), .B(n132), .Y(n123) );
  NAND3BX2 U231 ( .AN(n127), .B(n132), .C(n6), .Y(n121) );
  NOR2BXL U232 ( .AN(n109), .B(n103), .Y(n111) );
  XOR2X1 U233 ( .A(n12), .B(n119), .Y(SUM[24]) );
  INVX8 U234 ( .A(n90), .Y(n80) );
  AOI21X4 U235 ( .A0(n67), .A1(n68), .B0(n69), .Y(n66) );
  NOR2X4 U236 ( .A(A[30]), .B(B[30]), .Y(n70) );
  NOR2X4 U237 ( .A(n73), .B(n74), .Y(n67) );
  CLKINVX3 U238 ( .A(n75), .Y(n73) );
  AOI21X4 U239 ( .A0(n75), .A1(n68), .B0(n77), .Y(n76) );
  CLKINVX3 U240 ( .A(n78), .Y(n77) );
  OAI21X4 U241 ( .A0(n80), .A1(n79), .B0(n81), .Y(n68) );
  OR2X4 U242 ( .A(A[29]), .B(B[29]), .Y(n75) );
  OAI21X4 U243 ( .A0(n92), .A1(n93), .B0(n94), .Y(n90) );
  OAI211X2 U244 ( .A0(n99), .A1(n100), .B0(n101), .C0(n109), .Y(n96) );
  NOR2X4 U245 ( .A(A[25]), .B(B[25]), .Y(n99) );
  NOR2X4 U246 ( .A(n102), .B(n103), .Y(n95) );
  OR2X4 U247 ( .A(A[26]), .B(B[26]), .Y(n104) );
  NAND2X4 U248 ( .A(n117), .B(n118), .Y(n92) );
  OAI21X4 U249 ( .A0(n120), .A1(n121), .B0(n122), .Y(n117) );
  AOI21X4 U250 ( .A0(n123), .A1(n124), .B0(n125), .Y(n122) );
  CLKINVX3 U251 ( .A(n126), .Y(n125) );
  OAI211X2 U252 ( .A0(n127), .A1(n128), .B0(n129), .C0(n130), .Y(n124) );
  OR2X4 U253 ( .A(A[23]), .B(B[23]), .Y(n133) );
  OR2X4 U254 ( .A(A[22]), .B(B[22]), .Y(n132) );
  NAND2X4 U255 ( .A(B[22]), .B(A[22]), .Y(n130) );
  CLKINVX3 U256 ( .A(n139), .Y(n127) );
  OR2X4 U257 ( .A(A[21]), .B(B[21]), .Y(n139) );
  NAND2X4 U258 ( .A(n142), .B(n143), .Y(n120) );
  NAND2X4 U259 ( .A(n146), .B(n145), .Y(n142) );
  NAND3BX4 U260 ( .AN(n147), .B(n148), .C(n149), .Y(n146) );
  NOR2X4 U261 ( .A(n150), .B(n151), .Y(n149) );
  OAI211X2 U262 ( .A0(n158), .A1(n159), .B0(n160), .C0(n161), .Y(n155) );
  OR2X4 U263 ( .A(A[19]), .B(B[19]), .Y(n162) );
  OR2X4 U264 ( .A(A[18]), .B(B[18]), .Y(n168) );
  CLKINVX3 U265 ( .A(n153), .Y(n158) );
  OR2X4 U266 ( .A(A[17]), .B(B[17]), .Y(n153) );
  OR2X4 U267 ( .A(A[15]), .B(B[15]), .Y(n198) );
  OR2X4 U268 ( .A(A[14]), .B(B[14]), .Y(n197) );
  OR2X4 U269 ( .A(A[10]), .B(B[10]), .Y(n213) );
endmodule


module hash_core_DW01_add_16 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224;

  OAI21X2 U2 ( .A0(n196), .A1(n171), .B0(n176), .Y(n194) );
  CLKINVX8 U3 ( .A(n87), .Y(n85) );
  NAND2X1 U4 ( .A(n15), .B(n19), .Y(n202) );
  NAND2X2 U5 ( .A(B[8]), .B(A[8]), .Y(n19) );
  INVX4 U6 ( .A(n183), .Y(n169) );
  NAND3BX4 U7 ( .AN(n86), .B(n87), .C(n88), .Y(n74) );
  NAND2X1 U8 ( .A(B[9]), .B(A[9]), .Y(n15) );
  OAI21X1 U9 ( .A0(n32), .A1(n33), .B0(n34), .Y(n29) );
  NOR2X4 U10 ( .A(n113), .B(n114), .Y(n105) );
  INVX8 U11 ( .A(n116), .Y(n113) );
  INVX8 U12 ( .A(n115), .Y(n114) );
  NOR2X4 U13 ( .A(n169), .B(n170), .Y(n162) );
  OAI21X4 U14 ( .A0(n189), .A1(n9), .B0(n167), .Y(n187) );
  INVX4 U15 ( .A(n190), .Y(n189) );
  OAI21X1 U16 ( .A0(n186), .A1(n170), .B0(n168), .Y(n184) );
  AOI21X1 U17 ( .A0(n172), .A1(n177), .B0(n178), .Y(n175) );
  INVX2 U18 ( .A(n61), .Y(n71) );
  OR2X2 U19 ( .A(A[14]), .B(B[14]), .Y(n182) );
  OR2X2 U20 ( .A(A[9]), .B(B[9]), .Y(n201) );
  OR2X2 U21 ( .A(A[7]), .B(B[7]), .Y(n25) );
  NAND2X1 U22 ( .A(B[7]), .B(A[7]), .Y(n23) );
  OR2X2 U23 ( .A(A[21]), .B(B[21]), .Y(n122) );
  NAND2X1 U24 ( .A(B[14]), .B(A[14]), .Y(n168) );
  INVX1 U25 ( .A(n182), .Y(n170) );
  NAND2X1 U26 ( .A(B[12]), .B(A[12]), .Y(n166) );
  CLKINVX3 U27 ( .A(n201), .Y(n16) );
  INVX4 U28 ( .A(n122), .Y(n109) );
  NAND2X1 U29 ( .A(B[21]), .B(A[21]), .Y(n111) );
  NAND2X1 U30 ( .A(n64), .B(n220), .Y(n222) );
  OR2X2 U31 ( .A(A[3]), .B(B[3]), .Y(n220) );
  NAND2X1 U32 ( .A(B[2]), .B(A[2]), .Y(n45) );
  INVX4 U33 ( .A(n95), .Y(n86) );
  NAND2X1 U34 ( .A(n158), .B(n142), .Y(n156) );
  NAND2X2 U35 ( .A(B[20]), .B(A[20]), .Y(n110) );
  INVX1 U36 ( .A(n140), .Y(n139) );
  NAND2X4 U37 ( .A(B[26]), .B(A[26]), .Y(n83) );
  NAND2BX4 U38 ( .AN(n47), .B(n48), .Y(n6) );
  OAI21X2 U39 ( .A0(n175), .A1(n171), .B0(n176), .Y(n174) );
  AOI21X1 U40 ( .A0(n151), .A1(n152), .B0(n153), .Y(n150) );
  OAI2BB1X2 U41 ( .A0N(n122), .A1N(n123), .B0(n111), .Y(n120) );
  INVX2 U42 ( .A(n108), .Y(n107) );
  NAND2X2 U43 ( .A(B[11]), .B(A[11]), .Y(n204) );
  OR2X1 U44 ( .A(A[2]), .B(B[2]), .Y(n64) );
  CLKINVX3 U45 ( .A(n180), .Y(n172) );
  AOI21X4 U46 ( .A0(n162), .A1(n163), .B0(n164), .Y(n161) );
  NAND2X2 U47 ( .A(B[29]), .B(A[29]), .Y(n58) );
  NOR2BX1 U48 ( .AN(n15), .B(n16), .Y(n14) );
  NAND4BBX4 U49 ( .AN(n20), .BN(n16), .C(n200), .D(n199), .Y(n171) );
  INVX3 U50 ( .A(n136), .Y(n141) );
  NAND2X2 U51 ( .A(B[18]), .B(A[18]), .Y(n144) );
  AOI21X2 U52 ( .A0(n137), .A1(n138), .B0(n139), .Y(n128) );
  NOR2X4 U53 ( .A(n134), .B(n133), .Y(n137) );
  CLKBUFX2 U54 ( .A(n82), .Y(n1) );
  OAI211X2 U55 ( .A0(n9), .A1(n166), .B0(n167), .C0(n168), .Y(n163) );
  NAND2X2 U56 ( .A(n55), .B(n58), .Y(n68) );
  INVX2 U57 ( .A(n58), .Y(n57) );
  NOR2X4 U58 ( .A(n133), .B(n134), .Y(n132) );
  INVX8 U59 ( .A(n145), .Y(n134) );
  NAND2X1 U60 ( .A(B[19]), .B(A[19]), .Y(n140) );
  XOR2X1 U61 ( .A(n123), .B(n124), .Y(SUM[21]) );
  INVX2 U62 ( .A(n29), .Y(n26) );
  INVXL U63 ( .A(n99), .Y(n2) );
  INVX1 U64 ( .A(n2), .Y(n3) );
  INVX2 U65 ( .A(n179), .Y(n178) );
  CLKINVX8 U66 ( .A(n88), .Y(n84) );
  NAND2BX4 U67 ( .AN(n173), .B(n174), .Y(n160) );
  NAND2X1 U68 ( .A(n102), .B(n110), .Y(n123) );
  OAI21X4 U69 ( .A0(n52), .A1(n58), .B0(n53), .Y(n51) );
  NOR2X4 U70 ( .A(A[30]), .B(B[30]), .Y(n52) );
  AOI21X2 U71 ( .A0(n55), .A1(n50), .B0(n57), .Y(n56) );
  NAND2X4 U72 ( .A(n94), .B(n1), .Y(n92) );
  NAND2X4 U73 ( .A(n95), .B(n96), .Y(n94) );
  NAND2X4 U74 ( .A(B[28]), .B(A[28]), .Y(n61) );
  NAND2X4 U75 ( .A(B[25]), .B(A[25]), .Y(n82) );
  NAND2X4 U76 ( .A(n47), .B(n4), .Y(n5) );
  NAND2X4 U77 ( .A(n5), .B(n6), .Y(SUM[31]) );
  INVX4 U78 ( .A(n48), .Y(n4) );
  OR2X4 U79 ( .A(n119), .B(n114), .Y(n7) );
  NAND2X4 U80 ( .A(n7), .B(n112), .Y(n117) );
  INVX2 U81 ( .A(n120), .Y(n119) );
  NAND2X4 U82 ( .A(B[22]), .B(A[22]), .Y(n112) );
  XOR2X4 U83 ( .A(n117), .B(n118), .Y(SUM[23]) );
  OR2X4 U84 ( .A(n91), .B(n85), .Y(n8) );
  NAND2X4 U85 ( .A(n8), .B(n83), .Y(n89) );
  INVX4 U86 ( .A(n92), .Y(n91) );
  XOR2X4 U87 ( .A(n89), .B(n90), .Y(SUM[27]) );
  OAI21X2 U88 ( .A0(n155), .A1(n141), .B0(n143), .Y(n152) );
  CLKINVX4 U89 ( .A(n156), .Y(n155) );
  NOR2BX1 U90 ( .AN(n1), .B(n86), .Y(n97) );
  NAND3BX4 U91 ( .AN(n130), .B(n131), .C(n132), .Y(n129) );
  NAND2X2 U92 ( .A(B[30]), .B(A[30]), .Y(n53) );
  NOR2X2 U93 ( .A(A[25]), .B(B[25]), .Y(n80) );
  NAND2X4 U94 ( .A(B[5]), .B(A[5]), .Y(n34) );
  OR2X4 U95 ( .A(A[5]), .B(B[5]), .Y(n216) );
  AOI21X1 U96 ( .A0(n62), .A1(n70), .B0(n71), .Y(n69) );
  XNOR2X4 U97 ( .A(B[31]), .B(A[31]), .Y(n47) );
  OR2X4 U98 ( .A(A[6]), .B(B[6]), .Y(n31) );
  NAND2X4 U99 ( .A(B[6]), .B(A[6]), .Y(n28) );
  NAND4BX2 U100 ( .AN(n9), .B(n181), .C(n182), .D(n183), .Y(n173) );
  NOR2X4 U101 ( .A(A[13]), .B(B[13]), .Y(n9) );
  NAND2X1 U102 ( .A(B[17]), .B(A[17]), .Y(n143) );
  NAND2X2 U103 ( .A(B[13]), .B(A[13]), .Y(n167) );
  OR2X1 U104 ( .A(A[12]), .B(B[12]), .Y(n181) );
  INVX2 U105 ( .A(n205), .Y(n20) );
  NAND2XL U106 ( .A(n213), .B(n19), .Y(n13) );
  NAND2XL U107 ( .A(B[1]), .B(A[1]), .Y(n67) );
  NOR2XL U108 ( .A(A[4]), .B(B[4]), .Y(n10) );
  NAND4BBX2 U109 ( .AN(n33), .BN(n10), .C(n31), .D(n25), .Y(n180) );
  NAND2X4 U110 ( .A(n73), .B(n98), .Y(n96) );
  OAI21XL U111 ( .A0(n147), .A1(n148), .B0(n67), .Y(n224) );
  NOR2BX1 U112 ( .AN(n166), .B(n192), .Y(n195) );
  INVX1 U113 ( .A(n65), .Y(n147) );
  NAND2XL U114 ( .A(B[24]), .B(A[24]), .Y(n98) );
  NAND2X2 U115 ( .A(B[10]), .B(A[10]), .Y(n203) );
  OR2X2 U116 ( .A(A[24]), .B(B[24]), .Y(n100) );
  INVX2 U117 ( .A(n187), .Y(n186) );
  OAI21X2 U118 ( .A0(n192), .A1(n193), .B0(n166), .Y(n190) );
  INVX2 U119 ( .A(n194), .Y(n193) );
  NAND2XL U120 ( .A(n140), .B(n145), .Y(n149) );
  INVXL U121 ( .A(n144), .Y(n153) );
  AND2X2 U122 ( .A(n203), .B(n204), .Y(n197) );
  OAI21X2 U123 ( .A0(n221), .A1(n222), .B0(n41), .Y(n177) );
  AND2X1 U124 ( .A(n142), .B(n135), .Y(n159) );
  INVXL U125 ( .A(n31), .Y(n27) );
  NOR2BXL U126 ( .AN(n108), .B(n113), .Y(n118) );
  AND2X1 U127 ( .A(n110), .B(n126), .Y(n127) );
  NOR2BXL U128 ( .AN(n67), .B(n147), .Y(n146) );
  INVXL U129 ( .A(n220), .Y(n42) );
  INVXL U130 ( .A(n148), .Y(n66) );
  NAND2XL U131 ( .A(B[3]), .B(A[3]), .Y(n41) );
  NAND2X2 U132 ( .A(A[27]), .B(B[27]), .Y(n79) );
  OR2X4 U133 ( .A(A[16]), .B(B[16]), .Y(n135) );
  NOR2XL U134 ( .A(A[0]), .B(B[0]), .Y(n12) );
  OAI21X4 U135 ( .A0(n219), .A1(n180), .B0(n179), .Y(n17) );
  OAI2BB1X4 U136 ( .A0N(n214), .A1N(n215), .B0(n25), .Y(n179) );
  INVX1 U137 ( .A(n17), .Y(n196) );
  XOR2X1 U138 ( .A(n92), .B(n93), .Y(SUM[26]) );
  INVX1 U139 ( .A(n177), .Y(n219) );
  NOR2BXL U140 ( .AN(n83), .B(n85), .Y(n93) );
  INVX1 U141 ( .A(n79), .Y(n78) );
  INVX1 U142 ( .A(n216), .Y(n33) );
  NOR2BXL U143 ( .AN(n111), .B(n109), .Y(n124) );
  OAI2BB1X2 U144 ( .A0N(n197), .A1N(n198), .B0(n199), .Y(n176) );
  NAND3X1 U145 ( .A(n200), .B(n201), .C(n202), .Y(n198) );
  NAND3X1 U146 ( .A(n216), .B(n31), .C(n217), .Y(n215) );
  NOR2BX1 U147 ( .AN(n28), .B(n218), .Y(n214) );
  NAND2X1 U148 ( .A(n34), .B(n37), .Y(n217) );
  XOR2X1 U149 ( .A(n96), .B(n97), .Y(SUM[25]) );
  XOR2X1 U150 ( .A(n184), .B(n185), .Y(SUM[15]) );
  XOR2X1 U151 ( .A(n187), .B(n188), .Y(SUM[14]) );
  NOR2BXL U152 ( .AN(n168), .B(n170), .Y(n188) );
  INVX4 U153 ( .A(n151), .Y(n133) );
  XOR2X2 U154 ( .A(n68), .B(n69), .Y(SUM[29]) );
  XOR2X1 U155 ( .A(n149), .B(n150), .Y(SUM[19]) );
  INVX1 U156 ( .A(n23), .Y(n218) );
  AND2X2 U157 ( .A(n98), .B(n100), .Y(n101) );
  XOR2XL U158 ( .A(n72), .B(n60), .Y(SUM[28]) );
  NAND2XL U159 ( .A(n61), .B(n62), .Y(n72) );
  XOR2X1 U160 ( .A(n152), .B(n154), .Y(SUM[18]) );
  NAND2XL U161 ( .A(n135), .B(n136), .Y(n130) );
  XOR2X1 U162 ( .A(n120), .B(n121), .Y(SUM[22]) );
  XOR2X1 U163 ( .A(n125), .B(n127), .Y(SUM[20]) );
  XOR2X1 U164 ( .A(n156), .B(n157), .Y(SUM[17]) );
  OAI21XL U165 ( .A0(n212), .A1(n16), .B0(n15), .Y(n208) );
  INVX1 U166 ( .A(n13), .Y(n212) );
  NOR2X1 U167 ( .A(n223), .B(n224), .Y(n221) );
  INVX1 U168 ( .A(n45), .Y(n223) );
  AOI21XL U169 ( .A0(n200), .A1(n208), .B0(n209), .Y(n207) );
  INVX1 U170 ( .A(n203), .Y(n209) );
  INVX1 U171 ( .A(n181), .Y(n192) );
  NOR2BXL U172 ( .AN(n143), .B(n141), .Y(n157) );
  NOR2BXL U173 ( .AN(n144), .B(n133), .Y(n154) );
  NAND2X1 U174 ( .A(n17), .B(n205), .Y(n213) );
  XOR2X1 U175 ( .A(n208), .B(n210), .Y(SUM[10]) );
  NOR2BX1 U176 ( .AN(n203), .B(n211), .Y(n210) );
  INVXL U177 ( .A(n200), .Y(n211) );
  XOR2X1 U178 ( .A(n194), .B(n195), .Y(SUM[12]) );
  XOR2X1 U179 ( .A(n190), .B(n191), .Y(SUM[13]) );
  NOR2BX1 U180 ( .AN(n167), .B(n9), .Y(n191) );
  XOR2X1 U181 ( .A(n13), .B(n14), .Y(SUM[9]) );
  NAND2XL U182 ( .A(n199), .B(n204), .Y(n206) );
  XOR2X1 U183 ( .A(n206), .B(n207), .Y(SUM[11]) );
  NOR2BX1 U184 ( .AN(n148), .B(n12), .Y(SUM[0]) );
  OAI21XL U185 ( .A0(n10), .A1(n219), .B0(n37), .Y(n35) );
  INVX1 U186 ( .A(n35), .Y(n32) );
  XOR2X1 U187 ( .A(n35), .B(n36), .Y(SUM[5]) );
  NOR2BX1 U188 ( .AN(n34), .B(n33), .Y(n36) );
  XOR2X1 U189 ( .A(n29), .B(n30), .Y(SUM[6]) );
  NOR2BX1 U190 ( .AN(n28), .B(n27), .Y(n30) );
  INVX1 U191 ( .A(n25), .Y(n24) );
  XOR2X1 U192 ( .A(n17), .B(n18), .Y(SUM[8]) );
  NOR2BX1 U193 ( .AN(n19), .B(n20), .Y(n18) );
  XOR2X1 U194 ( .A(n21), .B(n22), .Y(SUM[7]) );
  OAI21XL U195 ( .A0(n26), .A1(n27), .B0(n28), .Y(n21) );
  NOR2BX1 U196 ( .AN(n23), .B(n24), .Y(n22) );
  INVX1 U197 ( .A(n64), .Y(n44) );
  XOR2X1 U198 ( .A(n46), .B(n63), .Y(SUM[2]) );
  NOR2BX1 U199 ( .AN(n45), .B(n44), .Y(n63) );
  OAI2BB1X1 U200 ( .A0N(n65), .A1N(n66), .B0(n67), .Y(n46) );
  XOR2X1 U201 ( .A(n177), .B(n38), .Y(SUM[4]) );
  NOR2BX1 U202 ( .AN(n37), .B(n10), .Y(n38) );
  XOR2X1 U203 ( .A(n39), .B(n40), .Y(SUM[3]) );
  OAI21XL U204 ( .A0(n43), .A1(n44), .B0(n45), .Y(n39) );
  NOR2BX1 U205 ( .AN(n41), .B(n42), .Y(n40) );
  INVX1 U206 ( .A(n46), .Y(n43) );
  XOR2X1 U207 ( .A(n66), .B(n146), .Y(SUM[1]) );
  OR2X2 U208 ( .A(A[20]), .B(B[20]), .Y(n126) );
  OR2X2 U209 ( .A(A[8]), .B(B[8]), .Y(n205) );
  XNOR2X4 U210 ( .A(n56), .B(n11), .Y(SUM[30]) );
  XOR2X1 U211 ( .A(B[30]), .B(A[30]), .Y(n11) );
  NAND2X1 U212 ( .A(B[4]), .B(A[4]), .Y(n37) );
  OR2X2 U213 ( .A(A[1]), .B(B[1]), .Y(n65) );
  NAND2X1 U214 ( .A(B[0]), .B(A[0]), .Y(n148) );
  NAND2X4 U215 ( .A(n160), .B(n161), .Y(n131) );
  NAND2X1 U216 ( .A(B[23]), .B(A[23]), .Y(n108) );
  NOR2BX1 U217 ( .AN(n112), .B(n114), .Y(n121) );
  NAND2X1 U218 ( .A(n131), .B(n135), .Y(n158) );
  XOR2X1 U219 ( .A(n131), .B(n159), .Y(SUM[16]) );
  INVX8 U220 ( .A(n70), .Y(n60) );
  NAND2XL U221 ( .A(B[15]), .B(A[15]), .Y(n165) );
  NOR2BXL U222 ( .AN(n165), .B(n169), .Y(n185) );
  NAND3BX2 U223 ( .AN(n109), .B(n115), .C(n116), .Y(n103) );
  NOR2BXL U224 ( .AN(n79), .B(n84), .Y(n90) );
  XOR2X1 U225 ( .A(n3), .B(n101), .Y(SUM[24]) );
  AOI21X4 U226 ( .A0(n49), .A1(n50), .B0(n51), .Y(n48) );
  NOR2X4 U227 ( .A(n52), .B(n54), .Y(n49) );
  CLKINVX3 U228 ( .A(n55), .Y(n54) );
  OAI21X4 U229 ( .A0(n59), .A1(n60), .B0(n61), .Y(n50) );
  CLKINVX3 U230 ( .A(n62), .Y(n59) );
  OR2X4 U231 ( .A(A[29]), .B(B[29]), .Y(n55) );
  OAI21X4 U232 ( .A0(n73), .A1(n74), .B0(n75), .Y(n70) );
  AOI21X4 U233 ( .A0(n76), .A1(n77), .B0(n78), .Y(n75) );
  OAI211X2 U234 ( .A0(n80), .A1(n81), .B0(n82), .C0(n83), .Y(n77) );
  NAND2X4 U235 ( .A(A[24]), .B(B[24]), .Y(n81) );
  NOR2X4 U236 ( .A(n84), .B(n85), .Y(n76) );
  OR2X4 U237 ( .A(A[28]), .B(B[28]), .Y(n62) );
  OR2X4 U238 ( .A(A[27]), .B(B[27]), .Y(n88) );
  OR2X4 U239 ( .A(A[26]), .B(B[26]), .Y(n87) );
  OR2X4 U240 ( .A(A[25]), .B(B[25]), .Y(n95) );
  NAND2X4 U241 ( .A(n99), .B(n100), .Y(n73) );
  OAI21X4 U242 ( .A0(n102), .A1(n103), .B0(n104), .Y(n99) );
  AOI21X4 U243 ( .A0(n105), .A1(n106), .B0(n107), .Y(n104) );
  OAI211X2 U244 ( .A0(n109), .A1(n110), .B0(n111), .C0(n112), .Y(n106) );
  OR2X4 U245 ( .A(A[23]), .B(B[23]), .Y(n116) );
  OR2X4 U246 ( .A(A[22]), .B(B[22]), .Y(n115) );
  NAND2X4 U247 ( .A(n125), .B(n126), .Y(n102) );
  NAND2X4 U248 ( .A(n128), .B(n129), .Y(n125) );
  OAI211X2 U249 ( .A0(n141), .A1(n142), .B0(n143), .C0(n144), .Y(n138) );
  OR2X4 U250 ( .A(A[19]), .B(B[19]), .Y(n145) );
  OR2X4 U251 ( .A(A[18]), .B(B[18]), .Y(n151) );
  OR2X4 U252 ( .A(A[17]), .B(B[17]), .Y(n136) );
  NAND2X4 U253 ( .A(B[16]), .B(A[16]), .Y(n142) );
  CLKINVX3 U254 ( .A(n165), .Y(n164) );
  OR2X4 U255 ( .A(A[15]), .B(B[15]), .Y(n183) );
  OR2X4 U256 ( .A(A[11]), .B(B[11]), .Y(n199) );
  OR2X4 U257 ( .A(A[10]), .B(B[10]), .Y(n200) );
endmodule


module hash_core_DW01_add_20 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n216, n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215;

  OR2X4 U2 ( .A(n206), .B(n27), .Y(n1) );
  NAND2X4 U3 ( .A(n1), .B(n26), .Y(n202) );
  INVX1 U4 ( .A(n202), .Y(n2) );
  NAND2XL U5 ( .A(n202), .B(n3), .Y(n4) );
  NAND2X1 U6 ( .A(n2), .B(n204), .Y(n5) );
  NAND2X1 U7 ( .A(n4), .B(n5), .Y(SUM[10]) );
  INVX1 U8 ( .A(n204), .Y(n3) );
  XOR2X2 U9 ( .A(n144), .B(n145), .Y(SUM[19]) );
  XOR2X2 U10 ( .A(n31), .B(n32), .Y(SUM[7]) );
  OAI21X4 U11 ( .A0(n16), .A1(n189), .B0(n30), .Y(n24) );
  NOR2X2 U12 ( .A(A[8]), .B(B[8]), .Y(n16) );
  INVX4 U13 ( .A(n187), .Y(n186) );
  OAI21X2 U14 ( .A0(n189), .A1(n168), .B0(n190), .Y(n187) );
  NOR2X2 U15 ( .A(A[13]), .B(B[13]), .Y(n15) );
  NAND3X1 U16 ( .A(n212), .B(n71), .C(n213), .Y(n177) );
  NAND2X1 U17 ( .A(n125), .B(n126), .Y(n105) );
  NAND2X1 U18 ( .A(n101), .B(n102), .Y(n81) );
  NOR2X1 U19 ( .A(n172), .B(n173), .Y(n156) );
  INVX1 U20 ( .A(n199), .Y(n27) );
  NAND3BX2 U21 ( .AN(n178), .B(n55), .C(n177), .Y(n45) );
  INVX1 U22 ( .A(n210), .Y(n36) );
  OAI21XL U23 ( .A0(n65), .A1(n66), .B0(n67), .Y(n63) );
  BUFX3 U24 ( .A(n216), .Y(SUM[14]) );
  NAND2X1 U25 ( .A(n98), .B(n93), .Y(n96) );
  NAND2X1 U26 ( .A(n82), .B(n99), .Y(n98) );
  AOI21X2 U27 ( .A0(n174), .A1(n175), .B0(n168), .Y(n172) );
  AOI21X2 U28 ( .A0(n75), .A1(n76), .B0(n77), .Y(n66) );
  OAI21X4 U29 ( .A0(n129), .A1(n130), .B0(n131), .Y(n125) );
  NAND2X4 U30 ( .A(n152), .B(n153), .Y(n129) );
  INVX4 U31 ( .A(n28), .Y(n189) );
  OAI21X4 U32 ( .A0(n18), .A1(n186), .B0(n166), .Y(n184) );
  XOR2X2 U33 ( .A(n179), .B(n180), .Y(SUM[15]) );
  NAND2XL U34 ( .A(B[13]), .B(A[13]), .Y(n167) );
  AOI21X1 U35 ( .A0(n84), .A1(n96), .B0(n97), .Y(n95) );
  OAI21X4 U36 ( .A0(n156), .A1(n157), .B0(n158), .Y(n152) );
  NAND3BXL U37 ( .AN(n19), .B(n141), .C(n142), .Y(n130) );
  OAI21XL U38 ( .A0(n35), .A1(n36), .B0(n37), .Y(n31) );
  XOR2X1 U39 ( .A(n69), .B(n57), .Y(SUM[2]) );
  NOR2BX1 U40 ( .AN(n140), .B(n132), .Y(n131) );
  XNOR2X1 U41 ( .A(n120), .B(n13), .Y(SUM[22]) );
  INVX1 U42 ( .A(n141), .Y(n135) );
  XNOR2X1 U43 ( .A(n63), .B(n10), .Y(SUM[30]) );
  OR2X1 U44 ( .A(A[1]), .B(B[1]), .Y(n71) );
  NOR2BX1 U45 ( .AN(n46), .B(n52), .Y(n51) );
  AOI21X1 U46 ( .A0(n108), .A1(n120), .B0(n121), .Y(n119) );
  OAI21XL U47 ( .A0(n57), .A1(n58), .B0(n59), .Y(n53) );
  NOR2BXL U48 ( .AN(n55), .B(n56), .Y(n54) );
  NAND2X1 U49 ( .A(n105), .B(n116), .Y(n123) );
  NAND4BXL U50 ( .AN(n16), .B(n199), .C(n194), .D(n195), .Y(n168) );
  NAND2X1 U51 ( .A(n89), .B(n84), .Y(n9) );
  NAND3XL U52 ( .A(n43), .B(n210), .C(n211), .Y(n208) );
  NOR2BXL U53 ( .AN(n55), .B(n178), .Y(n176) );
  INVX1 U54 ( .A(n89), .Y(n97) );
  INVX1 U55 ( .A(n165), .Y(n164) );
  NAND2X1 U56 ( .A(B[2]), .B(A[2]), .Y(n59) );
  NAND2X1 U57 ( .A(B[6]), .B(A[6]), .Y(n37) );
  NAND2X1 U58 ( .A(B[1]), .B(A[1]), .Y(n72) );
  OR2X2 U59 ( .A(A[5]), .B(B[5]), .Y(n43) );
  OR2X2 U60 ( .A(A[17]), .B(B[17]), .Y(n142) );
  AND2X2 U61 ( .A(n7), .B(n8), .Y(n14) );
  NOR2X1 U62 ( .A(n47), .B(n52), .Y(n7) );
  NOR2X1 U63 ( .A(n34), .B(n36), .Y(n8) );
  OAI2BB1X2 U64 ( .A0N(n14), .A1N(n45), .B0(n175), .Y(n28) );
  NAND2XL U65 ( .A(n59), .B(n73), .Y(n69) );
  XOR2X2 U66 ( .A(n94), .B(n95), .Y(SUM[27]) );
  XNOR2X2 U67 ( .A(n96), .B(n9), .Y(SUM[26]) );
  OAI21X2 U68 ( .A0(n191), .A1(n192), .B0(n193), .Y(n173) );
  OAI21X1 U69 ( .A0(n183), .A1(n15), .B0(n167), .Y(n181) );
  NAND2X1 U70 ( .A(n61), .B(n64), .Y(n10) );
  INVXL U71 ( .A(n195), .Y(n205) );
  NOR2BXL U72 ( .AN(n165), .B(n171), .Y(n182) );
  NOR2BXL U73 ( .AN(n33), .B(n34), .Y(n32) );
  NOR2XL U74 ( .A(n46), .B(n47), .Y(n40) );
  NAND3XL U75 ( .A(n43), .B(n44), .C(n45), .Y(n42) );
  AND2X2 U76 ( .A(n37), .B(n33), .Y(n207) );
  XNOR2X1 U77 ( .A(n101), .B(n11), .Y(SUM[24]) );
  NAND2X1 U78 ( .A(n92), .B(n102), .Y(n11) );
  XNOR2X1 U79 ( .A(n75), .B(n12), .Y(SUM[28]) );
  NAND2X1 U80 ( .A(n78), .B(n76), .Y(n12) );
  NAND2X1 U81 ( .A(n113), .B(n108), .Y(n13) );
  XOR2XL U82 ( .A(n74), .B(n66), .Y(SUM[29]) );
  NOR2BXL U83 ( .AN(n140), .B(n19), .Y(n145) );
  NOR2BXL U84 ( .AN(n26), .B(n27), .Y(n25) );
  OAI21X1 U85 ( .A0(n160), .A1(n17), .B0(n161), .Y(n159) );
  OAI21X1 U86 ( .A0(n15), .A1(n166), .B0(n167), .Y(n163) );
  NAND2XL U87 ( .A(n129), .B(n138), .Y(n150) );
  NAND2XL U88 ( .A(n63), .B(n64), .Y(n62) );
  NAND2XL U89 ( .A(B[0]), .B(A[0]), .Y(n23) );
  NAND2XL U90 ( .A(B[9]), .B(A[9]), .Y(n26) );
  NAND2XL U91 ( .A(B[7]), .B(A[7]), .Y(n33) );
  NOR2XL U92 ( .A(A[12]), .B(B[12]), .Y(n18) );
  NAND2XL U93 ( .A(B[11]), .B(A[11]), .Y(n193) );
  NAND2XL U94 ( .A(B[15]), .B(A[15]), .Y(n161) );
  NAND2XL U95 ( .A(B[18]), .B(A[18]), .Y(n134) );
  NAND2XL U96 ( .A(B[19]), .B(A[19]), .Y(n140) );
  OR2XL U97 ( .A(A[16]), .B(B[16]), .Y(n153) );
  INVX1 U98 ( .A(n173), .Y(n190) );
  NAND2X1 U99 ( .A(n169), .B(n170), .Y(n157) );
  INVX1 U100 ( .A(n159), .Y(n158) );
  INVX1 U101 ( .A(n24), .Y(n206) );
  NOR2BX1 U102 ( .AN(n161), .B(n17), .Y(n180) );
  OAI2BB1X1 U103 ( .A0N(n162), .A1N(n181), .B0(n165), .Y(n179) );
  INVX1 U104 ( .A(n73), .Y(n58) );
  INVX1 U105 ( .A(n214), .Y(n56) );
  XOR2X1 U106 ( .A(n200), .B(n201), .Y(SUM[11]) );
  NAND2X1 U107 ( .A(n193), .B(n194), .Y(n200) );
  AOI21X1 U108 ( .A0(n195), .A1(n202), .B0(n203), .Y(n201) );
  INVX1 U109 ( .A(n198), .Y(n203) );
  INVX1 U110 ( .A(n184), .Y(n183) );
  NAND2X1 U111 ( .A(n194), .B(n195), .Y(n192) );
  NOR2X1 U112 ( .A(n196), .B(n197), .Y(n191) );
  NAND2X1 U113 ( .A(n26), .B(n198), .Y(n197) );
  NAND3BX1 U114 ( .AN(n40), .B(n41), .C(n42), .Y(n38) );
  INVX1 U115 ( .A(n43), .Y(n47) );
  INVX1 U116 ( .A(n44), .Y(n52) );
  INVX1 U117 ( .A(n209), .Y(n34) );
  XOR2X1 U118 ( .A(n45), .B(n51), .Y(SUM[4]) );
  NOR2BX1 U119 ( .AN(n198), .B(n205), .Y(n204) );
  XOR2X1 U120 ( .A(n187), .B(n188), .Y(SUM[12]) );
  NOR2BX1 U121 ( .AN(n166), .B(n18), .Y(n188) );
  XOR2X1 U122 ( .A(n181), .B(n182), .Y(n216) );
  XOR2X1 U123 ( .A(n38), .B(n39), .Y(SUM[6]) );
  NOR2BX1 U124 ( .AN(n37), .B(n36), .Y(n39) );
  XOR2X1 U125 ( .A(n53), .B(n54), .Y(SUM[3]) );
  XOR2X1 U126 ( .A(n48), .B(n49), .Y(SUM[5]) );
  NAND2X1 U127 ( .A(n43), .B(n41), .Y(n48) );
  AOI21X1 U128 ( .A0(n45), .A1(n44), .B0(n50), .Y(n49) );
  INVX1 U129 ( .A(n46), .Y(n50) );
  XOR2X1 U130 ( .A(n28), .B(n29), .Y(SUM[8]) );
  NOR2BX1 U131 ( .AN(n30), .B(n16), .Y(n29) );
  OAI2BB1X1 U132 ( .A0N(n176), .A1N(n177), .B0(n14), .Y(n174) );
  AOI21X1 U133 ( .A0(n162), .A1(n163), .B0(n164), .Y(n160) );
  NAND2X1 U134 ( .A(n122), .B(n117), .Y(n120) );
  NAND2X1 U135 ( .A(n106), .B(n123), .Y(n122) );
  OAI2BB1X1 U136 ( .A0N(n207), .A1N(n208), .B0(n209), .Y(n175) );
  NOR2X1 U137 ( .A(n27), .B(n30), .Y(n196) );
  NAND2X1 U138 ( .A(n149), .B(n139), .Y(n147) );
  NAND2X1 U139 ( .A(n142), .B(n150), .Y(n149) );
  INVX1 U140 ( .A(n215), .Y(n178) );
  NAND2BX1 U141 ( .AN(n59), .B(n214), .Y(n215) );
  XOR2X1 U142 ( .A(n184), .B(n185), .Y(SUM[13]) );
  NOR2BX1 U143 ( .AN(n167), .B(n15), .Y(n185) );
  XOR2X1 U144 ( .A(n147), .B(n148), .Y(SUM[18]) );
  NOR2BX1 U145 ( .AN(n134), .B(n135), .Y(n148) );
  OAI21XL U146 ( .A0(n146), .A1(n135), .B0(n134), .Y(n144) );
  INVX1 U147 ( .A(n147), .Y(n146) );
  XOR2X1 U148 ( .A(n24), .B(n25), .Y(SUM[9]) );
  INVX1 U149 ( .A(n38), .Y(n35) );
  NAND2X1 U150 ( .A(n46), .B(n41), .Y(n211) );
  NAND2X1 U151 ( .A(n72), .B(n71), .Y(n143) );
  INVX1 U152 ( .A(n78), .Y(n77) );
  NAND2X1 U153 ( .A(n87), .B(n83), .Y(n94) );
  INVX1 U154 ( .A(n68), .Y(n65) );
  XOR2X1 U155 ( .A(n125), .B(n127), .Y(SUM[20]) );
  NOR2BX1 U156 ( .AN(n116), .B(n128), .Y(n127) );
  INVX1 U157 ( .A(n126), .Y(n128) );
  INVX1 U158 ( .A(n142), .Y(n137) );
  XOR2X1 U159 ( .A(n123), .B(n124), .Y(SUM[21]) );
  NOR2BX1 U160 ( .AN(n117), .B(n115), .Y(n124) );
  INVX1 U161 ( .A(n162), .Y(n171) );
  AOI21X1 U162 ( .A0(n133), .A1(n134), .B0(n19), .Y(n132) );
  NAND2BX1 U163 ( .AN(n135), .B(n136), .Y(n133) );
  OAI21XL U164 ( .A0(n137), .A1(n138), .B0(n139), .Y(n136) );
  XOR2X1 U165 ( .A(n152), .B(n154), .Y(SUM[16]) );
  NOR2BX1 U166 ( .AN(n138), .B(n155), .Y(n154) );
  INVX1 U167 ( .A(n153), .Y(n155) );
  NAND2X1 U168 ( .A(n103), .B(n104), .Y(n101) );
  AOI21X1 U169 ( .A0(n109), .A1(n107), .B0(n110), .Y(n103) );
  NAND4BXL U170 ( .AN(n105), .B(n106), .C(n107), .D(n108), .Y(n104) );
  INVX1 U171 ( .A(n111), .Y(n110) );
  XOR2X1 U172 ( .A(n150), .B(n151), .Y(SUM[17]) );
  NOR2BX1 U173 ( .AN(n139), .B(n137), .Y(n151) );
  NAND2X1 U174 ( .A(n67), .B(n68), .Y(n74) );
  XOR2X1 U175 ( .A(n118), .B(n119), .Y(SUM[23]) );
  NAND2X1 U176 ( .A(n111), .B(n107), .Y(n118) );
  INVX1 U177 ( .A(n113), .Y(n121) );
  NAND2X1 U178 ( .A(n81), .B(n92), .Y(n99) );
  NAND2X1 U179 ( .A(n79), .B(n80), .Y(n75) );
  AOI21X1 U180 ( .A0(n85), .A1(n83), .B0(n86), .Y(n79) );
  NAND4BXL U181 ( .AN(n81), .B(n82), .C(n83), .D(n84), .Y(n80) );
  INVX1 U182 ( .A(n87), .Y(n86) );
  NOR2X1 U183 ( .A(n15), .B(n18), .Y(n169) );
  XOR2X1 U184 ( .A(n99), .B(n100), .Y(SUM[25]) );
  NOR2BX1 U185 ( .AN(n93), .B(n91), .Y(n100) );
  NOR2X1 U186 ( .A(n17), .B(n171), .Y(n170) );
  INVX1 U187 ( .A(n106), .Y(n115) );
  NAND2X1 U188 ( .A(n112), .B(n113), .Y(n109) );
  NAND2X1 U189 ( .A(n108), .B(n114), .Y(n112) );
  OAI21XL U190 ( .A0(n115), .A1(n116), .B0(n117), .Y(n114) );
  NAND2X1 U191 ( .A(n61), .B(n62), .Y(n60) );
  INVX1 U192 ( .A(n82), .Y(n91) );
  NAND2X1 U193 ( .A(n88), .B(n89), .Y(n85) );
  NAND2X1 U194 ( .A(n84), .B(n90), .Y(n88) );
  OAI21XL U195 ( .A0(n91), .A1(n92), .B0(n93), .Y(n90) );
  OAI2BB1X1 U196 ( .A0N(B[0]), .A1N(A[0]), .B0(n72), .Y(n213) );
  NOR2X1 U197 ( .A(n56), .B(n58), .Y(n212) );
  OR2X2 U198 ( .A(A[3]), .B(B[3]), .Y(n214) );
  OR2X2 U199 ( .A(A[2]), .B(B[2]), .Y(n73) );
  XOR3X2 U200 ( .A(B[31]), .B(A[31]), .C(n60), .Y(SUM[31]) );
  AND2X2 U201 ( .A(n72), .B(n70), .Y(n57) );
  NAND3X1 U202 ( .A(A[0]), .B(B[0]), .C(n71), .Y(n70) );
  OR2X2 U203 ( .A(A[10]), .B(B[10]), .Y(n195) );
  NAND2X1 U204 ( .A(B[4]), .B(A[4]), .Y(n46) );
  NAND2X1 U205 ( .A(B[5]), .B(A[5]), .Y(n41) );
  NAND2X1 U206 ( .A(B[8]), .B(A[8]), .Y(n30) );
  OR2X2 U207 ( .A(A[11]), .B(B[11]), .Y(n194) );
  NAND2X1 U208 ( .A(B[10]), .B(A[10]), .Y(n198) );
  NAND2X1 U209 ( .A(B[3]), .B(A[3]), .Y(n55) );
  OR2X2 U210 ( .A(A[4]), .B(B[4]), .Y(n44) );
  XOR2X1 U211 ( .A(n23), .B(n143), .Y(SUM[1]) );
  OR2X2 U212 ( .A(A[9]), .B(B[9]), .Y(n199) );
  OR2X2 U213 ( .A(A[6]), .B(B[6]), .Y(n210) );
  OR2X2 U214 ( .A(A[7]), .B(B[7]), .Y(n209) );
  NOR2X1 U215 ( .A(A[15]), .B(B[15]), .Y(n17) );
  NOR2X1 U216 ( .A(A[19]), .B(B[19]), .Y(n19) );
  NAND2X1 U217 ( .A(B[12]), .B(A[12]), .Y(n166) );
  NAND2X1 U218 ( .A(B[17]), .B(A[17]), .Y(n139) );
  NAND2X1 U219 ( .A(B[14]), .B(A[14]), .Y(n165) );
  NOR2X1 U220 ( .A(n21), .B(n22), .Y(SUM[0]) );
  NOR2X1 U221 ( .A(A[0]), .B(B[0]), .Y(n21) );
  AND2X2 U222 ( .A(B[0]), .B(A[0]), .Y(n22) );
  OR2X2 U223 ( .A(A[14]), .B(B[14]), .Y(n162) );
  OR2X2 U224 ( .A(A[18]), .B(B[18]), .Y(n141) );
  OR2X2 U225 ( .A(A[22]), .B(B[22]), .Y(n108) );
  NAND2X1 U226 ( .A(B[22]), .B(A[22]), .Y(n113) );
  NAND2X1 U227 ( .A(B[16]), .B(A[16]), .Y(n138) );
  NAND2X1 U228 ( .A(B[20]), .B(A[20]), .Y(n116) );
  OR2X2 U229 ( .A(A[23]), .B(B[23]), .Y(n107) );
  NAND2X1 U230 ( .A(B[21]), .B(A[21]), .Y(n117) );
  OR2X2 U231 ( .A(A[21]), .B(B[21]), .Y(n106) );
  OR2X2 U232 ( .A(A[20]), .B(B[20]), .Y(n126) );
  OR2X2 U233 ( .A(A[26]), .B(B[26]), .Y(n84) );
  NAND2X1 U234 ( .A(B[24]), .B(A[24]), .Y(n92) );
  NAND2X1 U235 ( .A(B[26]), .B(A[26]), .Y(n89) );
  OR2X2 U236 ( .A(A[27]), .B(B[27]), .Y(n83) );
  NAND2X1 U237 ( .A(B[25]), .B(A[25]), .Y(n93) );
  OR2X2 U238 ( .A(A[25]), .B(B[25]), .Y(n82) );
  NAND2X1 U239 ( .A(B[23]), .B(A[23]), .Y(n111) );
  NAND2X1 U240 ( .A(B[27]), .B(A[27]), .Y(n87) );
  OR2X2 U241 ( .A(A[28]), .B(B[28]), .Y(n76) );
  OR2X2 U242 ( .A(A[24]), .B(B[24]), .Y(n102) );
  NAND2X1 U243 ( .A(B[30]), .B(A[30]), .Y(n61) );
  NAND2X1 U244 ( .A(B[29]), .B(A[29]), .Y(n67) );
  NAND2X1 U245 ( .A(B[28]), .B(A[28]), .Y(n78) );
  OR2X2 U246 ( .A(A[30]), .B(B[30]), .Y(n64) );
  OR2X2 U247 ( .A(A[29]), .B(B[29]), .Y(n68) );
endmodule


module hash_core_DW01_add_19 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n352, n353, n354, n1, n2, n3, n4, n6, n7, n9, n11, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351;

  INVX8 U2 ( .A(n262), .Y(n274) );
  INVX1 U3 ( .A(n242), .Y(n35) );
  INVX3 U4 ( .A(n192), .Y(n197) );
  NAND2X4 U5 ( .A(B[12]), .B(A[12]), .Y(n278) );
  NAND2X2 U6 ( .A(n85), .B(n86), .Y(n84) );
  NAND2BX4 U7 ( .AN(n220), .B(n221), .Y(n218) );
  OAI21X1 U8 ( .A0(n222), .A1(n223), .B0(n224), .Y(n220) );
  INVX4 U9 ( .A(n175), .Y(n163) );
  NAND2X4 U10 ( .A(n280), .B(n2), .Y(n3) );
  NAND2X2 U11 ( .A(n1), .B(n281), .Y(n4) );
  NAND2X4 U12 ( .A(n3), .B(n4), .Y(SUM[17]) );
  CLKINVX1 U13 ( .A(n280), .Y(n1) );
  INVX4 U14 ( .A(n281), .Y(n2) );
  NAND2X2 U15 ( .A(n248), .B(n229), .Y(n280) );
  NAND2X4 U16 ( .A(B[17]), .B(A[17]), .Y(n229) );
  CLKINVX8 U17 ( .A(n307), .Y(n311) );
  BUFX20 U18 ( .A(n67), .Y(SUM[14]) );
  OAI21X4 U19 ( .A0(n106), .A1(n107), .B0(n103), .Y(n104) );
  NOR2X4 U20 ( .A(n46), .B(n111), .Y(n106) );
  OAI2BB1X2 U21 ( .A0N(B[9]), .A1N(A[9]), .B0(n83), .Y(n336) );
  NOR2X4 U22 ( .A(n162), .B(n76), .Y(n161) );
  CLKINVX3 U23 ( .A(n167), .Y(n162) );
  CLKINVX3 U24 ( .A(n314), .Y(n43) );
  BUFX3 U25 ( .A(n126), .Y(n6) );
  OAI21X4 U26 ( .A0(n81), .A1(n83), .B0(n80), .Y(n347) );
  INVX1 U27 ( .A(n285), .Y(n290) );
  NAND2X4 U28 ( .A(n19), .B(A[15]), .Y(n285) );
  NOR3X4 U29 ( .A(n88), .B(n91), .C(n92), .Y(n90) );
  NAND4BXL U30 ( .AN(n91), .B(n109), .C(n94), .D(n93), .Y(n305) );
  CLKINVX3 U31 ( .A(n108), .Y(n91) );
  INVX2 U32 ( .A(n263), .Y(n275) );
  AOI21X4 U33 ( .A0(n256), .A1(n257), .B0(n258), .Y(n253) );
  NAND2X1 U34 ( .A(n151), .B(n251), .Y(n351) );
  NAND2X2 U35 ( .A(B[1]), .B(A[1]), .Y(n151) );
  OAI21X4 U36 ( .A0(n13), .A1(n165), .B0(n166), .Y(n156) );
  NAND2X4 U37 ( .A(n113), .B(n120), .Y(n345) );
  INVX2 U38 ( .A(n310), .Y(n340) );
  NOR2X2 U39 ( .A(n81), .B(n88), .Y(n334) );
  INVX8 U40 ( .A(n308), .Y(n81) );
  BUFX8 U41 ( .A(A[27]), .Y(n7) );
  BUFX8 U42 ( .A(n352), .Y(SUM[28]) );
  NAND2X4 U43 ( .A(B[14]), .B(A[14]), .Y(n276) );
  OAI21X4 U44 ( .A0(n339), .A1(n340), .B0(n329), .Y(n337) );
  INVX4 U45 ( .A(n179), .Y(n52) );
  AOI21X4 U46 ( .A0(n180), .A1(n181), .B0(n182), .Y(n179) );
  BUFX8 U47 ( .A(n186), .Y(n9) );
  NAND2XL U48 ( .A(B[23]), .B(A[23]), .Y(n186) );
  BUFX12 U49 ( .A(n353), .Y(SUM[27]) );
  INVX4 U50 ( .A(n266), .Y(n265) );
  NAND2X2 U51 ( .A(n226), .B(n255), .Y(n266) );
  INVX2 U52 ( .A(n354), .Y(n11) );
  CLKINVX4 U53 ( .A(n11), .Y(SUM[0]) );
  CLKINVX8 U54 ( .A(n321), .Y(n295) );
  OR2X4 U55 ( .A(A[12]), .B(B[12]), .Y(n321) );
  AOI21X2 U56 ( .A0(n300), .A1(n301), .B0(n302), .Y(n297) );
  INVX2 U57 ( .A(n202), .Y(n214) );
  AND2X2 U58 ( .A(n168), .B(n9), .Y(n185) );
  AOI31XL U59 ( .A0(n187), .A1(n188), .A2(n189), .B0(n190), .Y(n183) );
  OR2X2 U60 ( .A(A[11]), .B(B[11]), .Y(n26) );
  OAI21X1 U61 ( .A0(n206), .A1(n188), .B0(n215), .Y(n209) );
  INVX2 U62 ( .A(n120), .Y(n124) );
  INVX1 U63 ( .A(n303), .Y(n302) );
  NAND2X1 U64 ( .A(B[7]), .B(A[7]), .Y(n101) );
  NAND3X1 U65 ( .A(n187), .B(n188), .C(n204), .Y(n196) );
  CLKINVX3 U66 ( .A(n306), .Y(n277) );
  NAND2X1 U67 ( .A(n39), .B(n40), .Y(n41) );
  NAND2X1 U68 ( .A(n14), .B(n90), .Y(n82) );
  NOR2X2 U69 ( .A(n87), .B(n88), .Y(n85) );
  OAI2BB1X2 U70 ( .A0N(n234), .A1N(n235), .B0(n225), .Y(n233) );
  NAND2X1 U71 ( .A(n229), .B(n247), .Y(n258) );
  NAND2X1 U72 ( .A(B[18]), .B(A[18]), .Y(n255) );
  NOR2X1 U73 ( .A(n243), .B(n244), .Y(n267) );
  NAND3BX2 U74 ( .AN(n269), .B(n24), .C(n270), .Y(n268) );
  NAND2X1 U75 ( .A(n247), .B(n285), .Y(n269) );
  AND2X2 U76 ( .A(n140), .B(n143), .Y(n60) );
  NOR2X1 U77 ( .A(n214), .B(n213), .Y(n217) );
  INVX1 U78 ( .A(n188), .Y(n219) );
  NOR3X1 U79 ( .A(n206), .B(n213), .C(n214), .Y(n212) );
  INVX1 U80 ( .A(n178), .Y(n51) );
  NAND2X2 U81 ( .A(B[5]), .B(A[5]), .Y(n113) );
  AND2X2 U82 ( .A(n123), .B(n109), .Y(n55) );
  NAND3X2 U83 ( .A(n142), .B(n143), .C(n144), .Y(n141) );
  NOR2X2 U84 ( .A(n145), .B(n146), .Y(n139) );
  NOR2BX2 U85 ( .AN(n285), .B(n274), .Y(n313) );
  NAND2X2 U86 ( .A(B[27]), .B(n7), .Y(n157) );
  OR2X2 U87 ( .A(A[25]), .B(B[25]), .Y(n175) );
  OR2X2 U88 ( .A(A[26]), .B(B[26]), .Y(n167) );
  AOI21X2 U89 ( .A0(n176), .A1(n160), .B0(n177), .Y(n172) );
  BUFX3 U90 ( .A(n105), .Y(n25) );
  NAND3X2 U91 ( .A(n306), .B(n263), .C(n307), .Y(n292) );
  NAND3BX1 U92 ( .AN(n261), .B(n262), .C(n263), .Y(n259) );
  NOR2X2 U93 ( .A(n274), .B(n275), .Y(n273) );
  INVX1 U94 ( .A(n251), .Y(n150) );
  NAND2X2 U95 ( .A(B[0]), .B(A[0]), .Y(n251) );
  AND2X2 U96 ( .A(B[26]), .B(A[26]), .Y(n13) );
  AND2X2 U97 ( .A(n89), .B(n71), .Y(n14) );
  AND2X2 U98 ( .A(n227), .B(n225), .Y(n15) );
  AND2X2 U99 ( .A(n103), .B(n101), .Y(n16) );
  AND3X2 U100 ( .A(n201), .B(n77), .C(n192), .Y(n17) );
  NAND2X1 U101 ( .A(B[25]), .B(A[25]), .Y(n169) );
  OR2X2 U102 ( .A(A[3]), .B(B[3]), .Y(n128) );
  AOI21X2 U103 ( .A0(n135), .A1(n136), .B0(n137), .Y(n134) );
  NAND2BX4 U104 ( .AN(n30), .B(n330), .Y(n299) );
  CLKINVX2 U105 ( .A(B[15]), .Y(n18) );
  CLKINVX3 U106 ( .A(n18), .Y(n19) );
  NAND3BX2 U107 ( .AN(n139), .B(n140), .C(n141), .Y(n135) );
  CLKINVX3 U108 ( .A(n305), .Y(n300) );
  NAND3XL U109 ( .A(n308), .B(n309), .C(n310), .Y(n296) );
  OAI21XL U110 ( .A0(n163), .A1(n168), .B0(n169), .Y(n165) );
  NAND2XL U111 ( .A(n36), .B(n242), .Y(n37) );
  NAND2XL U112 ( .A(n329), .B(n330), .Y(n335) );
  CLKINVX2 U113 ( .A(n299), .Y(n298) );
  NAND2X1 U114 ( .A(n226), .B(n227), .Y(n223) );
  NAND2BX2 U115 ( .AN(n205), .B(n202), .Y(n187) );
  DLY1X1 U116 ( .A(B[11]), .Y(n20) );
  XOR2X4 U117 ( .A(n89), .B(n125), .Y(SUM[4]) );
  AOI31X1 U118 ( .A0(n286), .A1(n279), .A2(n276), .B0(n288), .Y(n284) );
  NAND2X1 U119 ( .A(B[13]), .B(A[13]), .Y(n279) );
  NOR2BX2 U120 ( .AN(n83), .B(n88), .Y(n96) );
  NAND2X2 U121 ( .A(n263), .B(n262), .Y(n288) );
  OAI21X2 U122 ( .A0(n211), .A1(n200), .B0(n212), .Y(n210) );
  NAND2X2 U123 ( .A(n200), .B(n32), .Y(n33) );
  INVX2 U124 ( .A(n200), .Y(n31) );
  BUFX8 U125 ( .A(n79), .Y(n56) );
  NOR2BX2 U126 ( .AN(n80), .B(n81), .Y(n79) );
  OAI21X2 U127 ( .A0(n271), .A1(n272), .B0(n273), .Y(n270) );
  NOR4BBX4 U128 ( .AN(n299), .BN(n21), .C(n295), .D(n311), .Y(n316) );
  OR2XL U129 ( .A(A[13]), .B(B[13]), .Y(n21) );
  XNOR2X4 U130 ( .A(n231), .B(n22), .Y(SUM[21]) );
  AND2X1 U131 ( .A(n202), .B(n188), .Y(n22) );
  NAND3BX2 U132 ( .AN(n70), .B(n9), .C(n184), .Y(n195) );
  NAND4BX4 U133 ( .AN(n350), .B(n351), .C(n149), .D(n148), .Y(n115) );
  NAND4X2 U134 ( .A(n23), .B(n309), .C(n93), .D(n86), .Y(n344) );
  OAI2BB1X2 U135 ( .A0N(n245), .A1N(n235), .B0(n225), .Y(n239) );
  NOR2X2 U136 ( .A(n236), .B(n237), .Y(n245) );
  AND2X4 U137 ( .A(n156), .B(n157), .Y(n73) );
  NAND3X1 U138 ( .A(n328), .B(n331), .C(n319), .Y(n64) );
  INVX3 U139 ( .A(n319), .Y(n324) );
  NAND2XL U140 ( .A(n108), .B(n113), .Y(n121) );
  OR2XL U141 ( .A(A[9]), .B(B[9]), .Y(n23) );
  CLKINVX3 U142 ( .A(n109), .Y(n92) );
  NAND2X1 U143 ( .A(A[29]), .B(B[29]), .Y(n140) );
  NAND3BX2 U144 ( .AN(n292), .B(n294), .C(n293), .Y(n24) );
  NAND3BX1 U145 ( .AN(n114), .B(n116), .C(n115), .Y(n110) );
  NAND2X4 U146 ( .A(B[4]), .B(A[4]), .Y(n120) );
  OAI2BB1X2 U147 ( .A0N(n203), .A1N(n196), .B0(n9), .Y(n199) );
  NOR2X2 U148 ( .A(n311), .B(n295), .Y(n327) );
  INVX4 U149 ( .A(n248), .Y(n243) );
  NAND2X2 U150 ( .A(n97), .B(n98), .Y(n95) );
  NOR2X2 U151 ( .A(n99), .B(n100), .Y(n97) );
  NAND2X1 U152 ( .A(n191), .B(n192), .Y(n190) );
  OAI21X1 U153 ( .A0(n129), .A1(n130), .B0(n131), .Y(n126) );
  NOR2BX4 U154 ( .AN(n9), .B(n197), .Y(n208) );
  NAND2X2 U155 ( .A(n335), .B(n307), .Y(n331) );
  NOR2X2 U156 ( .A(n243), .B(n244), .Y(n240) );
  NAND3BX4 U157 ( .AN(n348), .B(n89), .C(n349), .Y(n98) );
  NAND2X4 U158 ( .A(B[10]), .B(A[10]), .Y(n329) );
  XNOR2X4 U159 ( .A(n135), .B(n61), .Y(SUM[30]) );
  XOR2X4 U160 ( .A(n341), .B(n342), .Y(SUM[10]) );
  NAND2BX4 U161 ( .AN(n233), .B(n221), .Y(n232) );
  OAI21X2 U162 ( .A0(n278), .A1(n277), .B0(n318), .Y(n317) );
  INVX4 U163 ( .A(n341), .Y(n339) );
  OAI21X1 U164 ( .A0(A[9]), .A1(B[9]), .B0(n309), .Y(n346) );
  NAND2X1 U165 ( .A(B[9]), .B(A[9]), .Y(n80) );
  OR2X4 U166 ( .A(A[29]), .B(B[29]), .Y(n143) );
  AND2X2 U167 ( .A(n93), .B(n94), .Y(n71) );
  NAND3X4 U168 ( .A(n82), .B(n83), .C(n84), .Y(n78) );
  NAND2X1 U169 ( .A(B[26]), .B(A[26]), .Y(n174) );
  NAND2X1 U170 ( .A(n26), .B(n310), .Y(n332) );
  NAND2X2 U171 ( .A(n264), .B(n266), .Y(n28) );
  NAND2X4 U172 ( .A(n27), .B(n265), .Y(n29) );
  NAND2X4 U173 ( .A(n28), .B(n29), .Y(SUM[18]) );
  INVX3 U174 ( .A(n264), .Y(n27) );
  NAND2X2 U175 ( .A(n328), .B(n329), .Y(n30) );
  NAND2X2 U176 ( .A(B[11]), .B(A[11]), .Y(n328) );
  NAND2X2 U177 ( .A(n299), .B(n327), .Y(n326) );
  NAND2X4 U178 ( .A(n31), .B(n238), .Y(n34) );
  NAND2X4 U179 ( .A(n33), .B(n34), .Y(SUM[20]) );
  INVX2 U180 ( .A(n238), .Y(n32) );
  OR2X4 U181 ( .A(A[21]), .B(B[21]), .Y(n202) );
  NAND2X2 U182 ( .A(B[21]), .B(A[21]), .Y(n188) );
  NAND2X4 U183 ( .A(n16), .B(n102), .Y(n86) );
  NAND2X4 U184 ( .A(n93), .B(n86), .Y(n303) );
  NAND2X2 U185 ( .A(n35), .B(n287), .Y(n38) );
  NAND2X4 U186 ( .A(n37), .B(n38), .Y(SUM[16]) );
  INVX1 U187 ( .A(n287), .Y(n36) );
  NAND2X4 U188 ( .A(n41), .B(n289), .Y(n242) );
  INVXL U189 ( .A(n261), .Y(n39) );
  INVX1 U190 ( .A(n288), .Y(n40) );
  NAND2X4 U191 ( .A(n17), .B(n200), .Y(n184) );
  AND2X2 U192 ( .A(n191), .B(n202), .Y(n77) );
  OR2X4 U193 ( .A(A[20]), .B(B[20]), .Y(n201) );
  NAND3BX2 U194 ( .AN(n183), .B(n184), .C(n185), .Y(n181) );
  NAND2X2 U195 ( .A(n74), .B(n314), .Y(n44) );
  NAND2X4 U196 ( .A(n42), .B(n43), .Y(n45) );
  NAND2X4 U197 ( .A(n44), .B(n45), .Y(n67) );
  CLKINVX3 U198 ( .A(n74), .Y(n42) );
  AND2X2 U199 ( .A(n109), .B(n110), .Y(n46) );
  NAND2X2 U200 ( .A(n60), .B(n152), .Y(n49) );
  NAND2X4 U201 ( .A(n47), .B(n48), .Y(n50) );
  NAND2X4 U202 ( .A(n49), .B(n50), .Y(SUM[29]) );
  INVX4 U203 ( .A(n60), .Y(n47) );
  INVX4 U204 ( .A(n152), .Y(n48) );
  AOI21X4 U205 ( .A0(n153), .A1(n142), .B0(n154), .Y(n152) );
  NAND2X4 U206 ( .A(n178), .B(n52), .Y(n53) );
  NAND2X2 U207 ( .A(n51), .B(n179), .Y(n54) );
  NAND2X4 U208 ( .A(n53), .B(n54), .Y(SUM[26]) );
  NAND2X2 U209 ( .A(n167), .B(n174), .Y(n178) );
  NOR2X4 U210 ( .A(n55), .B(n124), .Y(n122) );
  NAND3BX2 U211 ( .AN(n114), .B(n116), .C(n115), .Y(n123) );
  NOR2BX2 U212 ( .AN(n131), .B(n130), .Y(n147) );
  NAND2X2 U213 ( .A(B[2]), .B(A[2]), .Y(n131) );
  NOR2X2 U214 ( .A(A[3]), .B(B[3]), .Y(n350) );
  NAND2BX2 U215 ( .AN(n118), .B(n119), .Y(n117) );
  NAND3X1 U216 ( .A(n108), .B(n109), .C(n89), .Y(n119) );
  NOR2BX4 U217 ( .AN(n94), .B(n87), .Y(n349) );
  AOI21X4 U218 ( .A0(n201), .A1(n232), .B0(n211), .Y(n231) );
  NOR2BX2 U219 ( .AN(n151), .B(n250), .Y(n249) );
  INVX4 U220 ( .A(n149), .Y(n250) );
  XOR2X4 U221 ( .A(n133), .B(n134), .Y(SUM[31]) );
  NAND3X2 U222 ( .A(n260), .B(n259), .C(n285), .Y(n257) );
  AOI2BB1X4 U223 ( .A0N(n98), .A1N(n346), .B0(n347), .Y(n343) );
  INVX2 U224 ( .A(n132), .Y(n129) );
  NAND2BX2 U225 ( .AN(n120), .B(n108), .Y(n112) );
  NOR2BX4 U226 ( .AN(n120), .B(n92), .Y(n125) );
  NOR2BX4 U227 ( .AN(n329), .B(n340), .Y(n342) );
  XOR2X4 U228 ( .A(n121), .B(n122), .Y(SUM[5]) );
  XOR2X2 U229 ( .A(n132), .B(n147), .Y(SUM[2]) );
  AOI21X2 U230 ( .A0(n20), .A1(A[11]), .B0(n311), .Y(n338) );
  INVX8 U231 ( .A(n176), .Y(n164) );
  OR2X4 U232 ( .A(A[24]), .B(B[24]), .Y(n176) );
  NAND2X4 U233 ( .A(n150), .B(n57), .Y(n58) );
  NAND2X2 U234 ( .A(n251), .B(n249), .Y(n59) );
  NAND2X4 U235 ( .A(n58), .B(n59), .Y(SUM[1]) );
  INVX2 U236 ( .A(n249), .Y(n57) );
  XOR2X4 U237 ( .A(n6), .B(n127), .Y(SUM[3]) );
  OR2X4 U238 ( .A(A[10]), .B(B[10]), .Y(n310) );
  NAND2X4 U239 ( .A(B[24]), .B(A[24]), .Y(n168) );
  NAND3BX2 U240 ( .AN(n284), .B(n24), .C(n285), .Y(n282) );
  NAND2X2 U241 ( .A(n73), .B(n155), .Y(n153) );
  NAND2X2 U242 ( .A(n138), .B(n136), .Y(n61) );
  OR2X2 U243 ( .A(A[28]), .B(B[28]), .Y(n142) );
  NAND2X1 U244 ( .A(B[28]), .B(A[28]), .Y(n145) );
  XOR2X4 U245 ( .A(n64), .B(n65), .Y(SUM[12]) );
  OAI2BB1X4 U246 ( .A0N(n194), .A1N(n195), .B0(n168), .Y(n193) );
  INVX8 U247 ( .A(n75), .Y(SUM[24]) );
  NOR2X2 U248 ( .A(n76), .B(n162), .Y(n166) );
  AND2X1 U249 ( .A(n175), .B(n169), .Y(n62) );
  INVXL U250 ( .A(n101), .Y(n100) );
  XNOR2X4 U251 ( .A(n160), .B(n198), .Y(n75) );
  NAND3X4 U252 ( .A(n159), .B(n160), .C(n161), .Y(n155) );
  NOR2XL U253 ( .A(n163), .B(n164), .Y(n159) );
  AND2X1 U254 ( .A(n191), .B(n215), .Y(n69) );
  INVX2 U255 ( .A(n143), .Y(n146) );
  INVXL U256 ( .A(n138), .Y(n137) );
  XOR2X4 U257 ( .A(n117), .B(n63), .Y(SUM[6]) );
  AND2X1 U258 ( .A(n103), .B(n94), .Y(n63) );
  INVX4 U259 ( .A(n201), .Y(n213) );
  AND2X2 U260 ( .A(n145), .B(n142), .Y(n158) );
  OAI21X4 U261 ( .A0(n296), .A1(n297), .B0(n298), .Y(n293) );
  AND2X1 U262 ( .A(n278), .B(n321), .Y(n65) );
  INVXL U263 ( .A(n276), .Y(n272) );
  AND3X4 U264 ( .A(n230), .B(n229), .C(n228), .Y(n222) );
  OR2X4 U265 ( .A(A[1]), .B(B[1]), .Y(n149) );
  OR2X4 U266 ( .A(A[2]), .B(B[2]), .Y(n148) );
  OR2X4 U267 ( .A(A[4]), .B(B[4]), .Y(n109) );
  OR2X4 U268 ( .A(B[5]), .B(A[5]), .Y(n108) );
  NAND2XL U269 ( .A(B[22]), .B(A[22]), .Y(n189) );
  NAND2X2 U270 ( .A(B[20]), .B(A[20]), .Y(n205) );
  NOR2BX1 U271 ( .AN(n251), .B(n68), .Y(n354) );
  NOR2XL U272 ( .A(A[0]), .B(B[0]), .Y(n68) );
  NOR2X1 U273 ( .A(n163), .B(n164), .Y(n180) );
  NOR2XL U274 ( .A(n197), .B(n164), .Y(n194) );
  INVX1 U275 ( .A(n169), .Y(n182) );
  NOR2BX1 U276 ( .AN(n205), .B(n213), .Y(n238) );
  XNOR2X4 U277 ( .A(n216), .B(n69), .Y(SUM[22]) );
  NOR2BX2 U278 ( .AN(n247), .B(n244), .Y(n287) );
  NOR2BX1 U279 ( .AN(n116), .B(n350), .Y(n127) );
  INVX1 U280 ( .A(n145), .Y(n154) );
  NAND2X1 U281 ( .A(n112), .B(n113), .Y(n111) );
  NAND2XL U282 ( .A(n306), .B(n318), .Y(n322) );
  AND2X1 U283 ( .A(n196), .B(n191), .Y(n70) );
  INVX1 U284 ( .A(n205), .Y(n211) );
  INVX1 U285 ( .A(n148), .Y(n130) );
  NAND2X1 U286 ( .A(n169), .B(n168), .Y(n177) );
  OAI2BB1X1 U287 ( .A0N(n149), .A1N(n150), .B0(n151), .Y(n132) );
  XNOR2X4 U288 ( .A(n312), .B(n313), .Y(n72) );
  INVX8 U289 ( .A(n72), .Y(SUM[15]) );
  OAI21XL U290 ( .A0(n277), .A1(n278), .B0(n279), .Y(n271) );
  INVXL U291 ( .A(n247), .Y(n283) );
  NAND2X2 U292 ( .A(n326), .B(n278), .Y(n325) );
  AND2X1 U293 ( .A(n276), .B(n263), .Y(n74) );
  NAND2X2 U294 ( .A(B[3]), .B(A[3]), .Y(n116) );
  OAI21XL U295 ( .A0(A[13]), .A1(B[13]), .B0(n321), .Y(n320) );
  NAND2X2 U296 ( .A(n303), .B(n98), .Y(n333) );
  NOR2X4 U297 ( .A(n7), .B(B[27]), .Y(n76) );
  NAND2XL U298 ( .A(B[13]), .B(A[13]), .Y(n318) );
  NAND2X2 U299 ( .A(B[19]), .B(A[19]), .Y(n225) );
  NAND2XL U300 ( .A(B[22]), .B(A[22]), .Y(n204) );
  NAND2XL U301 ( .A(B[22]), .B(A[22]), .Y(n215) );
  NAND3X2 U302 ( .A(n228), .B(n229), .C(n246), .Y(n235) );
  NAND2XL U303 ( .A(B[18]), .B(A[18]), .Y(n246) );
  NAND2XL U304 ( .A(B[18]), .B(A[18]), .Y(n230) );
  OR2X2 U305 ( .A(A[30]), .B(B[30]), .Y(n136) );
  NAND2X1 U306 ( .A(B[30]), .B(A[30]), .Y(n138) );
  XNOR2X1 U307 ( .A(B[31]), .B(A[31]), .Y(n133) );
  NAND3BX4 U308 ( .AN(n114), .B(n116), .C(n115), .Y(n89) );
  OAI21X2 U309 ( .A0(n314), .A1(n275), .B0(n276), .Y(n312) );
  INVX4 U310 ( .A(n260), .Y(n291) );
  NOR2X2 U311 ( .A(n197), .B(n206), .Y(n203) );
  INVX3 U312 ( .A(n191), .Y(n206) );
  INVX8 U313 ( .A(n226), .Y(n237) );
  INVX8 U314 ( .A(n227), .Y(n236) );
  NOR2X2 U315 ( .A(n236), .B(n237), .Y(n234) );
  INVX4 U316 ( .A(n256), .Y(n244) );
  NAND2X1 U317 ( .A(n248), .B(n226), .Y(n254) );
  AOI21X1 U318 ( .A0(B[7]), .A1(A[7]), .B0(n87), .Y(n105) );
  INVX4 U319 ( .A(n304), .Y(n114) );
  INVX8 U320 ( .A(n309), .Y(n88) );
  INVX8 U321 ( .A(n93), .Y(n87) );
  NAND2X1 U322 ( .A(n113), .B(n112), .Y(n118) );
  NAND2XL U323 ( .A(n109), .B(n108), .Y(n348) );
  NAND2XL U324 ( .A(n108), .B(n94), .Y(n107) );
  AOI21X1 U325 ( .A0(n102), .A1(n103), .B0(n87), .Y(n99) );
  NAND3XL U326 ( .A(n116), .B(n304), .C(n115), .Y(n301) );
  NAND2X2 U327 ( .A(B[6]), .B(A[6]), .Y(n103) );
  XOR2X4 U328 ( .A(n78), .B(n56), .Y(SUM[9]) );
  XOR2X4 U329 ( .A(n95), .B(n96), .Y(SUM[8]) );
  XOR2X4 U330 ( .A(n104), .B(n25), .Y(SUM[7]) );
  XOR2X4 U331 ( .A(n144), .B(n158), .Y(n352) );
  NAND3X4 U332 ( .A(n156), .B(n157), .C(n155), .Y(n144) );
  XOR2X4 U333 ( .A(n170), .B(n171), .Y(n353) );
  NOR2BX4 U334 ( .AN(n157), .B(n76), .Y(n171) );
  OAI21X4 U335 ( .A0(n172), .A1(n173), .B0(n174), .Y(n170) );
  NAND2X4 U336 ( .A(n175), .B(n167), .Y(n173) );
  XOR2X4 U337 ( .A(n193), .B(n62), .Y(SUM[25]) );
  NOR2BX4 U338 ( .AN(n168), .B(n164), .Y(n198) );
  NAND2BX4 U339 ( .AN(n199), .B(n184), .Y(n160) );
  XOR2X4 U340 ( .A(n207), .B(n208), .Y(SUM[23]) );
  OR2X4 U341 ( .A(A[23]), .B(B[23]), .Y(n192) );
  NAND2BX4 U342 ( .AN(n209), .B(n210), .Y(n207) );
  AOI21X4 U343 ( .A0(n217), .A1(n218), .B0(n219), .Y(n216) );
  AND2X2 U344 ( .A(n205), .B(n225), .Y(n224) );
  OR2X4 U345 ( .A(A[22]), .B(B[22]), .Y(n191) );
  NAND2BX4 U346 ( .AN(n239), .B(n221), .Y(n200) );
  NAND3X4 U347 ( .A(n242), .B(n241), .C(n240), .Y(n221) );
  NOR2X4 U348 ( .A(n236), .B(n237), .Y(n241) );
  NAND2BX4 U349 ( .AN(n247), .B(n248), .Y(n228) );
  XOR2X4 U350 ( .A(n252), .B(n15), .Y(SUM[19]) );
  OR2X4 U351 ( .A(A[19]), .B(B[19]), .Y(n227) );
  OAI21X4 U352 ( .A0(n253), .A1(n254), .B0(n255), .Y(n252) );
  OR2X4 U353 ( .A(A[18]), .B(B[18]), .Y(n226) );
  OAI2BB1X4 U354 ( .A0N(n267), .A1N(n268), .B0(n229), .Y(n264) );
  AOI21X4 U355 ( .A0(n256), .A1(n282), .B0(n283), .Y(n281) );
  OR2X4 U356 ( .A(A[17]), .B(B[17]), .Y(n248) );
  OR2X4 U357 ( .A(A[16]), .B(B[16]), .Y(n256) );
  NAND2X4 U358 ( .A(B[16]), .B(A[16]), .Y(n247) );
  NOR2X4 U359 ( .A(n290), .B(n291), .Y(n289) );
  NAND3BX4 U360 ( .AN(n292), .B(n293), .C(n294), .Y(n260) );
  NOR2X4 U361 ( .A(n295), .B(n274), .Y(n294) );
  AND3X4 U362 ( .A(n279), .B(n276), .C(n286), .Y(n261) );
  NAND2BX4 U363 ( .AN(n278), .B(n306), .Y(n286) );
  OR2X4 U364 ( .A(B[15]), .B(A[15]), .Y(n262) );
  NOR3X4 U365 ( .A(n315), .B(n316), .C(n317), .Y(n314) );
  NOR2X4 U366 ( .A(n319), .B(n320), .Y(n315) );
  OR2X4 U367 ( .A(A[14]), .B(B[14]), .Y(n263) );
  XOR2X4 U368 ( .A(n322), .B(n323), .Y(SUM[13]) );
  AOI21X4 U369 ( .A0(n324), .A1(n321), .B0(n325), .Y(n323) );
  OR2X4 U370 ( .A(A[13]), .B(B[13]), .Y(n306) );
  NAND3BX4 U371 ( .AN(n332), .B(n333), .C(n334), .Y(n319) );
  NAND3X4 U372 ( .A(n310), .B(n308), .C(n336), .Y(n330) );
  XOR2X4 U373 ( .A(n337), .B(n338), .Y(SUM[11]) );
  OR2X4 U374 ( .A(A[11]), .B(B[11]), .Y(n307) );
  NAND2X4 U375 ( .A(n343), .B(n344), .Y(n341) );
  NAND3X4 U376 ( .A(n108), .B(n94), .C(n345), .Y(n102) );
  NAND2X4 U377 ( .A(B[8]), .B(A[8]), .Y(n83) );
  OR2X4 U378 ( .A(A[9]), .B(B[9]), .Y(n308) );
  OR2X4 U379 ( .A(A[8]), .B(B[8]), .Y(n309) );
  OR2X4 U380 ( .A(A[7]), .B(B[7]), .Y(n93) );
  OR2X4 U381 ( .A(A[6]), .B(B[6]), .Y(n94) );
  NAND2BX4 U382 ( .AN(n131), .B(n128), .Y(n304) );
endmodule


module hash_core_DW01_add_26 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n265, n266, n267, n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264;

  INVX1 U2 ( .A(n224), .Y(n223) );
  CLKINVX3 U3 ( .A(n103), .Y(n102) );
  INVX3 U4 ( .A(n181), .Y(n15) );
  NOR2X4 U5 ( .A(n181), .B(n192), .Y(n191) );
  INVX2 U6 ( .A(n49), .Y(n238) );
  CLKINVX3 U7 ( .A(n161), .Y(n11) );
  NAND2X4 U8 ( .A(n104), .B(n103), .Y(n1) );
  NAND2X4 U9 ( .A(n2), .B(n86), .Y(n112) );
  CLKINVX3 U10 ( .A(n1), .Y(n2) );
  AOI21X2 U11 ( .A0(n112), .A1(n101), .B0(n113), .Y(n111) );
  NAND2X1 U12 ( .A(n59), .B(n4), .Y(n5) );
  NAND2X2 U13 ( .A(n3), .B(n60), .Y(n6) );
  NAND2X4 U14 ( .A(n5), .B(n6), .Y(SUM[6]) );
  INVX1 U15 ( .A(n59), .Y(n3) );
  INVX1 U16 ( .A(n60), .Y(n4) );
  INVX1 U17 ( .A(n33), .Y(n59) );
  NOR2BX2 U18 ( .AN(n58), .B(n57), .Y(n60) );
  OR2X4 U19 ( .A(A[17]), .B(B[17]), .Y(n189) );
  NAND4BBX2 U20 ( .AN(n37), .BN(n38), .C(n61), .D(n259), .Y(n225) );
  NOR2X2 U21 ( .A(A[4]), .B(B[4]), .Y(n38) );
  NAND2X2 U22 ( .A(n62), .B(n66), .Y(n258) );
  BUFX8 U23 ( .A(n267), .Y(SUM[13]) );
  AOI21X4 U24 ( .A0(n143), .A1(n119), .B0(n144), .Y(n142) );
  OAI21X4 U25 ( .A0(n145), .A1(n146), .B0(n147), .Y(n143) );
  NOR2BX2 U26 ( .AN(n147), .B(n145), .Y(n153) );
  CLKINVX8 U27 ( .A(n120), .Y(n145) );
  NOR2X2 U28 ( .A(n148), .B(n149), .Y(n146) );
  BUFX4 U29 ( .A(n266), .Y(SUM[20]) );
  NOR2X4 U30 ( .A(B[27]), .B(A[27]), .Y(n118) );
  NOR2X4 U31 ( .A(n117), .B(n118), .Y(n116) );
  NOR2X2 U32 ( .A(A[26]), .B(B[26]), .Y(n117) );
  NOR2X2 U33 ( .A(n44), .B(n43), .Y(n210) );
  INVX4 U34 ( .A(n186), .Y(n181) );
  NAND2X2 U35 ( .A(n157), .B(n137), .Y(n138) );
  NAND3X2 U36 ( .A(A[24]), .B(B[24]), .C(n119), .Y(n132) );
  OR2X2 U37 ( .A(A[6]), .B(B[6]), .Y(n61) );
  NOR2BX1 U38 ( .AN(n169), .B(n173), .Y(n172) );
  INVX1 U39 ( .A(n171), .Y(n173) );
  INVX4 U40 ( .A(n185), .Y(n182) );
  INVX4 U41 ( .A(n203), .Y(n202) );
  INVX4 U42 ( .A(n189), .Y(n183) );
  AND2X2 U43 ( .A(n167), .B(n157), .Y(n168) );
  NAND2X1 U44 ( .A(B[10]), .B(A[10]), .Y(n245) );
  INVX1 U45 ( .A(n41), .Y(n16) );
  BUFX3 U46 ( .A(n43), .Y(n14) );
  INVX1 U47 ( .A(n259), .Y(n56) );
  AOI21X2 U48 ( .A0(n63), .A1(n34), .B0(n35), .Y(n33) );
  NAND2X1 U49 ( .A(B[5]), .B(A[5]), .Y(n62) );
  NAND2X1 U50 ( .A(B[4]), .B(A[4]), .Y(n66) );
  NAND2X1 U51 ( .A(B[0]), .B(A[0]), .Y(n196) );
  NAND2X1 U52 ( .A(n98), .B(n84), .Y(n110) );
  XOR2X1 U53 ( .A(B[31]), .B(A[31]), .Y(n77) );
  NOR2BX2 U54 ( .AN(n104), .B(n118), .Y(n126) );
  CLKBUFX8 U55 ( .A(n265), .Y(SUM[22]) );
  XOR2X2 U56 ( .A(n46), .B(n47), .Y(SUM[9]) );
  NOR2BX1 U57 ( .AN(n51), .B(n52), .Y(n50) );
  INVX1 U58 ( .A(n226), .Y(n235) );
  NOR2BX2 U59 ( .AN(n135), .B(n140), .Y(n161) );
  NOR2X2 U60 ( .A(n29), .B(n100), .Y(n95) );
  NOR2BX1 U61 ( .AN(n215), .B(n41), .Y(n234) );
  XOR2X1 U62 ( .A(n68), .B(n69), .Y(SUM[3]) );
  OAI21X1 U63 ( .A0(n72), .A1(n73), .B0(n74), .Y(n68) );
  XOR2X1 U64 ( .A(n75), .B(n105), .Y(SUM[2]) );
  NAND2X2 U65 ( .A(n205), .B(n184), .Y(n203) );
  NOR2BX2 U66 ( .AN(n184), .B(n207), .Y(n206) );
  OR2X2 U67 ( .A(A[26]), .B(B[26]), .Y(n91) );
  XOR2X1 U68 ( .A(n63), .B(n64), .Y(SUM[5]) );
  NAND2X2 U69 ( .A(B[9]), .B(A[9]), .Y(n8) );
  AND2X2 U70 ( .A(B[26]), .B(A[26]), .Y(n9) );
  NAND2X4 U71 ( .A(B[14]), .B(A[14]), .Y(n216) );
  INVX1 U72 ( .A(n225), .Y(n218) );
  NAND2X1 U73 ( .A(B[30]), .B(A[30]), .Y(n79) );
  NOR2X4 U74 ( .A(A[15]), .B(B[15]), .Y(n44) );
  OR2X4 U75 ( .A(A[15]), .B(B[15]), .Y(n42) );
  AND2X4 U76 ( .A(n128), .B(n91), .Y(n36) );
  NAND2X2 U77 ( .A(A[16]), .B(B[16]), .Y(n184) );
  CLKINVX3 U78 ( .A(n188), .Y(n207) );
  NAND2X4 U79 ( .A(n10), .B(n219), .Y(n208) );
  AND3X4 U80 ( .A(n42), .B(n226), .C(n227), .Y(n10) );
  NAND3X4 U81 ( .A(n174), .B(n175), .C(n176), .Y(n170) );
  NAND3X2 U82 ( .A(n175), .B(n174), .C(n176), .Y(n17) );
  XOR2X4 U83 ( .A(n164), .B(n165), .Y(n265) );
  OAI2BB1X4 U84 ( .A0N(n120), .A1N(n121), .B0(n147), .Y(n151) );
  XNOR2X4 U85 ( .A(n160), .B(n11), .Y(SUM[23]) );
  CLKINVX3 U86 ( .A(n46), .Y(n254) );
  XOR2X2 U87 ( .A(n251), .B(n253), .Y(SUM[10]) );
  NAND3X4 U88 ( .A(A[20]), .B(n18), .C(n157), .Y(n156) );
  NOR2X1 U89 ( .A(n138), .B(n19), .Y(n133) );
  OAI2BB1X4 U90 ( .A0N(n226), .A1N(n236), .B0(n214), .Y(n233) );
  XOR2X4 U91 ( .A(n199), .B(n201), .Y(SUM[18]) );
  NAND2X2 U92 ( .A(B[23]), .B(A[23]), .Y(n135) );
  NAND4X4 U93 ( .A(n12), .B(n185), .C(n15), .D(n187), .Y(n175) );
  AND2X4 U94 ( .A(n188), .B(n189), .Y(n12) );
  CLKINVX4 U95 ( .A(n180), .Y(n179) );
  NAND2X1 U96 ( .A(B[19]), .B(A[19]), .Y(n180) );
  NAND2X4 U97 ( .A(n208), .B(n209), .Y(n13) );
  XOR2X1 U98 ( .A(n13), .B(n206), .Y(SUM[16]) );
  OAI2BB1X4 U99 ( .A0N(n233), .A1N(n16), .B0(n215), .Y(n231) );
  CLKBUFX3 U100 ( .A(B[21]), .Y(n20) );
  NAND2XL U101 ( .A(B[26]), .B(A[26]), .Y(n128) );
  NAND2X2 U102 ( .A(B[17]), .B(A[17]), .Y(n193) );
  AOI21X4 U103 ( .A0(n20), .A1(A[21]), .B0(n158), .Y(n155) );
  BUFX4 U104 ( .A(B[20]), .Y(n18) );
  NAND2X4 U105 ( .A(n170), .B(n171), .Y(n19) );
  NOR2X4 U106 ( .A(n43), .B(n41), .Y(n227) );
  NOR2BXL U107 ( .AN(n216), .B(n14), .Y(n232) );
  INVX4 U108 ( .A(n159), .Y(n158) );
  NAND2X2 U109 ( .A(B[25]), .B(A[25]), .Y(n124) );
  NOR2BX1 U110 ( .AN(n193), .B(n183), .Y(n204) );
  NAND2X4 U111 ( .A(B[8]), .B(A[8]), .Y(n51) );
  AOI21X4 U112 ( .A0(n190), .A1(n185), .B0(n191), .Y(n174) );
  NAND2X2 U113 ( .A(B[2]), .B(A[2]), .Y(n74) );
  OR2X2 U114 ( .A(B[2]), .B(A[2]), .Y(n106) );
  INVX4 U115 ( .A(n154), .Y(n140) );
  INVX2 U116 ( .A(n75), .Y(n72) );
  INVX4 U117 ( .A(n106), .Y(n73) );
  XOR2X2 U118 ( .A(n166), .B(n168), .Y(SUM[21]) );
  INVX4 U119 ( .A(n222), .Y(n65) );
  INVX3 U120 ( .A(n213), .Y(n212) );
  NAND2X2 U121 ( .A(B[15]), .B(A[15]), .Y(n213) );
  NOR2X4 U122 ( .A(n181), .B(n193), .Y(n190) );
  NAND2X4 U123 ( .A(B[13]), .B(A[13]), .Y(n215) );
  NAND2BX2 U124 ( .AN(n40), .B(n79), .Y(n93) );
  OR2X4 U125 ( .A(n65), .B(n225), .Y(n21) );
  NAND2X4 U126 ( .A(n21), .B(n224), .Y(n49) );
  NAND2X4 U127 ( .A(n49), .B(n248), .Y(n255) );
  NAND2X1 U128 ( .A(A[18]), .B(B[18]), .Y(n192) );
  NAND2X4 U129 ( .A(n249), .B(n23), .Y(n24) );
  NAND2X4 U130 ( .A(n22), .B(n250), .Y(n25) );
  NAND2X4 U131 ( .A(n24), .B(n25), .Y(SUM[11]) );
  CLKINVX3 U132 ( .A(n249), .Y(n22) );
  INVX2 U133 ( .A(n250), .Y(n23) );
  NAND2X4 U134 ( .A(n26), .B(n27), .Y(n28) );
  NAND2X4 U135 ( .A(n28), .B(n221), .Y(n236) );
  CLKINVX3 U136 ( .A(n238), .Y(n26) );
  CLKINVX3 U137 ( .A(n217), .Y(n27) );
  NAND4BBX4 U138 ( .AN(n52), .BN(n48), .C(n242), .D(n241), .Y(n217) );
  XOR2X2 U139 ( .A(n236), .B(n237), .Y(SUM[12]) );
  NAND2X4 U140 ( .A(n18), .B(A[20]), .Y(n169) );
  AND2X2 U141 ( .A(n99), .B(n86), .Y(n29) );
  NOR2X2 U142 ( .A(n90), .B(n102), .Y(n99) );
  NAND2X2 U143 ( .A(n98), .B(n101), .Y(n100) );
  NOR2X4 U144 ( .A(n95), .B(n96), .Y(n94) );
  NOR2X4 U145 ( .A(A[14]), .B(B[14]), .Y(n43) );
  NAND2X4 U146 ( .A(B[29]), .B(A[29]), .Y(n84) );
  NAND2X2 U147 ( .A(n20), .B(A[21]), .Y(n167) );
  NAND2X2 U148 ( .A(B[24]), .B(A[24]), .Y(n147) );
  OAI211X2 U149 ( .A0(n41), .A1(n214), .B0(n215), .C0(n216), .Y(n211) );
  NOR2X4 U150 ( .A(A[13]), .B(B[13]), .Y(n41) );
  OR2X2 U151 ( .A(B[27]), .B(A[27]), .Y(n39) );
  OAI21X2 U152 ( .A0(n80), .A1(n81), .B0(n82), .Y(n78) );
  AOI21X2 U153 ( .A0(n85), .A1(n86), .B0(n87), .Y(n80) );
  INVX4 U154 ( .A(n137), .Y(n163) );
  NOR2X2 U155 ( .A(n83), .B(n40), .Y(n82) );
  NOR2X2 U156 ( .A(A[30]), .B(B[30]), .Y(n40) );
  NAND2X4 U157 ( .A(n255), .B(n51), .Y(n46) );
  NAND2X4 U158 ( .A(n8), .B(n51), .Y(n244) );
  OAI21X2 U159 ( .A0(n33), .A1(n57), .B0(n58), .Y(n53) );
  NAND3BX2 U160 ( .AN(n133), .B(n134), .C(n135), .Y(n130) );
  NAND2X4 U161 ( .A(n135), .B(n150), .Y(n149) );
  AOI21X4 U162 ( .A0(n242), .A1(n251), .B0(n252), .Y(n250) );
  OAI21X4 U163 ( .A0(n254), .A1(n48), .B0(n8), .Y(n251) );
  NAND2X4 U164 ( .A(B[1]), .B(A[1]), .Y(n109) );
  OR2X4 U165 ( .A(A[1]), .B(B[1]), .Y(n107) );
  XOR2X4 U166 ( .A(n53), .B(n54), .Y(SUM[7]) );
  OR2X4 U167 ( .A(A[3]), .B(B[3]), .Y(n260) );
  NAND2X1 U168 ( .A(B[3]), .B(A[3]), .Y(n70) );
  NOR2X2 U169 ( .A(A[5]), .B(B[5]), .Y(n37) );
  NOR3BX4 U170 ( .AN(n154), .B(n19), .C(n138), .Y(n148) );
  NAND2X1 U171 ( .A(B[6]), .B(A[6]), .Y(n58) );
  OAI2BB1X1 U172 ( .A0N(n107), .A1N(n108), .B0(n109), .Y(n75) );
  OAI2BB1X4 U173 ( .A0N(n157), .A1N(n166), .B0(n167), .Y(n164) );
  INVXL U174 ( .A(n62), .Y(n35) );
  INVX2 U175 ( .A(n98), .Y(n83) );
  INVXL U176 ( .A(n92), .Y(n88) );
  NAND3X1 U177 ( .A(n242), .B(n243), .C(n244), .Y(n240) );
  XOR2X2 U178 ( .A(n231), .B(n232), .Y(SUM[14]) );
  NOR2BX1 U179 ( .AN(n159), .B(n163), .Y(n165) );
  NAND3X4 U180 ( .A(n119), .B(n120), .C(n121), .Y(n31) );
  NAND3X4 U181 ( .A(n39), .B(n91), .C(n92), .Y(n103) );
  OAI21X4 U182 ( .A0(n261), .A1(n262), .B0(n70), .Y(n222) );
  NOR2X2 U183 ( .A(n263), .B(n264), .Y(n261) );
  NAND2X4 U184 ( .A(n106), .B(n260), .Y(n262) );
  CLKINVX3 U185 ( .A(n74), .Y(n263) );
  NOR2BX1 U186 ( .AN(n55), .B(n56), .Y(n54) );
  OAI21X2 U187 ( .A0(n195), .A1(n196), .B0(n109), .Y(n264) );
  INVXL U188 ( .A(n245), .Y(n252) );
  NOR2BXL U189 ( .AN(n109), .B(n195), .Y(n194) );
  NAND3BX4 U190 ( .AN(n148), .B(n135), .C(n150), .Y(n121) );
  AND2X1 U191 ( .A(n124), .B(n119), .Y(n152) );
  AND2X1 U192 ( .A(n245), .B(n242), .Y(n253) );
  INVX4 U193 ( .A(n231), .Y(n230) );
  INVXL U194 ( .A(n260), .Y(n71) );
  INVX4 U195 ( .A(n243), .Y(n48) );
  INVX1 U196 ( .A(n37), .Y(n34) );
  XOR2X2 U197 ( .A(n76), .B(n77), .Y(SUM[31]) );
  AOI2BB1X2 U198 ( .A0N(n88), .A1N(n89), .B0(n90), .Y(n85) );
  NAND2BX4 U199 ( .AN(n31), .B(n116), .Y(n86) );
  OAI2BB1X4 U200 ( .A0N(n122), .A1N(n119), .B0(n123), .Y(n92) );
  NOR2BX1 U201 ( .AN(n196), .B(n32), .Y(SUM[0]) );
  NOR2XL U202 ( .A(A[0]), .B(B[0]), .Y(n32) );
  OAI21X4 U203 ( .A0(n38), .A1(n65), .B0(n66), .Y(n63) );
  AOI21X1 U204 ( .A0(n218), .A1(n222), .B0(n223), .Y(n220) );
  NOR2BX1 U205 ( .AN(n214), .B(n235), .Y(n237) );
  XOR2X1 U206 ( .A(n49), .B(n50), .Y(SUM[8]) );
  NOR2BX1 U207 ( .AN(n192), .B(n182), .Y(n201) );
  XOR2X1 U208 ( .A(n233), .B(n234), .Y(n267) );
  NOR2BX1 U209 ( .AN(n62), .B(n37), .Y(n64) );
  NOR2BX1 U210 ( .AN(n8), .B(n48), .Y(n47) );
  NAND2XL U211 ( .A(n180), .B(n186), .Y(n197) );
  INVXL U212 ( .A(n192), .Y(n200) );
  NAND2XL U213 ( .A(n241), .B(n247), .Y(n249) );
  XOR2X1 U214 ( .A(n222), .B(n67), .Y(SUM[4]) );
  NOR2BX1 U215 ( .AN(n66), .B(n38), .Y(n67) );
  INVX1 U216 ( .A(n114), .Y(n113) );
  XNOR2X4 U217 ( .A(n36), .B(n142), .Y(SUM[26]) );
  INVXL U218 ( .A(n61), .Y(n57) );
  INVX1 U219 ( .A(n104), .Y(n90) );
  INVX1 U220 ( .A(n107), .Y(n195) );
  XOR2X2 U221 ( .A(n121), .B(n153), .Y(SUM[24]) );
  OAI21X2 U222 ( .A0(n83), .A1(n97), .B0(n84), .Y(n96) );
  NOR2BX1 U223 ( .AN(n213), .B(n44), .Y(n229) );
  NAND3X2 U224 ( .A(n257), .B(n58), .C(n55), .Y(n256) );
  NAND3BX2 U225 ( .AN(n37), .B(n258), .C(n61), .Y(n257) );
  NOR2BX2 U226 ( .AN(n245), .B(n246), .Y(n239) );
  NAND2XL U227 ( .A(n136), .B(n137), .Y(n134) );
  NOR2BX1 U228 ( .AN(n70), .B(n71), .Y(n69) );
  NOR2BX1 U229 ( .AN(n74), .B(n73), .Y(n105) );
  XOR2X1 U230 ( .A(n108), .B(n194), .Y(SUM[1]) );
  INVX1 U231 ( .A(n196), .Y(n108) );
  NAND2X2 U232 ( .A(n78), .B(n79), .Y(n76) );
  NAND2X2 U233 ( .A(B[12]), .B(A[12]), .Y(n214) );
  NAND2X1 U234 ( .A(B[7]), .B(A[7]), .Y(n55) );
  NAND2XL U235 ( .A(B[28]), .B(A[28]), .Y(n114) );
  NAND2XL U236 ( .A(A[28]), .B(B[28]), .Y(n97) );
  OAI2BB1X1 U237 ( .A0N(B[28]), .A1N(A[28]), .B0(n84), .Y(n81) );
  NAND2X4 U238 ( .A(n208), .B(n209), .Y(n187) );
  NAND2X4 U239 ( .A(n13), .B(n188), .Y(n205) );
  OAI21X2 U240 ( .A0(n220), .A1(n217), .B0(n221), .Y(n219) );
  XOR2X1 U241 ( .A(n170), .B(n172), .Y(n266) );
  NAND2X2 U242 ( .A(n120), .B(n119), .Y(n141) );
  NAND2X2 U243 ( .A(B[11]), .B(A[11]), .Y(n247) );
  OAI21XL U244 ( .A0(B[27]), .A1(A[27]), .B0(n91), .Y(n89) );
  XNOR2X4 U245 ( .A(n202), .B(n204), .Y(SUM[17]) );
  INVX4 U246 ( .A(n164), .Y(n162) );
  AND2X1 U247 ( .A(A[24]), .B(B[24]), .Y(n122) );
  XOR2X4 U248 ( .A(n93), .B(n94), .Y(SUM[30]) );
  XOR2X4 U249 ( .A(n111), .B(n110), .Y(SUM[29]) );
  OR2X4 U250 ( .A(A[29]), .B(B[29]), .Y(n98) );
  XOR2X4 U251 ( .A(n112), .B(n115), .Y(SUM[28]) );
  NOR2BX4 U252 ( .AN(n114), .B(n87), .Y(n115) );
  CLKINVX3 U253 ( .A(n101), .Y(n87) );
  OR2X4 U254 ( .A(A[28]), .B(B[28]), .Y(n101) );
  NOR2BX4 U255 ( .AN(n124), .B(n9), .Y(n123) );
  XOR2X4 U256 ( .A(n125), .B(n126), .Y(SUM[27]) );
  NAND2X4 U257 ( .A(B[27]), .B(A[27]), .Y(n104) );
  OAI21X4 U258 ( .A0(n127), .A1(n117), .B0(n128), .Y(n125) );
  AOI21X4 U259 ( .A0(n129), .A1(n130), .B0(n131), .Y(n127) );
  NAND2BX4 U260 ( .AN(n144), .B(n132), .Y(n131) );
  NOR2X4 U261 ( .A(n140), .B(n141), .Y(n129) );
  CLKINVX3 U262 ( .A(n124), .Y(n144) );
  XOR2X4 U263 ( .A(n151), .B(n152), .Y(SUM[25]) );
  OR2X4 U264 ( .A(B[25]), .B(A[25]), .Y(n119) );
  OR2X4 U265 ( .A(A[24]), .B(B[24]), .Y(n120) );
  NAND3X4 U266 ( .A(n137), .B(n154), .C(n136), .Y(n150) );
  NAND2X4 U267 ( .A(n155), .B(n156), .Y(n136) );
  OR2X4 U268 ( .A(B[23]), .B(A[23]), .Y(n154) );
  OAI21X4 U269 ( .A0(n162), .A1(n163), .B0(n159), .Y(n160) );
  OR2X4 U270 ( .A(B[22]), .B(A[22]), .Y(n137) );
  NAND2X4 U271 ( .A(A[22]), .B(B[22]), .Y(n159) );
  OR2X4 U272 ( .A(B[21]), .B(A[21]), .Y(n157) );
  NAND2X4 U273 ( .A(n139), .B(n169), .Y(n166) );
  NAND2X4 U274 ( .A(n17), .B(n171), .Y(n139) );
  OR2X4 U275 ( .A(A[20]), .B(B[20]), .Y(n171) );
  AOI21X4 U276 ( .A0(n178), .A1(n177), .B0(n179), .Y(n176) );
  NOR2X4 U277 ( .A(n181), .B(n182), .Y(n178) );
  NOR2X4 U278 ( .A(n183), .B(n184), .Y(n177) );
  XOR2X4 U279 ( .A(n198), .B(n197), .Y(SUM[19]) );
  AOI21X4 U280 ( .A0(n199), .A1(n185), .B0(n200), .Y(n198) );
  OR2X4 U281 ( .A(B[19]), .B(A[19]), .Y(n186) );
  OR2X4 U282 ( .A(B[18]), .B(A[18]), .Y(n185) );
  OAI21X4 U283 ( .A0(n202), .A1(n183), .B0(n193), .Y(n199) );
  OR2X4 U284 ( .A(B[16]), .B(A[16]), .Y(n188) );
  AOI21X4 U285 ( .A0(n210), .A1(n211), .B0(n212), .Y(n209) );
  XOR2X4 U286 ( .A(n228), .B(n229), .Y(SUM[15]) );
  OAI21X4 U287 ( .A0(n230), .A1(n14), .B0(n216), .Y(n228) );
  OR2X4 U288 ( .A(A[12]), .B(B[12]), .Y(n226) );
  OAI2BB1X4 U289 ( .A0N(n239), .A1N(n240), .B0(n241), .Y(n221) );
  CLKINVX3 U290 ( .A(n247), .Y(n246) );
  CLKINVX3 U291 ( .A(n248), .Y(n52) );
  OR2X4 U292 ( .A(B[11]), .B(A[11]), .Y(n241) );
  OR2X4 U293 ( .A(A[10]), .B(B[10]), .Y(n242) );
  OR2X4 U294 ( .A(A[9]), .B(B[9]), .Y(n243) );
  OR2X4 U295 ( .A(A[8]), .B(B[8]), .Y(n248) );
  NAND2BX4 U296 ( .AN(n56), .B(n256), .Y(n224) );
  OR2X4 U297 ( .A(A[7]), .B(B[7]), .Y(n259) );
endmodule


module hash_core_DW01_add_27 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n267, n268, n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266;

  CLKINVX3 U2 ( .A(n166), .Y(n12) );
  NOR2X4 U3 ( .A(n149), .B(n148), .Y(n146) );
  NAND2X4 U4 ( .A(n1), .B(n2), .Y(n3) );
  NAND2X4 U5 ( .A(n3), .B(n216), .Y(n229) );
  INVX4 U6 ( .A(n231), .Y(n1) );
  INVX20 U7 ( .A(n43), .Y(n2) );
  NAND2X4 U8 ( .A(B[14]), .B(A[14]), .Y(n216) );
  NAND2X1 U9 ( .A(B[10]), .B(A[10]), .Y(n247) );
  NAND2X2 U10 ( .A(n187), .B(n186), .Y(n4) );
  NAND3X4 U11 ( .A(n5), .B(n188), .C(n19), .Y(n176) );
  CLKINVX3 U12 ( .A(n4), .Y(n5) );
  AND2X2 U13 ( .A(n189), .B(n190), .Y(n19) );
  NAND3X1 U14 ( .A(n175), .B(n176), .C(n177), .Y(n171) );
  NOR2BXL U15 ( .AN(n8), .B(n47), .Y(n46) );
  NAND2X4 U16 ( .A(n8), .B(n50), .Y(n246) );
  XOR2X2 U17 ( .A(n45), .B(n46), .Y(SUM[9]) );
  OR2X4 U18 ( .A(A[7]), .B(B[7]), .Y(n261) );
  NAND2X2 U19 ( .A(B[7]), .B(A[7]), .Y(n54) );
  NAND2X2 U20 ( .A(B[29]), .B(A[29]), .Y(n83) );
  INVX2 U21 ( .A(n268), .Y(n6) );
  CLKINVX4 U22 ( .A(n6), .Y(SUM[12]) );
  INVX8 U23 ( .A(n223), .Y(n64) );
  OAI21X4 U24 ( .A0(n263), .A1(n264), .B0(n69), .Y(n223) );
  OAI21X1 U25 ( .A0(n79), .A1(n80), .B0(n81), .Y(n77) );
  INVX1 U26 ( .A(n227), .Y(n236) );
  INVX2 U27 ( .A(n156), .Y(n139) );
  INVX1 U28 ( .A(n167), .Y(n14) );
  INVX4 U29 ( .A(n187), .Y(n182) );
  AOI2BB1X1 U30 ( .A0N(n87), .A1N(n88), .B0(n89), .Y(n84) );
  OR2X2 U31 ( .A(A[1]), .B(B[1]), .Y(n106) );
  OR2X2 U32 ( .A(A[8]), .B(B[8]), .Y(n250) );
  NOR2BX2 U33 ( .AN(n247), .B(n248), .Y(n241) );
  OR2X2 U34 ( .A(A[12]), .B(B[12]), .Y(n227) );
  INVX1 U35 ( .A(n73), .Y(n265) );
  AOI21X2 U36 ( .A0(B[21]), .A1(A[21]), .B0(n160), .Y(n157) );
  NAND3X2 U37 ( .A(A[20]), .B(B[20]), .C(n159), .Y(n158) );
  INVX2 U38 ( .A(n161), .Y(n160) );
  INVX1 U39 ( .A(n261), .Y(n55) );
  NAND2X1 U40 ( .A(A[0]), .B(B[0]), .Y(n197) );
  NAND2X1 U41 ( .A(B[1]), .B(A[1]), .Y(n108) );
  NOR2X2 U42 ( .A(A[15]), .B(B[15]), .Y(n40) );
  INVX1 U43 ( .A(n42), .Y(n15) );
  INVX1 U44 ( .A(n250), .Y(n51) );
  NOR2BX1 U45 ( .AN(n194), .B(n184), .Y(n205) );
  NOR2BX1 U46 ( .AN(n170), .B(n174), .Y(n173) );
  INVX1 U47 ( .A(n172), .Y(n174) );
  BUFX3 U48 ( .A(n38), .Y(n31) );
  OR2X2 U49 ( .A(A[3]), .B(B[3]), .Y(n262) );
  NAND2X1 U50 ( .A(B[2]), .B(A[2]), .Y(n73) );
  NAND2X1 U51 ( .A(n97), .B(n100), .Y(n99) );
  XOR2X1 U52 ( .A(B[31]), .B(A[31]), .Y(n76) );
  NOR2BX1 U53 ( .AN(n161), .B(n164), .Y(n165) );
  INVX2 U54 ( .A(n13), .Y(n21) );
  BUFX3 U55 ( .A(n267), .Y(SUM[13]) );
  XOR2X2 U56 ( .A(n200), .B(n202), .Y(SUM[18]) );
  INVX1 U57 ( .A(n247), .Y(n254) );
  XOR2X1 U58 ( .A(n238), .B(n239), .Y(n268) );
  NOR2BX1 U59 ( .AN(n214), .B(n236), .Y(n239) );
  AND2X2 U60 ( .A(n247), .B(n244), .Y(n255) );
  NOR2BX1 U61 ( .AN(n65), .B(n29), .Y(n66) );
  NOR2BX2 U62 ( .AN(n103), .B(n127), .Y(n126) );
  NAND2X1 U63 ( .A(n124), .B(n90), .Y(n141) );
  INVX1 U64 ( .A(n152), .Y(n24) );
  NOR2BX2 U65 ( .AN(n30), .B(n139), .Y(n163) );
  OAI21X2 U66 ( .A0(n13), .A1(n164), .B0(n161), .Y(n162) );
  XOR2X2 U67 ( .A(n58), .B(n59), .Y(SUM[6]) );
  INVX1 U68 ( .A(n34), .Y(n58) );
  NOR2BX1 U69 ( .AN(n54), .B(n55), .Y(n53) );
  OR2X2 U70 ( .A(A[26]), .B(B[26]), .Y(n90) );
  NOR2X1 U71 ( .A(A[26]), .B(B[26]), .Y(n116) );
  NAND2X2 U72 ( .A(B[9]), .B(A[9]), .Y(n8) );
  INVX1 U73 ( .A(n118), .Y(n153) );
  NAND2X1 U74 ( .A(B[5]), .B(A[5]), .Y(n61) );
  AND2X2 U75 ( .A(n57), .B(n54), .Y(n9) );
  NAND2X2 U76 ( .A(B[17]), .B(A[17]), .Y(n194) );
  AND2X2 U77 ( .A(n103), .B(n102), .Y(n10) );
  NAND3X2 U78 ( .A(n136), .B(n156), .C(n135), .Y(n11) );
  AOI21X4 U79 ( .A0(n166), .A1(n159), .B0(n14), .Y(n13) );
  NAND2X4 U80 ( .A(n188), .B(n189), .Y(n206) );
  NAND2X2 U81 ( .A(B[16]), .B(A[16]), .Y(n185) );
  INVX3 U82 ( .A(n48), .Y(n240) );
  NOR2XL U83 ( .A(B[27]), .B(A[27]), .Y(n117) );
  NOR2X1 U84 ( .A(B[27]), .B(A[27]), .Y(n32) );
  OAI21XL U85 ( .A0(B[27]), .A1(A[27]), .B0(n90), .Y(n88) );
  NAND2X2 U86 ( .A(B[27]), .B(A[27]), .Y(n103) );
  AOI21X1 U87 ( .A0(n84), .A1(n85), .B0(n86), .Y(n79) );
  AOI21X2 U88 ( .A0(n98), .A1(n85), .B0(n99), .Y(n94) );
  OAI2BB1X4 U89 ( .A0N(n234), .A1N(n15), .B0(n215), .Y(n232) );
  BUFX4 U90 ( .A(B[4]), .Y(n16) );
  AOI21X2 U91 ( .A0(n218), .A1(n223), .B0(n224), .Y(n221) );
  XOR2X1 U92 ( .A(n48), .B(n49), .Y(SUM[8]) );
  AOI21X4 U93 ( .A0(n210), .A1(n211), .B0(n212), .Y(n209) );
  NOR2BXL U94 ( .AN(n50), .B(n51), .Y(n49) );
  CLKINVX8 U95 ( .A(n119), .Y(n145) );
  OR2X4 U96 ( .A(A[24]), .B(B[24]), .Y(n119) );
  XOR2X1 U97 ( .A(n188), .B(n207), .Y(SUM[16]) );
  NOR2BX2 U98 ( .AN(n113), .B(n86), .Y(n114) );
  INVX1 U99 ( .A(n100), .Y(n86) );
  NOR2BX1 U100 ( .AN(n216), .B(n43), .Y(n233) );
  NAND2X4 U101 ( .A(n17), .B(n115), .Y(n85) );
  AND3X2 U102 ( .A(n118), .B(n119), .C(n120), .Y(n17) );
  NAND3X2 U103 ( .A(n44), .B(n227), .C(n228), .Y(n219) );
  NOR2X2 U104 ( .A(n43), .B(n42), .Y(n228) );
  NAND2X2 U105 ( .A(B[30]), .B(A[30]), .Y(n78) );
  AOI21X4 U106 ( .A0(n244), .A1(n253), .B0(n254), .Y(n252) );
  NAND3X4 U107 ( .A(n175), .B(n176), .C(n177), .Y(n18) );
  NAND2X4 U108 ( .A(B[26]), .B(A[26]), .Y(n124) );
  XOR2X1 U109 ( .A(n171), .B(n173), .Y(SUM[20]) );
  INVX1 U110 ( .A(n120), .Y(n154) );
  INVX2 U111 ( .A(n123), .Y(n144) );
  NAND2X2 U112 ( .A(n119), .B(n118), .Y(n140) );
  NAND3X2 U113 ( .A(n20), .B(n133), .C(n30), .Y(n130) );
  OR2X1 U114 ( .A(n137), .B(n138), .Y(n20) );
  BUFX8 U115 ( .A(n39), .Y(n29) );
  NOR2X1 U116 ( .A(A[4]), .B(n16), .Y(n39) );
  AOI21X4 U117 ( .A0(n62), .A1(n35), .B0(n36), .Y(n34) );
  OAI21X4 U118 ( .A0(n29), .A1(n64), .B0(n65), .Y(n62) );
  OAI21X4 U119 ( .A0(n203), .A1(n184), .B0(n194), .Y(n22) );
  CLKINVX8 U120 ( .A(n204), .Y(n203) );
  NOR2BXL U121 ( .AN(n215), .B(n42), .Y(n235) );
  NAND2X2 U122 ( .A(B[25]), .B(A[25]), .Y(n123) );
  OAI2BB1X4 U123 ( .A0N(n119), .A1N(n120), .B0(n28), .Y(n151) );
  OR2X2 U124 ( .A(A[2]), .B(B[2]), .Y(n105) );
  XOR2X4 U125 ( .A(n251), .B(n252), .Y(SUM[11]) );
  NAND2X4 U126 ( .A(n250), .B(n48), .Y(n257) );
  NAND2BXL U127 ( .AN(n41), .B(n78), .Y(n92) );
  NOR2X2 U128 ( .A(n40), .B(n43), .Y(n210) );
  NAND2X2 U129 ( .A(n77), .B(n78), .Y(n75) );
  NAND2X2 U130 ( .A(n151), .B(n24), .Y(n25) );
  NAND2X4 U131 ( .A(n23), .B(n152), .Y(n26) );
  NAND2X4 U132 ( .A(n25), .B(n26), .Y(SUM[25]) );
  INVX4 U133 ( .A(n151), .Y(n23) );
  NAND2X4 U134 ( .A(n10), .B(n85), .Y(n111) );
  NAND2X4 U135 ( .A(B[20]), .B(A[20]), .Y(n170) );
  NAND2X4 U136 ( .A(n9), .B(n259), .Y(n258) );
  NAND3BX2 U137 ( .AN(n31), .B(n260), .C(n60), .Y(n259) );
  NAND2X1 U138 ( .A(B[6]), .B(A[6]), .Y(n57) );
  NOR2X4 U139 ( .A(n94), .B(n95), .Y(n93) );
  OAI21X2 U140 ( .A0(n82), .A1(n96), .B0(n83), .Y(n95) );
  NAND4BBX4 U141 ( .AN(n51), .BN(n47), .C(n244), .D(n243), .Y(n217) );
  NOR2X2 U142 ( .A(n89), .B(n101), .Y(n98) );
  BUFX8 U143 ( .A(n147), .Y(n28) );
  INVX8 U144 ( .A(n190), .Y(n184) );
  NAND4BBX2 U145 ( .AN(n31), .BN(n29), .C(n60), .D(n261), .Y(n226) );
  OAI21X4 U146 ( .A0(n64), .A1(n226), .B0(n225), .Y(n48) );
  XOR2X2 U147 ( .A(n62), .B(n63), .Y(SUM[5]) );
  NAND2X2 U148 ( .A(B[4]), .B(A[4]), .Y(n65) );
  OAI21X2 U149 ( .A0(n34), .A1(n56), .B0(n57), .Y(n52) );
  NAND2BX4 U150 ( .AN(n219), .B(n220), .Y(n208) );
  OAI21X2 U151 ( .A0(n221), .A1(n217), .B0(n222), .Y(n220) );
  INVX4 U152 ( .A(n136), .Y(n164) );
  AOI21X4 U153 ( .A0(n186), .A1(n22), .B0(n201), .Y(n199) );
  OAI21X4 U154 ( .A0(n203), .A1(n184), .B0(n194), .Y(n200) );
  XOR2X4 U155 ( .A(n92), .B(n93), .Y(SUM[30]) );
  NAND2X2 U156 ( .A(B[13]), .B(A[13]), .Y(n215) );
  BUFX8 U157 ( .A(n134), .Y(n30) );
  XOR2X4 U158 ( .A(n75), .B(n76), .Y(SUM[31]) );
  NOR2X4 U159 ( .A(B[14]), .B(A[14]), .Y(n43) );
  NAND2X2 U160 ( .A(B[15]), .B(A[15]), .Y(n213) );
  OR2X4 U161 ( .A(A[15]), .B(B[15]), .Y(n44) );
  OAI211X2 U162 ( .A0(n42), .A1(n214), .B0(n215), .C0(n216), .Y(n211) );
  NOR2X4 U163 ( .A(A[13]), .B(B[13]), .Y(n42) );
  NOR2XL U164 ( .A(A[5]), .B(B[5]), .Y(n38) );
  NAND2X2 U165 ( .A(B[8]), .B(A[8]), .Y(n50) );
  XOR2X4 U166 ( .A(n52), .B(n53), .Y(SUM[7]) );
  NAND2X1 U167 ( .A(B[3]), .B(A[3]), .Y(n69) );
  NAND2X4 U168 ( .A(B[12]), .B(A[12]), .Y(n214) );
  OR2X4 U169 ( .A(A[17]), .B(B[17]), .Y(n190) );
  NOR2X2 U170 ( .A(A[30]), .B(B[30]), .Y(n41) );
  OR2X2 U171 ( .A(A[6]), .B(B[6]), .Y(n60) );
  INVXL U172 ( .A(n61), .Y(n36) );
  XOR2X2 U173 ( .A(n154), .B(n155), .Y(n37) );
  NAND3BX2 U174 ( .AN(n32), .B(n90), .C(n91), .Y(n102) );
  AND2X2 U175 ( .A(A[24]), .B(B[24]), .Y(n121) );
  OAI2BB1XL U176 ( .A0N(n106), .A1N(n107), .B0(n108), .Y(n74) );
  NOR2X4 U177 ( .A(n184), .B(n185), .Y(n178) );
  CLKINVX3 U178 ( .A(n181), .Y(n180) );
  INVX4 U179 ( .A(n37), .Y(SUM[24]) );
  AND2X2 U180 ( .A(n123), .B(n124), .Y(n122) );
  NOR2X2 U181 ( .A(n265), .B(n266), .Y(n263) );
  NAND2X4 U182 ( .A(n105), .B(n262), .Y(n264) );
  NOR2BXL U183 ( .AN(n57), .B(n56), .Y(n59) );
  INVXL U184 ( .A(n262), .Y(n70) );
  AND2X1 U185 ( .A(n185), .B(n189), .Y(n207) );
  INVXL U186 ( .A(n159), .Y(n169) );
  INVXL U187 ( .A(n193), .Y(n201) );
  NAND3X1 U188 ( .A(n244), .B(n245), .C(n246), .Y(n242) );
  INVX1 U189 ( .A(n31), .Y(n35) );
  OAI21X1 U190 ( .A0(n196), .A1(n197), .B0(n108), .Y(n266) );
  NOR2BXL U191 ( .AN(n108), .B(n196), .Y(n195) );
  NAND2XL U192 ( .A(B[24]), .B(A[24]), .Y(n147) );
  NAND2XL U193 ( .A(B[23]), .B(A[23]), .Y(n134) );
  OR2X4 U194 ( .A(A[28]), .B(B[28]), .Y(n100) );
  NOR2BX1 U195 ( .AN(n197), .B(n33), .Y(SUM[0]) );
  NOR2XL U196 ( .A(A[0]), .B(B[0]), .Y(n33) );
  INVX1 U197 ( .A(n226), .Y(n218) );
  INVXL U198 ( .A(n225), .Y(n224) );
  XOR2X1 U199 ( .A(n234), .B(n235), .Y(n267) );
  NOR2BXL U200 ( .AN(n193), .B(n183), .Y(n202) );
  NOR2BX1 U201 ( .AN(n61), .B(n31), .Y(n63) );
  XOR2X2 U202 ( .A(n204), .B(n205), .Y(SUM[17]) );
  NAND2XL U203 ( .A(n243), .B(n249), .Y(n251) );
  XNOR2X4 U204 ( .A(n12), .B(n168), .Y(SUM[21]) );
  XOR2X1 U205 ( .A(n223), .B(n66), .Y(SUM[4]) );
  NAND2X1 U206 ( .A(n97), .B(n83), .Y(n109) );
  INVX1 U207 ( .A(n113), .Y(n112) );
  INVX1 U208 ( .A(n60), .Y(n56) );
  INVX1 U209 ( .A(n103), .Y(n89) );
  NOR2BX1 U210 ( .AN(n213), .B(n40), .Y(n230) );
  NOR2X2 U211 ( .A(n182), .B(n193), .Y(n192) );
  INVX1 U212 ( .A(n102), .Y(n101) );
  NAND2X1 U213 ( .A(n61), .B(n65), .Y(n260) );
  INVX4 U214 ( .A(n245), .Y(n47) );
  NAND2XL U215 ( .A(n135), .B(n136), .Y(n133) );
  INVX1 U216 ( .A(n213), .Y(n212) );
  XOR2X1 U217 ( .A(n67), .B(n68), .Y(SUM[3]) );
  OAI21XL U218 ( .A0(n71), .A1(n72), .B0(n73), .Y(n67) );
  NOR2BX1 U219 ( .AN(n69), .B(n70), .Y(n68) );
  INVX1 U220 ( .A(n74), .Y(n71) );
  XOR2X1 U221 ( .A(n74), .B(n104), .Y(SUM[2]) );
  NOR2BX1 U222 ( .AN(n73), .B(n72), .Y(n104) );
  INVX1 U223 ( .A(n105), .Y(n72) );
  NOR2X2 U224 ( .A(n116), .B(n117), .Y(n115) );
  INVX1 U225 ( .A(n106), .Y(n196) );
  OAI2BB1X1 U226 ( .A0N(B[28]), .A1N(A[28]), .B0(n83), .Y(n80) );
  NOR2X1 U227 ( .A(n82), .B(n41), .Y(n81) );
  INVXL U228 ( .A(n91), .Y(n87) );
  NAND2XL U229 ( .A(B[28]), .B(A[28]), .Y(n113) );
  NAND2XL U230 ( .A(A[28]), .B(B[28]), .Y(n96) );
  XOR2X1 U231 ( .A(n107), .B(n195), .Y(SUM[1]) );
  INVX1 U232 ( .A(n197), .Y(n107) );
  NAND2X4 U233 ( .A(n208), .B(n209), .Y(n188) );
  NAND2X2 U234 ( .A(n159), .B(n136), .Y(n137) );
  NAND2X4 U235 ( .A(n138), .B(n170), .Y(n166) );
  NOR2BX4 U236 ( .AN(n28), .B(n145), .Y(n155) );
  OR2X2 U237 ( .A(A[9]), .B(B[9]), .Y(n245) );
  NAND2X1 U238 ( .A(B[18]), .B(A[18]), .Y(n193) );
  NAND2X2 U239 ( .A(B[11]), .B(A[11]), .Y(n249) );
  NAND2XL U240 ( .A(B[19]), .B(A[19]), .Y(n181) );
  NOR2X1 U241 ( .A(B[27]), .B(A[27]), .Y(n127) );
  NAND2XL U242 ( .A(B[21]), .B(A[21]), .Y(n167) );
  NAND2XL U243 ( .A(n181), .B(n187), .Y(n198) );
  NAND3X2 U244 ( .A(A[24]), .B(B[24]), .C(n118), .Y(n132) );
  INVX4 U245 ( .A(n238), .Y(n237) );
  INVX4 U246 ( .A(n232), .Y(n231) );
  INVX4 U247 ( .A(n186), .Y(n183) );
  CLKINVX3 U248 ( .A(n97), .Y(n82) );
  XOR2X4 U249 ( .A(n109), .B(n110), .Y(SUM[29]) );
  AOI21X4 U250 ( .A0(n111), .A1(n100), .B0(n112), .Y(n110) );
  OR2X4 U251 ( .A(A[29]), .B(B[29]), .Y(n97) );
  XOR2X4 U252 ( .A(n111), .B(n114), .Y(SUM[28]) );
  OAI2BB1X4 U253 ( .A0N(n121), .A1N(n118), .B0(n122), .Y(n91) );
  XOR2X4 U254 ( .A(n125), .B(n126), .Y(SUM[27]) );
  OAI21X4 U255 ( .A0(n128), .A1(n116), .B0(n124), .Y(n125) );
  AOI21X4 U256 ( .A0(n130), .A1(n129), .B0(n131), .Y(n128) );
  NAND2BX4 U257 ( .AN(n144), .B(n132), .Y(n131) );
  NOR2X4 U258 ( .A(n139), .B(n140), .Y(n129) );
  XOR2X4 U259 ( .A(n141), .B(n142), .Y(SUM[26]) );
  AOI21X4 U260 ( .A0(n143), .A1(n118), .B0(n144), .Y(n142) );
  OAI21X4 U261 ( .A0(n145), .A1(n146), .B0(n28), .Y(n143) );
  NAND2X4 U262 ( .A(n150), .B(n30), .Y(n149) );
  NOR2BX4 U263 ( .AN(n123), .B(n153), .Y(n152) );
  OR2X4 U264 ( .A(A[25]), .B(B[25]), .Y(n118) );
  NAND3BX4 U265 ( .AN(n148), .B(n30), .C(n11), .Y(n120) );
  NAND3X4 U266 ( .A(n136), .B(n156), .C(n135), .Y(n150) );
  NAND2X4 U267 ( .A(n157), .B(n158), .Y(n135) );
  NOR3BX4 U268 ( .AN(n156), .B(n138), .C(n137), .Y(n148) );
  XOR2X4 U269 ( .A(n162), .B(n163), .Y(SUM[23]) );
  OR2X4 U270 ( .A(A[23]), .B(B[23]), .Y(n156) );
  XOR2X4 U271 ( .A(n21), .B(n165), .Y(SUM[22]) );
  OR2X4 U272 ( .A(A[22]), .B(B[22]), .Y(n136) );
  NAND2X4 U273 ( .A(B[22]), .B(A[22]), .Y(n161) );
  NOR2BX4 U274 ( .AN(n167), .B(n169), .Y(n168) );
  OR2X4 U275 ( .A(B[21]), .B(A[21]), .Y(n159) );
  NAND2X4 U276 ( .A(n18), .B(n172), .Y(n138) );
  OR2X4 U277 ( .A(A[20]), .B(B[20]), .Y(n172) );
  AOI21X4 U278 ( .A0(n178), .A1(n179), .B0(n180), .Y(n177) );
  NOR2X4 U279 ( .A(n182), .B(n183), .Y(n179) );
  AOI21X4 U280 ( .A0(n191), .A1(n186), .B0(n192), .Y(n175) );
  NOR2X4 U281 ( .A(n182), .B(n194), .Y(n191) );
  XOR2X4 U282 ( .A(n199), .B(n198), .Y(SUM[19]) );
  OR2X4 U283 ( .A(B[19]), .B(A[19]), .Y(n187) );
  OR2X4 U284 ( .A(A[18]), .B(B[18]), .Y(n186) );
  NAND2X4 U285 ( .A(n206), .B(n185), .Y(n204) );
  OR2X4 U286 ( .A(A[16]), .B(B[16]), .Y(n189) );
  XOR2X4 U287 ( .A(n229), .B(n230), .Y(SUM[15]) );
  XOR2X4 U288 ( .A(n232), .B(n233), .Y(SUM[14]) );
  OAI21X4 U289 ( .A0(n237), .A1(n236), .B0(n214), .Y(n234) );
  OAI21X4 U290 ( .A0(n240), .A1(n217), .B0(n222), .Y(n238) );
  OAI2BB1X4 U291 ( .A0N(n241), .A1N(n242), .B0(n243), .Y(n222) );
  CLKINVX3 U292 ( .A(n249), .Y(n248) );
  OR2X4 U293 ( .A(B[11]), .B(A[11]), .Y(n243) );
  XOR2X4 U294 ( .A(n253), .B(n255), .Y(SUM[10]) );
  OR2X4 U295 ( .A(A[10]), .B(B[10]), .Y(n244) );
  OAI21X4 U296 ( .A0(n256), .A1(n47), .B0(n8), .Y(n253) );
  CLKINVX3 U297 ( .A(n45), .Y(n256) );
  NAND2X4 U298 ( .A(n257), .B(n50), .Y(n45) );
  NAND2BX4 U299 ( .AN(n55), .B(n258), .Y(n225) );
endmodule


module hash_core_DW01_add_30 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n240, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239;

  NAND3X2 U2 ( .A(n147), .B(n148), .C(n149), .Y(n146) );
  CLKINVX3 U3 ( .A(n141), .Y(n140) );
  AOI21X2 U4 ( .A0(n214), .A1(n215), .B0(n216), .Y(n212) );
  XOR2X4 U5 ( .A(n56), .B(n57), .Y(SUM[6]) );
  BUFX3 U6 ( .A(n27), .Y(n1) );
  NOR2X2 U7 ( .A(A[17]), .B(B[17]), .Y(n26) );
  XOR2X2 U8 ( .A(n107), .B(n108), .Y(SUM[27]) );
  NOR2X2 U9 ( .A(n22), .B(n1), .Y(n194) );
  OAI21X4 U10 ( .A0(n22), .A1(n181), .B0(n182), .Y(n179) );
  NOR2X2 U11 ( .A(A[13]), .B(B[13]), .Y(n22) );
  OAI21X4 U12 ( .A0(n1), .A1(n206), .B0(n181), .Y(n204) );
  INVX4 U13 ( .A(n207), .Y(n206) );
  BUFX4 U14 ( .A(n34), .Y(n2) );
  AOI2BB1XL U15 ( .A0N(n50), .A1N(n51), .B0(n52), .Y(n49) );
  NOR2X2 U16 ( .A(n23), .B(n50), .Y(n239) );
  NOR2X2 U17 ( .A(n23), .B(n50), .Y(n232) );
  NOR2BX1 U18 ( .AN(n53), .B(n50), .Y(n57) );
  INVX4 U19 ( .A(n55), .Y(n50) );
  AOI21X2 U20 ( .A0(n51), .A1(n60), .B0(n58), .Y(n231) );
  OAI21X1 U21 ( .A0(n62), .A1(n58), .B0(n51), .Y(n56) );
  INVX4 U22 ( .A(n54), .Y(n58) );
  NAND2X4 U23 ( .A(B[1]), .B(A[1]), .Y(n85) );
  OR2X4 U24 ( .A(A[1]), .B(B[1]), .Y(n83) );
  OAI21X4 U25 ( .A0(n203), .A1(n22), .B0(n182), .Y(n200) );
  INVX4 U26 ( .A(n204), .Y(n203) );
  AOI2BB1X2 U27 ( .A0N(n23), .A1N(n53), .B0(n234), .Y(n233) );
  INVXL U28 ( .A(n161), .Y(n15) );
  INVXL U29 ( .A(n26), .Y(n14) );
  XOR2X2 U30 ( .A(n200), .B(n202), .Y(SUM[14]) );
  NAND2X1 U31 ( .A(B[26]), .B(A[26]), .Y(n98) );
  NOR2BX1 U32 ( .AN(n98), .B(n99), .Y(n111) );
  OAI21X2 U33 ( .A0(n70), .A1(n25), .B0(n71), .Y(n66) );
  OR2X2 U34 ( .A(A[3]), .B(B[3]), .Y(n237) );
  INVX1 U35 ( .A(n201), .Y(n180) );
  NAND2X1 U36 ( .A(B[8]), .B(A[8]), .Y(n38) );
  INVX1 U37 ( .A(n174), .Y(n173) );
  AOI21X1 U38 ( .A0(n32), .A1(n219), .B0(n224), .Y(n226) );
  NAND2X1 U39 ( .A(n114), .B(n115), .Y(n93) );
  OR2X2 U40 ( .A(A[23]), .B(B[23]), .Y(n125) );
  OR2X2 U41 ( .A(A[22]), .B(B[22]), .Y(n131) );
  OAI2BB1X1 U42 ( .A0N(n209), .A1N(n41), .B0(n210), .Y(n207) );
  AOI21X1 U43 ( .A0(n211), .A1(n43), .B0(n189), .Y(n210) );
  OR2X2 U44 ( .A(A[4]), .B(B[4]), .Y(n59) );
  NAND2X1 U45 ( .A(B[5]), .B(A[5]), .Y(n51) );
  NAND2X1 U46 ( .A(B[3]), .B(A[3]), .Y(n68) );
  NOR2X1 U47 ( .A(A[11]), .B(B[11]), .Y(n24) );
  NAND2X1 U48 ( .A(B[10]), .B(A[10]), .Y(n217) );
  XOR2X2 U49 ( .A(n167), .B(n168), .Y(SUM[18]) );
  INVX1 U50 ( .A(n13), .Y(n167) );
  NOR2X2 U51 ( .A(A[7]), .B(B[7]), .Y(n23) );
  OR2X2 U52 ( .A(A[6]), .B(B[6]), .Y(n55) );
  OR2X2 U53 ( .A(A[5]), .B(B[5]), .Y(n54) );
  NAND2X1 U54 ( .A(n7), .B(n98), .Y(n107) );
  NAND2X1 U55 ( .A(n110), .B(n105), .Y(n7) );
  NAND2X2 U56 ( .A(n4), .B(n5), .Y(SUM[26]) );
  NAND2X1 U57 ( .A(n109), .B(n111), .Y(n5) );
  NOR2BX2 U58 ( .AN(n164), .B(n20), .Y(SUM[0]) );
  INVX1 U59 ( .A(n110), .Y(n109) );
  INVX2 U60 ( .A(n83), .Y(n163) );
  OR2X2 U61 ( .A(n39), .B(n35), .Y(n18) );
  CLKINVX3 U62 ( .A(n219), .Y(n35) );
  XOR2X2 U63 ( .A(n135), .B(n136), .Y(SUM[23]) );
  OAI2BB1X2 U64 ( .A0N(n227), .A1N(n41), .B0(n228), .Y(n32) );
  OR2X4 U65 ( .A(A[8]), .B(B[8]), .Y(n229) );
  XOR2X4 U66 ( .A(n198), .B(n199), .Y(SUM[15]) );
  AOI21X2 U67 ( .A0(n178), .A1(n200), .B0(n180), .Y(n199) );
  INVX2 U68 ( .A(n122), .Y(n143) );
  NAND2X4 U69 ( .A(n145), .B(n146), .Y(n122) );
  NAND2X1 U70 ( .A(n110), .B(n3), .Y(n4) );
  INVX1 U71 ( .A(n111), .Y(n3) );
  OR2X4 U72 ( .A(n222), .B(n218), .Y(n6) );
  NAND2X4 U73 ( .A(n6), .B(n217), .Y(n220) );
  AOI21XL U74 ( .A0(n32), .A1(n219), .B0(n224), .Y(n222) );
  NAND2X2 U75 ( .A(n225), .B(n9), .Y(n10) );
  NAND2X1 U76 ( .A(n8), .B(n226), .Y(n11) );
  NAND2X4 U77 ( .A(n10), .B(n11), .Y(SUM[10]) );
  INVXL U78 ( .A(n225), .Y(n8) );
  INVX2 U79 ( .A(n226), .Y(n9) );
  NAND2XL U80 ( .A(n217), .B(n223), .Y(n225) );
  OAI21X4 U81 ( .A0(n30), .A1(n143), .B0(n133), .Y(n141) );
  BUFX4 U82 ( .A(n240), .Y(SUM[22]) );
  AOI21X4 U83 ( .A0(n41), .A1(n59), .B0(n63), .Y(n62) );
  XOR2X2 U84 ( .A(n32), .B(n33), .Y(SUM[9]) );
  XOR2X4 U85 ( .A(n220), .B(n221), .Y(SUM[11]) );
  AOI21X4 U86 ( .A0(n169), .A1(n14), .B0(n15), .Y(n13) );
  OAI21X4 U87 ( .A0(n28), .A1(n171), .B0(n160), .Y(n169) );
  NOR2X4 U88 ( .A(A[2]), .B(B[2]), .Y(n25) );
  NAND2X4 U89 ( .A(B[2]), .B(A[2]), .Y(n71) );
  XOR2X4 U90 ( .A(n66), .B(n67), .Y(SUM[3]) );
  NAND2XL U91 ( .A(B[13]), .B(A[13]), .Y(n182) );
  NAND2XL U92 ( .A(B[4]), .B(A[4]), .Y(n60) );
  NAND2BX4 U93 ( .AN(n71), .B(n237), .Y(n238) );
  NOR2BX2 U94 ( .AN(n85), .B(n163), .Y(n162) );
  XNOR2X1 U95 ( .A(n76), .B(n19), .Y(SUM[30]) );
  INVX2 U96 ( .A(n158), .Y(n150) );
  NOR2XL U97 ( .A(A[20]), .B(B[20]), .Y(n30) );
  NAND2XL U98 ( .A(B[21]), .B(A[21]), .Y(n134) );
  NAND2XL U99 ( .A(B[17]), .B(A[17]), .Y(n161) );
  INVXL U100 ( .A(n184), .Y(n211) );
  NOR2XL U101 ( .A(n192), .B(n193), .Y(n190) );
  NAND2XL U102 ( .A(n190), .B(n191), .Y(n188) );
  NAND2XL U103 ( .A(n54), .B(n51), .Y(n61) );
  OAI21X2 U104 ( .A0(n140), .A1(n29), .B0(n134), .Y(n137) );
  OR2X4 U105 ( .A(n58), .B(n65), .Y(n16) );
  AOI21X1 U106 ( .A0(n178), .A1(n179), .B0(n180), .Y(n175) );
  XOR2X1 U107 ( .A(n207), .B(n208), .Y(SUM[12]) );
  OR2X4 U108 ( .A(n218), .B(n24), .Y(n17) );
  INVX2 U109 ( .A(n223), .Y(n218) );
  NAND2XL U110 ( .A(B[6]), .B(A[6]), .Y(n53) );
  NAND2XL U111 ( .A(B[9]), .B(A[9]), .Y(n34) );
  NAND2X1 U112 ( .A(B[24]), .B(A[24]), .Y(n102) );
  NOR2X1 U113 ( .A(A[21]), .B(B[21]), .Y(n29) );
  OAI21X4 U114 ( .A0(n183), .A1(n21), .B0(n173), .Y(n149) );
  INVXL U115 ( .A(n43), .Y(n42) );
  OAI2BB1X2 U116 ( .A0N(n83), .A1N(n84), .B0(n85), .Y(n72) );
  NOR2BX2 U117 ( .AN(n60), .B(n65), .Y(n64) );
  NAND3BX4 U118 ( .AN(n193), .B(n68), .C(n191), .Y(n41) );
  NOR2BXL U119 ( .AN(n130), .B(n123), .Y(n139) );
  NAND2XL U120 ( .A(n128), .B(n125), .Y(n135) );
  INVXL U121 ( .A(n130), .Y(n138) );
  OAI21X2 U122 ( .A0(n212), .A1(n24), .B0(n213), .Y(n189) );
  NOR2BXL U123 ( .AN(n103), .B(n101), .Y(n113) );
  INVX2 U124 ( .A(n229), .Y(n39) );
  OAI2BB1X2 U125 ( .A0N(n106), .A1N(n112), .B0(n103), .Y(n110) );
  NAND2BX4 U126 ( .AN(n16), .B(n239), .Y(n44) );
  OR2X4 U127 ( .A(n17), .B(n18), .Y(n184) );
  NOR2BXL U128 ( .AN(n155), .B(n151), .Y(n166) );
  OAI21X1 U129 ( .A0(n13), .A1(n150), .B0(n157), .Y(n165) );
  NOR2BXL U130 ( .AN(n2), .B(n35), .Y(n33) );
  NOR2BX1 U131 ( .AN(n104), .B(n96), .Y(n95) );
  NAND2X1 U132 ( .A(n74), .B(n77), .Y(n19) );
  XOR2XL U133 ( .A(n86), .B(n79), .Y(SUM[29]) );
  NOR2XL U134 ( .A(n44), .B(n39), .Y(n227) );
  AOI21XL U135 ( .A0(n43), .A1(n229), .B0(n230), .Y(n228) );
  NAND2XL U136 ( .A(n76), .B(n77), .Y(n75) );
  NAND2X4 U137 ( .A(B[0]), .B(A[0]), .Y(n164) );
  NOR2XL U138 ( .A(A[0]), .B(B[0]), .Y(n20) );
  NAND2X2 U139 ( .A(B[12]), .B(A[12]), .Y(n181) );
  OR2X4 U140 ( .A(A[9]), .B(B[9]), .Y(n219) );
  NOR2XL U141 ( .A(A[12]), .B(B[12]), .Y(n27) );
  NAND2XL U142 ( .A(B[18]), .B(A[18]), .Y(n157) );
  NAND2XL U143 ( .A(B[15]), .B(A[15]), .Y(n177) );
  NAND2XL U144 ( .A(B[11]), .B(A[11]), .Y(n213) );
  NAND2XL U145 ( .A(B[7]), .B(A[7]), .Y(n47) );
  NOR2XL U146 ( .A(A[16]), .B(B[16]), .Y(n28) );
  NAND2XL U147 ( .A(B[19]), .B(A[19]), .Y(n155) );
  NAND2XL U148 ( .A(B[25]), .B(A[25]), .Y(n103) );
  AOI21X1 U149 ( .A0(n187), .A1(n188), .B0(n189), .Y(n185) );
  NOR2X1 U150 ( .A(n184), .B(n44), .Y(n187) );
  NOR2X1 U151 ( .A(n35), .B(n218), .Y(n214) );
  NOR2X1 U152 ( .A(n184), .B(n44), .Y(n209) );
  NAND2BX1 U153 ( .AN(n184), .B(n43), .Y(n186) );
  AND2X2 U154 ( .A(n185), .B(n186), .Y(n21) );
  NOR2X1 U155 ( .A(n150), .B(n151), .Y(n147) );
  XOR2X2 U156 ( .A(n204), .B(n205), .Y(SUM[13]) );
  NOR2BX1 U157 ( .AN(n182), .B(n22), .Y(n205) );
  NOR2BX1 U158 ( .AN(n213), .B(n24), .Y(n221) );
  INVX1 U159 ( .A(n217), .Y(n216) );
  NAND2X1 U160 ( .A(n2), .B(n38), .Y(n215) );
  NOR2BX1 U161 ( .AN(n157), .B(n150), .Y(n168) );
  NOR2BX1 U162 ( .AN(n68), .B(n69), .Y(n67) );
  INVX1 U163 ( .A(n72), .Y(n70) );
  XOR2X1 U164 ( .A(n137), .B(n139), .Y(n240) );
  INVX1 U165 ( .A(n38), .Y(n230) );
  NAND2X1 U166 ( .A(n177), .B(n197), .Y(n198) );
  NOR2BX1 U167 ( .AN(n201), .B(n196), .Y(n202) );
  AOI21X1 U168 ( .A0(n131), .A1(n137), .B0(n138), .Y(n136) );
  INVX1 U169 ( .A(n59), .Y(n65) );
  INVX1 U170 ( .A(n178), .Y(n196) );
  XOR2X2 U171 ( .A(n45), .B(n46), .Y(SUM[7]) );
  NOR2BX1 U172 ( .AN(n47), .B(n23), .Y(n46) );
  OAI21X2 U173 ( .A0(n62), .A1(n48), .B0(n49), .Y(n45) );
  NAND2X1 U174 ( .A(n54), .B(n55), .Y(n48) );
  XOR2X1 U175 ( .A(n41), .B(n64), .Y(SUM[4]) );
  XOR2X1 U176 ( .A(n169), .B(n170), .Y(SUM[17]) );
  NOR2BX1 U177 ( .AN(n161), .B(n26), .Y(n170) );
  XOR2X1 U178 ( .A(n165), .B(n166), .Y(SUM[19]) );
  NOR2BX1 U179 ( .AN(n181), .B(n1), .Y(n208) );
  XOR2X1 U180 ( .A(n84), .B(n162), .Y(SUM[1]) );
  XOR2X1 U181 ( .A(n36), .B(n37), .Y(SUM[8]) );
  NOR2BX1 U182 ( .AN(n38), .B(n39), .Y(n37) );
  OAI2BB1X1 U183 ( .A0N(n40), .A1N(n41), .B0(n42), .Y(n36) );
  INVX1 U184 ( .A(n44), .Y(n40) );
  XOR2X1 U185 ( .A(n72), .B(n82), .Y(SUM[2]) );
  NOR2BX1 U186 ( .AN(n71), .B(n25), .Y(n82) );
  XOR2X2 U187 ( .A(n61), .B(n62), .Y(SUM[5]) );
  INVX1 U188 ( .A(n60), .Y(n63) );
  OAI21XL U189 ( .A0(n175), .A1(n176), .B0(n177), .Y(n174) );
  AOI21X1 U190 ( .A0(n152), .A1(n153), .B0(n154), .Y(n145) );
  INVX1 U191 ( .A(n155), .Y(n154) );
  INVX1 U192 ( .A(n53), .Y(n52) );
  INVX1 U193 ( .A(n164), .Y(n84) );
  INVX1 U194 ( .A(n149), .Y(n171) );
  INVX1 U195 ( .A(n47), .Y(n234) );
  NAND2X1 U196 ( .A(n194), .B(n195), .Y(n183) );
  NOR2X1 U197 ( .A(n176), .B(n196), .Y(n195) );
  OAI21XL U198 ( .A0(n93), .A1(n94), .B0(n95), .Y(n87) );
  NAND3BX1 U199 ( .AN(n31), .B(n105), .C(n106), .Y(n94) );
  INVX1 U200 ( .A(n197), .Y(n176) );
  INVX1 U201 ( .A(n2), .Y(n224) );
  INVX1 U202 ( .A(n153), .Y(n151) );
  XOR2X1 U203 ( .A(n87), .B(n91), .Y(SUM[28]) );
  NOR2BX1 U204 ( .AN(n90), .B(n92), .Y(n91) );
  INVX1 U205 ( .A(n88), .Y(n92) );
  XOR2X1 U206 ( .A(n141), .B(n142), .Y(SUM[21]) );
  NOR2BX1 U207 ( .AN(n134), .B(n29), .Y(n142) );
  XOR2X1 U208 ( .A(n122), .B(n144), .Y(SUM[20]) );
  NOR2BX1 U209 ( .AN(n133), .B(n30), .Y(n144) );
  XOR2X1 U210 ( .A(n149), .B(n172), .Y(SUM[16]) );
  NOR2BX1 U211 ( .AN(n160), .B(n28), .Y(n172) );
  NOR2BX1 U212 ( .AN(n104), .B(n31), .Y(n108) );
  XOR2X1 U213 ( .A(n114), .B(n116), .Y(SUM[24]) );
  NOR2BX1 U214 ( .AN(n102), .B(n117), .Y(n116) );
  INVX1 U215 ( .A(n115), .Y(n117) );
  XOR2X1 U216 ( .A(n112), .B(n113), .Y(SUM[25]) );
  NAND2X1 U217 ( .A(n118), .B(n119), .Y(n114) );
  AOI21X1 U218 ( .A0(n126), .A1(n125), .B0(n127), .Y(n118) );
  NAND3X1 U219 ( .A(n120), .B(n121), .C(n122), .Y(n119) );
  INVX1 U220 ( .A(n128), .Y(n127) );
  NOR2X1 U221 ( .A(n26), .B(n28), .Y(n148) );
  NAND2X1 U222 ( .A(n93), .B(n102), .Y(n112) );
  NAND2X1 U223 ( .A(n156), .B(n157), .Y(n152) );
  NAND2X1 U224 ( .A(n158), .B(n159), .Y(n156) );
  OAI21XL U225 ( .A0(n26), .A1(n160), .B0(n161), .Y(n159) );
  INVX1 U226 ( .A(n68), .Y(n192) );
  AOI21X1 U227 ( .A0(n87), .A1(n88), .B0(n89), .Y(n79) );
  INVX1 U228 ( .A(n90), .Y(n89) );
  OAI21XL U229 ( .A0(n78), .A1(n79), .B0(n80), .Y(n76) );
  INVX1 U230 ( .A(n81), .Y(n78) );
  INVX1 U231 ( .A(n131), .Y(n123) );
  NAND2X1 U232 ( .A(n129), .B(n130), .Y(n126) );
  NAND2X1 U233 ( .A(n131), .B(n132), .Y(n129) );
  OAI21XL U234 ( .A0(n29), .A1(n133), .B0(n134), .Y(n132) );
  NAND2X1 U235 ( .A(n80), .B(n81), .Y(n86) );
  NOR2X1 U236 ( .A(n29), .B(n30), .Y(n121) );
  NOR2X1 U237 ( .A(n123), .B(n124), .Y(n120) );
  INVX1 U238 ( .A(n125), .Y(n124) );
  NAND2X1 U239 ( .A(n74), .B(n75), .Y(n73) );
  INVX1 U240 ( .A(n105), .Y(n99) );
  INVX1 U241 ( .A(n106), .Y(n101) );
  AOI21X1 U242 ( .A0(n97), .A1(n98), .B0(n31), .Y(n96) );
  NAND2BX1 U243 ( .AN(n99), .B(n100), .Y(n97) );
  OAI21XL U244 ( .A0(n101), .A1(n102), .B0(n103), .Y(n100) );
  XOR3X2 U245 ( .A(B[31]), .B(A[31]), .C(n73), .Y(SUM[31]) );
  OR2X2 U246 ( .A(A[14]), .B(B[14]), .Y(n178) );
  NAND2X1 U247 ( .A(B[14]), .B(A[14]), .Y(n201) );
  OR2X2 U248 ( .A(A[10]), .B(B[10]), .Y(n223) );
  NAND2X1 U249 ( .A(B[16]), .B(A[16]), .Y(n160) );
  OR2X2 U250 ( .A(A[19]), .B(B[19]), .Y(n153) );
  OR2X2 U251 ( .A(A[18]), .B(B[18]), .Y(n158) );
  OR2X2 U252 ( .A(A[15]), .B(B[15]), .Y(n197) );
  NAND2X1 U253 ( .A(B[20]), .B(A[20]), .Y(n133) );
  NAND2X1 U254 ( .A(B[22]), .B(A[22]), .Y(n130) );
  NAND2X1 U255 ( .A(B[23]), .B(A[23]), .Y(n128) );
  OR2X2 U256 ( .A(A[24]), .B(B[24]), .Y(n115) );
  NOR2X1 U257 ( .A(A[27]), .B(B[27]), .Y(n31) );
  OR2X2 U258 ( .A(A[25]), .B(B[25]), .Y(n106) );
  NAND2X1 U259 ( .A(B[27]), .B(A[27]), .Y(n104) );
  OR2X2 U260 ( .A(A[28]), .B(B[28]), .Y(n88) );
  OR2X2 U261 ( .A(A[26]), .B(B[26]), .Y(n105) );
  NAND2X1 U262 ( .A(B[29]), .B(A[29]), .Y(n80) );
  NAND2X1 U263 ( .A(B[28]), .B(A[28]), .Y(n90) );
  OR2X2 U264 ( .A(A[30]), .B(B[30]), .Y(n77) );
  OR2X2 U265 ( .A(A[29]), .B(B[29]), .Y(n81) );
  NAND2X1 U266 ( .A(B[30]), .B(A[30]), .Y(n74) );
  OAI2BB1X4 U267 ( .A0N(n231), .A1N(n232), .B0(n233), .Y(n43) );
  NAND2X4 U268 ( .A(n235), .B(n236), .Y(n191) );
  NOR2X4 U269 ( .A(n69), .B(n25), .Y(n236) );
  CLKINVX3 U270 ( .A(n237), .Y(n69) );
  AOI21X4 U271 ( .A0(n85), .A1(n164), .B0(n163), .Y(n235) );
  CLKINVX3 U272 ( .A(n238), .Y(n193) );
endmodule


module hash_core_DW01_add_32 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n275, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n22, n23, n24, n25, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274;

  NOR3X4 U2 ( .A(n193), .B(n194), .C(n195), .Y(n192) );
  INVX1 U3 ( .A(n88), .Y(n176) );
  NAND2X4 U4 ( .A(B[16]), .B(A[16]), .Y(n170) );
  OAI21X4 U5 ( .A0(n258), .A1(n259), .B0(n260), .Y(n257) );
  NOR2BXL U6 ( .AN(n210), .B(n221), .Y(n242) );
  AOI21X1 U7 ( .A0(n114), .A1(n126), .B0(n127), .Y(n125) );
  NAND2X1 U8 ( .A(B[12]), .B(A[12]), .Y(n210) );
  NAND2X4 U9 ( .A(n79), .B(n60), .Y(n77) );
  AND3X4 U10 ( .A(n54), .B(n55), .C(n56), .Y(n33) );
  OAI21X4 U11 ( .A0(n265), .A1(n261), .B0(n262), .Y(n263) );
  NAND2X4 U12 ( .A(n1), .B(n2), .Y(n3) );
  NAND2X4 U13 ( .A(n3), .B(n75), .Y(n70) );
  INVX4 U14 ( .A(n74), .Y(n1) );
  INVX4 U15 ( .A(n9), .Y(n2) );
  INVX3 U16 ( .A(n198), .Y(n74) );
  OAI2BB1X2 U17 ( .A0N(n45), .A1N(n34), .B0(n262), .Y(n258) );
  AOI21X4 U18 ( .A0(n199), .A1(n200), .B0(n201), .Y(n189) );
  NOR2X2 U19 ( .A(n195), .B(n194), .Y(n199) );
  NOR2BX4 U20 ( .AN(n76), .B(n83), .Y(n82) );
  NOR2BX1 U21 ( .AN(n76), .B(n197), .Y(n196) );
  NAND2X2 U22 ( .A(B[3]), .B(A[3]), .Y(n76) );
  NOR2X1 U23 ( .A(A[0]), .B(B[0]), .Y(n101) );
  NOR2X2 U24 ( .A(n209), .B(n221), .Y(n217) );
  NAND2BX4 U25 ( .AN(n221), .B(n216), .Y(n233) );
  CLKINVX3 U26 ( .A(n239), .Y(n221) );
  NAND2X4 U27 ( .A(B[2]), .B(A[2]), .Y(n86) );
  NAND2BX4 U28 ( .AN(n243), .B(n240), .Y(n215) );
  INVX4 U29 ( .A(n238), .Y(n243) );
  BUFX8 U30 ( .A(n63), .Y(n4) );
  BUFX8 U31 ( .A(n65), .Y(n5) );
  OAI21X4 U32 ( .A0(n80), .A1(n193), .B0(n254), .Y(n10) );
  NAND2X2 U33 ( .A(n213), .B(n214), .Y(n188) );
  CLKINVX8 U34 ( .A(n193), .Y(n50) );
  NOR3BX4 U35 ( .AN(n38), .B(n261), .C(n193), .Y(n259) );
  NAND2X1 U36 ( .A(n61), .B(n62), .Y(n57) );
  OR2X4 U37 ( .A(A[6]), .B(B[6]), .Y(n62) );
  INVX4 U38 ( .A(n261), .Y(n34) );
  NAND2X4 U39 ( .A(n253), .B(n46), .Y(n261) );
  CLKINVX2 U40 ( .A(n45), .Y(n254) );
  NAND2X4 U41 ( .A(n212), .B(n53), .Y(n45) );
  OAI2BB1X4 U42 ( .A0N(n244), .A1N(n245), .B0(n246), .Y(n240) );
  NOR2X2 U43 ( .A(n42), .B(n250), .Y(n244) );
  NOR2BX4 U44 ( .AN(n7), .B(n248), .Y(n246) );
  BUFX4 U45 ( .A(n41), .Y(n6) );
  BUFX4 U46 ( .A(n247), .Y(n7) );
  CLKINVX8 U47 ( .A(n61), .Y(n72) );
  OR2X4 U48 ( .A(A[5]), .B(B[5]), .Y(n61) );
  INVX2 U49 ( .A(n208), .Y(n207) );
  INVX1 U50 ( .A(n194), .Y(n214) );
  OR2X2 U51 ( .A(A[21]), .B(B[21]), .Y(n149) );
  NAND3BXL U52 ( .AN(n36), .B(n173), .C(n174), .Y(n162) );
  NAND2X1 U53 ( .A(B[20]), .B(A[20]), .Y(n145) );
  OR2X2 U54 ( .A(A[25]), .B(B[25]), .Y(n112) );
  NAND3BX2 U55 ( .AN(n57), .B(n58), .C(n38), .Y(n56) );
  INVX1 U56 ( .A(n249), .Y(n248) );
  OAI21XL U57 ( .A0(n169), .A1(n170), .B0(n171), .Y(n168) );
  INVX1 U58 ( .A(n172), .Y(n163) );
  OAI21XL U59 ( .A0(n144), .A1(n145), .B0(n146), .Y(n143) );
  NAND2X1 U60 ( .A(n6), .B(n48), .Y(n245) );
  OR2X2 U61 ( .A(A[12]), .B(B[12]), .Y(n239) );
  INVX1 U62 ( .A(n103), .Y(n12) );
  INVX1 U63 ( .A(n148), .Y(n142) );
  NOR2X1 U64 ( .A(A[23]), .B(B[23]), .Y(n37) );
  NOR2BX1 U65 ( .AN(n141), .B(n142), .Y(n153) );
  OR2X2 U66 ( .A(A[24]), .B(B[24]), .Y(n132) );
  NOR2X2 U67 ( .A(n20), .B(n89), .Y(n84) );
  NAND2X1 U68 ( .A(n204), .B(n220), .Y(n222) );
  AOI21X2 U69 ( .A0(n224), .A1(n11), .B0(n226), .Y(n223) );
  OAI21XL U70 ( .A0(n219), .A1(n211), .B0(n208), .Y(n226) );
  INVX1 U71 ( .A(n211), .Y(n230) );
  OR2X2 U72 ( .A(A[11]), .B(B[11]), .Y(n238) );
  INVX1 U73 ( .A(n48), .Y(n47) );
  OAI2BB1X1 U74 ( .A0N(n6), .A1N(n48), .B0(n253), .Y(n262) );
  XOR2X1 U75 ( .A(n157), .B(n159), .Y(SUM[20]) );
  XOR2X2 U76 ( .A(n182), .B(n183), .Y(SUM[17]) );
  XOR2X2 U77 ( .A(n180), .B(n181), .Y(SUM[18]) );
  XOR2X2 U78 ( .A(n177), .B(n178), .Y(SUM[19]) );
  INVX1 U79 ( .A(n180), .Y(n179) );
  NOR2BX1 U80 ( .AN(n211), .B(n209), .Y(n231) );
  XOR2X1 U81 ( .A(n129), .B(n130), .Y(SUM[25]) );
  CLKINVX3 U82 ( .A(n175), .Y(n13) );
  NOR2BX4 U83 ( .AN(n90), .B(n176), .Y(n175) );
  OAI2BB1X2 U84 ( .A0N(B[0]), .A1N(A[0]), .B0(n90), .Y(n198) );
  INVX1 U85 ( .A(n90), .Y(n89) );
  NAND2X1 U86 ( .A(n100), .B(n90), .Y(n22) );
  AND3X4 U87 ( .A(n87), .B(n271), .C(n88), .Y(n8) );
  OAI21X4 U88 ( .A0(n232), .A1(n233), .B0(n234), .Y(n225) );
  OAI21X2 U89 ( .A0(n232), .A1(n233), .B0(n234), .Y(n11) );
  INVX4 U90 ( .A(n8), .Y(n9) );
  NAND2XL U91 ( .A(n212), .B(n53), .Y(n200) );
  OAI21X4 U92 ( .A0(n69), .A1(n70), .B0(n71), .Y(n68) );
  AOI21X2 U93 ( .A0(n50), .A1(n38), .B0(n45), .Y(n265) );
  OAI21X4 U94 ( .A0(n232), .A1(n195), .B0(n215), .Y(n241) );
  AOI21X2 U95 ( .A0(n229), .A1(n225), .B0(n230), .Y(n228) );
  CLKINVX4 U96 ( .A(n103), .Y(n102) );
  NAND2X2 U97 ( .A(A[1]), .B(B[1]), .Y(n90) );
  AOI2BB1X4 U98 ( .A0N(n235), .A1N(n236), .B0(n237), .Y(n234) );
  CLKINVX4 U99 ( .A(n240), .Y(n235) );
  NAND2X4 U100 ( .A(B[8]), .B(A[8]), .Y(n48) );
  INVX8 U101 ( .A(n229), .Y(n209) );
  NAND2X4 U102 ( .A(n111), .B(n122), .Y(n129) );
  NAND2X4 U103 ( .A(n131), .B(n132), .Y(n111) );
  XOR2X4 U104 ( .A(n155), .B(n156), .Y(SUM[21]) );
  NAND2X4 U105 ( .A(n135), .B(n145), .Y(n155) );
  INVX8 U106 ( .A(n38), .Y(n80) );
  BUFX16 U107 ( .A(n59), .Y(n38) );
  NOR2BX1 U108 ( .AN(n48), .B(n49), .Y(n51) );
  NAND2X2 U109 ( .A(n103), .B(n175), .Y(n14) );
  NAND2X4 U110 ( .A(n12), .B(n13), .Y(n15) );
  NAND2X4 U111 ( .A(n14), .B(n15), .Y(n275) );
  NAND2X4 U112 ( .A(B[0]), .B(A[0]), .Y(n103) );
  BUFX12 U113 ( .A(n275), .Y(SUM[1]) );
  NAND2X2 U114 ( .A(n152), .B(n17), .Y(n18) );
  NAND2X4 U115 ( .A(n16), .B(n153), .Y(n19) );
  NAND2X4 U116 ( .A(n18), .B(n19), .Y(SUM[22]) );
  INVX4 U117 ( .A(n152), .Y(n16) );
  INVX1 U118 ( .A(n153), .Y(n17) );
  AND2X2 U119 ( .A(n88), .B(n102), .Y(n20) );
  OAI21X4 U120 ( .A0(n84), .A1(n85), .B0(n86), .Y(n81) );
  NAND2X1 U121 ( .A(n58), .B(n38), .Y(n79) );
  AOI21X2 U122 ( .A0(n205), .A1(n206), .B0(n207), .Y(n202) );
  NAND3BXL U123 ( .AN(n101), .B(n102), .C(n88), .Y(n100) );
  NAND2X2 U124 ( .A(B[6]), .B(A[6]), .Y(n63) );
  OAI21X1 U125 ( .A0(n209), .A1(n210), .B0(n211), .Y(n206) );
  NAND2X2 U126 ( .A(B[13]), .B(A[13]), .Y(n211) );
  OAI21X4 U127 ( .A0(n135), .A1(n136), .B0(n137), .Y(n131) );
  XNOR2X2 U128 ( .A(n126), .B(n25), .Y(SUM[26]) );
  CLKINVX8 U129 ( .A(n31), .Y(n157) );
  XOR2XL U130 ( .A(n104), .B(n97), .Y(SUM[29]) );
  NAND2X2 U131 ( .A(B[5]), .B(A[5]), .Y(n65) );
  NOR2BXL U132 ( .AN(n172), .B(n36), .Y(n178) );
  NAND2XL U133 ( .A(B[19]), .B(A[19]), .Y(n172) );
  OR2XL U134 ( .A(A[20]), .B(B[20]), .Y(n158) );
  NOR2BXL U135 ( .AN(n146), .B(n144), .Y(n156) );
  AOI2BB1X4 U136 ( .A0N(n161), .A1N(n162), .B0(n32), .Y(n31) );
  NAND3BXL U137 ( .AN(n37), .B(n148), .C(n149), .Y(n136) );
  NAND2X1 U138 ( .A(n119), .B(n114), .Y(n25) );
  NOR2X1 U139 ( .A(A[19]), .B(B[19]), .Y(n36) );
  NAND2XL U140 ( .A(B[18]), .B(A[18]), .Y(n166) );
  NAND2X1 U141 ( .A(B[17]), .B(A[17]), .Y(n171) );
  NAND2X1 U142 ( .A(B[21]), .B(A[21]), .Y(n146) );
  NAND2X1 U143 ( .A(B[25]), .B(A[25]), .Y(n123) );
  NAND2X1 U144 ( .A(B[24]), .B(A[24]), .Y(n122) );
  NOR2X4 U145 ( .A(n72), .B(n73), .Y(n273) );
  NOR2X4 U146 ( .A(n269), .B(n66), .Y(n274) );
  NAND2X2 U147 ( .A(n191), .B(n192), .Y(n190) );
  XOR2X4 U148 ( .A(n22), .B(n23), .Y(SUM[2]) );
  AND2X1 U149 ( .A(n87), .B(n86), .Y(n23) );
  XOR2X4 U150 ( .A(n80), .B(n24), .Y(SUM[4]) );
  NAND2XL U151 ( .A(n60), .B(n58), .Y(n24) );
  INVXL U152 ( .A(n119), .Y(n127) );
  OR2X4 U153 ( .A(n163), .B(n164), .Y(n32) );
  NAND2X2 U154 ( .A(n128), .B(n123), .Y(n126) );
  NAND2X2 U155 ( .A(n112), .B(n129), .Y(n128) );
  NAND2X4 U156 ( .A(n157), .B(n158), .Y(n135) );
  XNOR2X4 U157 ( .A(n77), .B(n78), .Y(SUM[5]) );
  XOR2X2 U158 ( .A(n94), .B(n35), .Y(SUM[30]) );
  XNOR2X1 U159 ( .A(n105), .B(n27), .Y(SUM[28]) );
  NAND2X1 U160 ( .A(n108), .B(n106), .Y(n27) );
  NOR2BXL U161 ( .AN(n171), .B(n169), .Y(n183) );
  NOR2BXL U162 ( .AN(n166), .B(n167), .Y(n181) );
  XNOR2X4 U163 ( .A(n33), .B(n28), .Y(SUM[7]) );
  AND2X1 U164 ( .A(n52), .B(n53), .Y(n28) );
  AOI21XL U165 ( .A0(n45), .A1(n46), .B0(n47), .Y(n44) );
  AND2X1 U166 ( .A(n249), .B(n238), .Y(n29) );
  AND2X1 U167 ( .A(n4), .B(n62), .Y(n30) );
  OAI21X4 U168 ( .A0(n16), .A1(n142), .B0(n141), .Y(n150) );
  NAND2XL U169 ( .A(n94), .B(n95), .Y(n93) );
  INVXL U170 ( .A(n7), .Y(n256) );
  OR2X4 U171 ( .A(A[17]), .B(B[17]), .Y(n174) );
  OR2X4 U172 ( .A(A[18]), .B(B[18]), .Y(n173) );
  NAND2XL U173 ( .A(B[22]), .B(A[22]), .Y(n141) );
  OR2XL U174 ( .A(A[16]), .B(B[16]), .Y(n185) );
  NAND2XL U175 ( .A(B[23]), .B(A[23]), .Y(n147) );
  INVXL U176 ( .A(n195), .Y(n216) );
  NOR2XL U177 ( .A(n209), .B(n219), .Y(n224) );
  NAND2XL U178 ( .A(n208), .B(n205), .Y(n227) );
  OAI21XL U179 ( .A0(n9), .A1(n74), .B0(n196), .Y(n191) );
  NOR2X1 U180 ( .A(n138), .B(n139), .Y(n137) );
  INVX1 U181 ( .A(n147), .Y(n138) );
  INVX1 U182 ( .A(n173), .Y(n167) );
  INVX1 U183 ( .A(n174), .Y(n169) );
  NOR2BXL U184 ( .AN(n6), .B(n42), .Y(n40) );
  NOR2BX1 U185 ( .AN(n145), .B(n160), .Y(n159) );
  INVX1 U186 ( .A(n158), .Y(n160) );
  XOR2X1 U187 ( .A(n184), .B(n186), .Y(SUM[16]) );
  NOR2BX1 U188 ( .AN(n170), .B(n187), .Y(n186) );
  INVX1 U189 ( .A(n185), .Y(n187) );
  NOR2BX1 U190 ( .AN(n147), .B(n37), .Y(n151) );
  NOR2BXL U191 ( .AN(n7), .B(n250), .Y(n264) );
  NOR2BX1 U192 ( .AN(n123), .B(n121), .Y(n130) );
  XOR2X1 U193 ( .A(n124), .B(n125), .Y(SUM[27]) );
  NAND2X1 U194 ( .A(n117), .B(n113), .Y(n124) );
  NAND2XL U195 ( .A(n60), .B(n76), .Y(n69) );
  AOI21X1 U196 ( .A0(n165), .A1(n166), .B0(n36), .Y(n164) );
  NAND2BX1 U197 ( .AN(n167), .B(n168), .Y(n165) );
  INVXL U198 ( .A(n271), .Y(n83) );
  NOR2BX1 U199 ( .AN(n4), .B(n64), .Y(n54) );
  NOR2XL U200 ( .A(n5), .B(n66), .Y(n64) );
  INVXL U201 ( .A(n87), .Y(n85) );
  INVX1 U202 ( .A(n210), .Y(n237) );
  OR2XL U203 ( .A(n57), .B(n60), .Y(n55) );
  NAND2XL U204 ( .A(n61), .B(n5), .Y(n78) );
  NAND2XL U205 ( .A(n238), .B(n239), .Y(n236) );
  AOI21X1 U206 ( .A0(n105), .A1(n106), .B0(n107), .Y(n97) );
  INVX1 U207 ( .A(n108), .Y(n107) );
  OAI21XL U208 ( .A0(n96), .A1(n97), .B0(n98), .Y(n94) );
  INVX1 U209 ( .A(n99), .Y(n96) );
  INVX1 U210 ( .A(n149), .Y(n144) );
  XOR2X1 U211 ( .A(n131), .B(n133), .Y(SUM[24]) );
  NOR2BX1 U212 ( .AN(n122), .B(n134), .Y(n133) );
  INVX1 U213 ( .A(n132), .Y(n134) );
  NAND2X1 U214 ( .A(n98), .B(n99), .Y(n104) );
  NAND2X1 U215 ( .A(n109), .B(n110), .Y(n105) );
  AOI21X1 U216 ( .A0(n115), .A1(n113), .B0(n116), .Y(n109) );
  NAND4BXL U217 ( .AN(n111), .B(n112), .C(n113), .D(n114), .Y(n110) );
  INVX1 U218 ( .A(n117), .Y(n116) );
  AOI21X1 U219 ( .A0(n140), .A1(n141), .B0(n37), .Y(n139) );
  NAND2BX1 U220 ( .AN(n142), .B(n143), .Y(n140) );
  AND2X2 U221 ( .A(n92), .B(n95), .Y(n35) );
  INVX1 U222 ( .A(n112), .Y(n121) );
  NAND2X1 U223 ( .A(n92), .B(n93), .Y(n91) );
  NAND2X1 U224 ( .A(n118), .B(n119), .Y(n115) );
  NAND2X1 U225 ( .A(n114), .B(n120), .Y(n118) );
  OAI21XL U226 ( .A0(n121), .A1(n122), .B0(n123), .Y(n120) );
  AND2X2 U227 ( .A(n103), .B(n272), .Y(SUM[0]) );
  OR2XL U228 ( .A(A[0]), .B(B[0]), .Y(n272) );
  NAND2XL U229 ( .A(B[7]), .B(A[7]), .Y(n53) );
  NAND2XL U230 ( .A(B[14]), .B(A[14]), .Y(n208) );
  NAND2XL U231 ( .A(B[9]), .B(A[9]), .Y(n41) );
  NAND2XL U232 ( .A(B[10]), .B(A[10]), .Y(n247) );
  NAND2XL U233 ( .A(B[15]), .B(A[15]), .Y(n204) );
  NAND2XL U234 ( .A(B[11]), .B(A[11]), .Y(n249) );
  XOR3X2 U235 ( .A(B[31]), .B(A[31]), .C(n91), .Y(SUM[31]) );
  OR2X2 U236 ( .A(A[22]), .B(B[22]), .Y(n148) );
  OR2X2 U237 ( .A(A[26]), .B(B[26]), .Y(n114) );
  NAND2X1 U238 ( .A(B[26]), .B(A[26]), .Y(n119) );
  OR2X2 U239 ( .A(A[27]), .B(B[27]), .Y(n113) );
  NAND2X1 U240 ( .A(B[27]), .B(A[27]), .Y(n117) );
  NAND2X1 U241 ( .A(B[28]), .B(A[28]), .Y(n108) );
  OR2X2 U242 ( .A(A[28]), .B(B[28]), .Y(n106) );
  NAND2X1 U243 ( .A(B[30]), .B(A[30]), .Y(n92) );
  NAND2X1 U244 ( .A(B[29]), .B(A[29]), .Y(n98) );
  OR2X2 U245 ( .A(A[30]), .B(B[30]), .Y(n95) );
  OR2X2 U246 ( .A(A[29]), .B(B[29]), .Y(n99) );
  NAND3BX4 U247 ( .AN(n197), .B(n76), .C(n270), .Y(n59) );
  NAND3X4 U248 ( .A(n189), .B(n190), .C(n188), .Y(n184) );
  NOR2X1 U249 ( .A(n72), .B(n73), .Y(n71) );
  INVX8 U250 ( .A(n62), .Y(n66) );
  OAI21X2 U251 ( .A0(n80), .A1(n43), .B0(n44), .Y(n39) );
  NAND2X4 U252 ( .A(n8), .B(n198), .Y(n270) );
  INVX8 U253 ( .A(n10), .Y(n232) );
  XOR2X4 U254 ( .A(n10), .B(n51), .Y(SUM[8]) );
  XOR2X4 U255 ( .A(n39), .B(n40), .Y(SUM[9]) );
  NAND2BX4 U256 ( .AN(n49), .B(n50), .Y(n43) );
  XOR2X4 U257 ( .A(n67), .B(n30), .Y(SUM[6]) );
  NAND2X4 U258 ( .A(n68), .B(n5), .Y(n67) );
  XOR2X4 U259 ( .A(n81), .B(n82), .Y(SUM[3]) );
  XOR2X4 U260 ( .A(n150), .B(n151), .Y(SUM[23]) );
  NAND2X4 U261 ( .A(n154), .B(n146), .Y(n152) );
  NAND2X4 U262 ( .A(n149), .B(n155), .Y(n154) );
  OAI21X4 U263 ( .A0(n179), .A1(n167), .B0(n166), .Y(n177) );
  OAI2BB1X4 U264 ( .A0N(n174), .A1N(n182), .B0(n171), .Y(n180) );
  NAND2X4 U265 ( .A(n161), .B(n170), .Y(n182) );
  NAND2X4 U266 ( .A(n184), .B(n185), .Y(n161) );
  OAI21X4 U267 ( .A0(n202), .A1(n203), .B0(n204), .Y(n201) );
  CLKINVX3 U268 ( .A(n215), .Y(n213) );
  NAND2X4 U269 ( .A(n217), .B(n218), .Y(n194) );
  NOR2X4 U270 ( .A(n203), .B(n219), .Y(n218) );
  CLKINVX3 U271 ( .A(n220), .Y(n203) );
  XOR2X4 U272 ( .A(n222), .B(n223), .Y(SUM[15]) );
  CLKINVX3 U273 ( .A(n205), .Y(n219) );
  OR2X4 U274 ( .A(A[15]), .B(B[15]), .Y(n220) );
  XOR2X4 U275 ( .A(n228), .B(n227), .Y(SUM[14]) );
  OR2X4 U276 ( .A(A[14]), .B(B[14]), .Y(n205) );
  XOR2X4 U277 ( .A(n225), .B(n231), .Y(SUM[13]) );
  OR2X4 U278 ( .A(A[13]), .B(B[13]), .Y(n229) );
  XOR2X4 U279 ( .A(n241), .B(n242), .Y(SUM[12]) );
  NAND2X4 U280 ( .A(n251), .B(n252), .Y(n195) );
  NOR2X4 U281 ( .A(n49), .B(n42), .Y(n252) );
  CLKINVX3 U282 ( .A(n253), .Y(n42) );
  CLKINVX3 U283 ( .A(n46), .Y(n49) );
  NOR2X4 U284 ( .A(n250), .B(n243), .Y(n251) );
  XOR2X4 U285 ( .A(n255), .B(n29), .Y(SUM[11]) );
  NAND2BX4 U286 ( .AN(n256), .B(n257), .Y(n255) );
  XOR2X4 U287 ( .A(n263), .B(n264), .Y(SUM[10]) );
  CLKINVX3 U288 ( .A(n260), .Y(n250) );
  OR2X4 U289 ( .A(A[10]), .B(B[10]), .Y(n260) );
  OR2X4 U290 ( .A(A[8]), .B(B[8]), .Y(n46) );
  OR2X4 U291 ( .A(A[9]), .B(B[9]), .Y(n253) );
  NAND3X4 U292 ( .A(n266), .B(n267), .C(n268), .Y(n212) );
  NAND3X4 U293 ( .A(n5), .B(n4), .C(n60), .Y(n268) );
  NAND2X4 U294 ( .A(B[4]), .B(A[4]), .Y(n60) );
  NOR2X4 U295 ( .A(n269), .B(n66), .Y(n267) );
  NAND2X4 U296 ( .A(n72), .B(n4), .Y(n266) );
  OR2X4 U297 ( .A(A[1]), .B(B[1]), .Y(n88) );
  OR2X4 U298 ( .A(A[2]), .B(B[2]), .Y(n87) );
  CLKINVX3 U299 ( .A(n75), .Y(n197) );
  NAND2BX4 U300 ( .AN(n86), .B(n271), .Y(n75) );
  OR2X4 U301 ( .A(A[3]), .B(B[3]), .Y(n271) );
  NAND2X4 U302 ( .A(n273), .B(n274), .Y(n193) );
  CLKINVX3 U303 ( .A(n52), .Y(n269) );
  OR2X4 U304 ( .A(A[7]), .B(B[7]), .Y(n52) );
  CLKINVX3 U305 ( .A(n58), .Y(n73) );
  OR2X4 U306 ( .A(A[4]), .B(B[4]), .Y(n58) );
endmodule


module hash_core_DW01_add_38 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n274, n275, n276, n277, n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273;

  CLKINVX8 U2 ( .A(n161), .Y(n160) );
  NAND2X1 U3 ( .A(n45), .B(n70), .Y(n68) );
  INVX4 U4 ( .A(n93), .Y(n91) );
  XOR2X2 U5 ( .A(n93), .B(n104), .Y(n277) );
  INVX8 U6 ( .A(n186), .Y(n185) );
  NAND2X2 U7 ( .A(B[13]), .B(A[13]), .Y(n222) );
  INVX2 U8 ( .A(n164), .Y(n25) );
  NAND2X4 U9 ( .A(n111), .B(n112), .Y(n109) );
  AOI21X4 U10 ( .A0(n71), .A1(n49), .B0(n73), .Y(n67) );
  BUFX16 U11 ( .A(n72), .Y(n49) );
  NAND2X2 U12 ( .A(n223), .B(n222), .Y(n1) );
  NAND2X4 U13 ( .A(n2), .B(n224), .Y(n219) );
  INVX4 U14 ( .A(n1), .Y(n2) );
  AOI21X4 U15 ( .A0(n218), .A1(n219), .B0(n220), .Y(n195) );
  NAND2X2 U16 ( .A(n37), .B(n192), .Y(n5) );
  NAND2X4 U17 ( .A(n3), .B(n4), .Y(n6) );
  NAND2X4 U18 ( .A(n5), .B(n6), .Y(SUM[17]) );
  CLKINVX3 U19 ( .A(n37), .Y(n3) );
  INVX4 U20 ( .A(n192), .Y(n4) );
  NAND2X4 U21 ( .A(n169), .B(n170), .Y(n168) );
  NAND2X1 U22 ( .A(n71), .B(n270), .Y(n80) );
  OAI21X4 U23 ( .A0(n67), .A1(n68), .B0(n69), .Y(n65) );
  NAND2X4 U24 ( .A(B[0]), .B(A[0]), .Y(n182) );
  INVX3 U25 ( .A(n247), .Y(n246) );
  NOR2X1 U26 ( .A(A[20]), .B(B[20]), .Y(n44) );
  NAND2X4 U27 ( .A(B[20]), .B(A[20]), .Y(n152) );
  NOR2BX2 U28 ( .AN(n177), .B(n172), .Y(n194) );
  NAND2X2 U29 ( .A(B[16]), .B(A[16]), .Y(n177) );
  BUFX4 U30 ( .A(n274), .Y(SUM[24]) );
  OAI21X4 U31 ( .A0(n171), .A1(n177), .B0(n178), .Y(n176) );
  NOR4X4 U32 ( .A(n43), .B(n42), .C(n171), .D(n172), .Y(n170) );
  INVX4 U33 ( .A(n190), .Y(n171) );
  INVX2 U34 ( .A(n156), .Y(n151) );
  INVX2 U35 ( .A(n216), .Y(n261) );
  INVX1 U36 ( .A(n58), .Y(n259) );
  NAND3BX2 U37 ( .AN(n211), .B(n205), .C(n206), .Y(n207) );
  INVXL U38 ( .A(A[12]), .Y(n13) );
  NAND2X1 U39 ( .A(n36), .B(n28), .Y(n29) );
  NAND4BX2 U40 ( .AN(n14), .B(n64), .C(n249), .D(n250), .Y(n211) );
  OAI2BB1X2 U41 ( .A0N(n210), .A1N(n199), .B0(n62), .Y(n237) );
  AOI21X2 U42 ( .A0(n174), .A1(n175), .B0(n43), .Y(n173) );
  AOI21X2 U43 ( .A0(n58), .A1(n63), .B0(n14), .Y(n243) );
  NOR2BX2 U44 ( .AN(n230), .B(n225), .Y(n231) );
  OAI21X2 U45 ( .A0(n91), .A1(n46), .B0(n92), .Y(n87) );
  AOI2BB1X2 U46 ( .A0N(n51), .A1N(n52), .B0(n265), .Y(n66) );
  INVX1 U47 ( .A(n152), .Y(n28) );
  INVX4 U48 ( .A(n105), .Y(n181) );
  NAND2X1 U49 ( .A(B[21]), .B(A[21]), .Y(n153) );
  NOR2BX2 U50 ( .AN(n107), .B(n181), .Y(n180) );
  NAND2X1 U51 ( .A(n64), .B(n210), .Y(n266) );
  OR2X2 U52 ( .A(A[17]), .B(B[17]), .Y(n190) );
  OR2X2 U53 ( .A(A[16]), .B(B[16]), .Y(n191) );
  NAND2X1 U54 ( .A(B[19]), .B(A[19]), .Y(n179) );
  INVX1 U55 ( .A(n14), .Y(n251) );
  OAI2BB1X2 U56 ( .A0N(n12), .A1N(n165), .B0(n152), .Y(n163) );
  INVX1 U57 ( .A(n44), .Y(n12) );
  NOR2X1 U58 ( .A(n118), .B(n119), .Y(n117) );
  INVX1 U59 ( .A(n128), .Y(n118) );
  INVX1 U60 ( .A(n165), .Y(n144) );
  INVX4 U61 ( .A(n234), .Y(n232) );
  NOR2BX1 U62 ( .AN(n206), .B(n211), .Y(n236) );
  AOI21X2 U63 ( .A0(n201), .A1(n206), .B0(n239), .Y(n238) );
  NAND2BX2 U64 ( .AN(n54), .B(A[3]), .Y(n89) );
  CLKINVX3 U65 ( .A(n250), .Y(n248) );
  INVX1 U66 ( .A(n129), .Y(n123) );
  INVX1 U67 ( .A(n149), .Y(n20) );
  XNOR2X2 U68 ( .A(n38), .B(n33), .Y(SUM[12]) );
  NOR2X2 U69 ( .A(n241), .B(n201), .Y(n33) );
  INVX1 U70 ( .A(n270), .Y(n84) );
  BUFX3 U71 ( .A(n277), .Y(SUM[2]) );
  XOR2X1 U72 ( .A(n97), .B(n99), .Y(SUM[30]) );
  NAND2X4 U73 ( .A(n260), .B(n49), .Y(n62) );
  AOI21X4 U74 ( .A0(n209), .A1(n228), .B0(n229), .Y(n227) );
  NOR2X4 U75 ( .A(A[21]), .B(B[21]), .Y(n41) );
  CLKINVX3 U76 ( .A(n182), .Y(n106) );
  AND2X2 U77 ( .A(n190), .B(n191), .Y(n8) );
  OR2X2 U78 ( .A(A[7]), .B(B[7]), .Y(n210) );
  AND2X2 U79 ( .A(n64), .B(n49), .Y(n9) );
  AND2X2 U80 ( .A(n29), .B(n153), .Y(n10) );
  NOR2XL U81 ( .A(A[15]), .B(B[15]), .Y(n11) );
  NAND3BX1 U82 ( .AN(n13), .B(B[12]), .C(n205), .Y(n224) );
  NOR2X2 U83 ( .A(n248), .B(n16), .Y(n242) );
  NOR2X4 U84 ( .A(A[9]), .B(B[9]), .Y(n14) );
  NAND3X2 U85 ( .A(n63), .B(n256), .C(n257), .Y(n255) );
  XOR2X1 U86 ( .A(n103), .B(n108), .Y(SUM[29]) );
  NAND2X2 U87 ( .A(n109), .B(n110), .Y(n103) );
  NAND2X2 U88 ( .A(n24), .B(n164), .Y(n27) );
  NAND2XL U89 ( .A(n163), .B(n25), .Y(n26) );
  INVXL U90 ( .A(n163), .Y(n24) );
  NAND4BX2 U91 ( .AN(n14), .B(n64), .C(n249), .D(n250), .Y(n15) );
  NOR3BX4 U92 ( .AN(n201), .B(n202), .C(n203), .Y(n200) );
  NAND2X2 U93 ( .A(n74), .B(n75), .Y(n73) );
  NOR2BX4 U94 ( .AN(n179), .B(n173), .Y(n167) );
  NOR2X2 U95 ( .A(A[11]), .B(B[11]), .Y(n16) );
  CLKINVX4 U96 ( .A(n232), .Y(n17) );
  BUFX12 U97 ( .A(B[5]), .Y(n18) );
  AOI21X4 U98 ( .A0(n107), .A1(n182), .B0(n181), .Y(n262) );
  NOR3BX2 U99 ( .AN(n206), .B(n15), .C(n215), .Y(n214) );
  NOR2BX1 U100 ( .AN(n58), .B(n14), .Y(n57) );
  OR2X4 U101 ( .A(A[5]), .B(B[5]), .Y(n270) );
  OR2X4 U102 ( .A(A[5]), .B(B[5]), .Y(n45) );
  AOI21X2 U103 ( .A0(n198), .A1(n199), .B0(n200), .Y(n197) );
  NAND3X4 U104 ( .A(n204), .B(n209), .C(n210), .Y(n208) );
  OAI21X1 U105 ( .A0(B[14]), .A1(A[14]), .B0(n206), .Y(n202) );
  NOR2X2 U106 ( .A(n81), .B(n49), .Y(n79) );
  OAI2BB1X2 U107 ( .A0N(n71), .A1N(n49), .B0(n75), .Y(n82) );
  INVX2 U108 ( .A(n240), .Y(n239) );
  NAND2X2 U109 ( .A(B[12]), .B(A[12]), .Y(n240) );
  OAI2BB1X2 U110 ( .A0N(B[7]), .A1N(A[7]), .B0(n273), .Y(n267) );
  NOR2BX2 U111 ( .AN(n182), .B(n35), .Y(SUM[0]) );
  NAND2X4 U112 ( .A(n9), .B(n260), .Y(n257) );
  NOR2BX4 U113 ( .AN(n50), .B(n84), .Y(n83) );
  NAND2X2 U114 ( .A(n8), .B(n169), .Y(n189) );
  NAND2X4 U115 ( .A(n18), .B(A[5]), .Y(n74) );
  NAND3X1 U116 ( .A(n155), .B(n156), .C(n157), .Y(n143) );
  INVX1 U117 ( .A(n136), .Y(n125) );
  NAND2BX4 U118 ( .AN(n265), .B(n199), .Y(n61) );
  BUFX8 U119 ( .A(n276), .Y(SUM[4]) );
  OR2X4 U120 ( .A(A[27]), .B(B[27]), .Y(n130) );
  CLKINVX8 U121 ( .A(n215), .Y(n260) );
  NOR2X4 U122 ( .A(n160), .B(n151), .Y(n19) );
  OR2X4 U123 ( .A(n19), .B(n20), .Y(n158) );
  NAND2X4 U124 ( .A(B[22]), .B(A[22]), .Y(n149) );
  NAND3BX4 U125 ( .AN(n188), .B(n178), .C(n189), .Y(n186) );
  NAND2X4 U126 ( .A(n106), .B(n21), .Y(n22) );
  NAND2X2 U127 ( .A(n182), .B(n180), .Y(n23) );
  NAND2X4 U128 ( .A(n22), .B(n23), .Y(SUM[1]) );
  INVX3 U129 ( .A(n180), .Y(n21) );
  NAND2X4 U130 ( .A(n26), .B(n27), .Y(SUM[21]) );
  NOR2BXL U131 ( .AN(n153), .B(n41), .Y(n164) );
  NAND4BX4 U132 ( .AN(n265), .B(n45), .C(n70), .D(n71), .Y(n215) );
  OAI21X4 U133 ( .A0(n47), .A1(n101), .B0(n102), .Y(n97) );
  XOR2X2 U134 ( .A(n137), .B(n138), .Y(SUM[25]) );
  XOR2X4 U135 ( .A(n111), .B(n113), .Y(SUM[28]) );
  OAI21X2 U136 ( .A0(n115), .A1(n116), .B0(n117), .Y(n111) );
  OAI21X2 U137 ( .A0(n79), .A1(n80), .B0(n50), .Y(n76) );
  NOR2BX4 U138 ( .AN(n149), .B(n151), .Y(n162) );
  XOR2X4 U139 ( .A(n134), .B(n135), .Y(SUM[26]) );
  OAI2BB1X2 U140 ( .A0N(n136), .A1N(n137), .B0(n127), .Y(n134) );
  XOR2X4 U141 ( .A(n82), .B(n83), .Y(SUM[5]) );
  NOR2BX2 U142 ( .AN(n75), .B(n86), .Y(n85) );
  XOR2X4 U143 ( .A(n76), .B(n77), .Y(SUM[6]) );
  NAND2XL U144 ( .A(B[25]), .B(A[25]), .Y(n127) );
  NAND2X1 U145 ( .A(B[24]), .B(A[24]), .Y(n126) );
  OAI2BB1X4 U146 ( .A0N(n163), .A1N(n36), .B0(n153), .Y(n161) );
  INVX2 U147 ( .A(n157), .Y(n150) );
  OR2X2 U148 ( .A(A[24]), .B(B[24]), .Y(n140) );
  NOR2BXL U149 ( .AN(n128), .B(n122), .Y(n132) );
  NAND2X1 U150 ( .A(B[18]), .B(A[18]), .Y(n175) );
  NAND2XL U151 ( .A(B[23]), .B(A[23]), .Y(n154) );
  NOR2X4 U152 ( .A(n90), .B(n46), .Y(n263) );
  NOR2X2 U153 ( .A(n146), .B(n147), .Y(n145) );
  NOR2XL U154 ( .A(n41), .B(n44), .Y(n155) );
  NOR2BX1 U155 ( .AN(n152), .B(n44), .Y(n166) );
  INVX1 U156 ( .A(n130), .Y(n122) );
  NOR2X4 U157 ( .A(A[2]), .B(B[2]), .Y(n46) );
  NAND2X2 U158 ( .A(B[4]), .B(A[4]), .Y(n75) );
  NAND2X2 U159 ( .A(B[1]), .B(A[1]), .Y(n107) );
  NAND2X1 U160 ( .A(B[17]), .B(A[17]), .Y(n178) );
  NOR2X4 U161 ( .A(A[18]), .B(B[18]), .Y(n42) );
  BUFX8 U162 ( .A(n90), .Y(n53) );
  INVXL U163 ( .A(n112), .Y(n114) );
  NOR2BXL U164 ( .AN(n121), .B(n123), .Y(n135) );
  NOR2BXL U165 ( .AN(n127), .B(n125), .Y(n138) );
  NAND2XL U166 ( .A(n97), .B(n98), .Y(n96) );
  OR2X4 U167 ( .A(n151), .B(n10), .Y(n148) );
  INVXL U168 ( .A(n134), .Y(n133) );
  NOR2BX4 U169 ( .AN(n69), .B(n78), .Y(n77) );
  INVX1 U170 ( .A(n41), .Y(n36) );
  CLKINVX3 U171 ( .A(n221), .Y(n220) );
  NAND2X2 U172 ( .A(n61), .B(n62), .Y(n60) );
  NOR2BXL U173 ( .AN(n154), .B(n150), .Y(n159) );
  XOR2X4 U174 ( .A(n252), .B(n34), .Y(SUM[11]) );
  AND2X1 U175 ( .A(n247), .B(n249), .Y(n34) );
  NOR2XL U176 ( .A(n177), .B(n171), .Y(n188) );
  NOR2BXL U177 ( .AN(n179), .B(n43), .Y(n184) );
  OR2X4 U178 ( .A(A[4]), .B(B[4]), .Y(n71) );
  NOR2XL U179 ( .A(A[0]), .B(B[0]), .Y(n35) );
  NAND2XL U180 ( .A(B[27]), .B(A[27]), .Y(n128) );
  OR2X4 U181 ( .A(A[22]), .B(B[22]), .Y(n156) );
  NAND2XL U182 ( .A(B[30]), .B(A[30]), .Y(n95) );
  NAND2XL U183 ( .A(B[28]), .B(A[28]), .Y(n110) );
  INVXL U184 ( .A(A[7]), .Y(n52) );
  NAND2XL U185 ( .A(B[4]), .B(A[4]), .Y(n272) );
  INVXL U186 ( .A(A[5]), .Y(n55) );
  NAND3X2 U187 ( .A(n212), .B(n213), .C(n214), .Y(n196) );
  INVX1 U188 ( .A(n103), .Y(n101) );
  NAND3BX1 U189 ( .AN(n125), .B(n129), .C(n130), .Y(n116) );
  NOR2BX1 U190 ( .AN(n175), .B(n42), .Y(n187) );
  AND2X1 U191 ( .A(n178), .B(n190), .Y(n37) );
  NAND2XL U192 ( .A(n221), .B(n204), .Y(n226) );
  INVX1 U193 ( .A(n230), .Y(n229) );
  OAI21XL U194 ( .A0(n248), .A1(n58), .B0(n245), .Y(n253) );
  INVX1 U195 ( .A(n191), .Y(n172) );
  NAND2BX1 U196 ( .AN(n42), .B(n176), .Y(n174) );
  NAND2XL U197 ( .A(n63), .B(n64), .Y(n59) );
  XOR2X1 U198 ( .A(n139), .B(n141), .Y(n274) );
  NOR2BX1 U199 ( .AN(n126), .B(n142), .Y(n141) );
  INVX1 U200 ( .A(n140), .Y(n142) );
  NOR2BX1 U201 ( .AN(n95), .B(n100), .Y(n99) );
  INVX1 U202 ( .A(n98), .Y(n100) );
  NOR2BX1 U203 ( .AN(n110), .B(n114), .Y(n113) );
  XOR2X1 U204 ( .A(n165), .B(n166), .Y(SUM[20]) );
  AND2X1 U205 ( .A(n240), .B(n206), .Y(n38) );
  XOR2X1 U206 ( .A(n49), .B(n85), .Y(n276) );
  INVX1 U207 ( .A(n71), .Y(n86) );
  NOR2BX1 U208 ( .AN(n102), .B(n47), .Y(n108) );
  NOR2BX1 U209 ( .AN(n92), .B(n46), .Y(n104) );
  AOI21X1 U210 ( .A0(n120), .A1(n121), .B0(n122), .Y(n119) );
  NAND2BX1 U211 ( .AN(n123), .B(n124), .Y(n120) );
  OAI21XL U212 ( .A0(n125), .A1(n126), .B0(n127), .Y(n124) );
  AOI21X2 U213 ( .A0(n148), .A1(n149), .B0(n150), .Y(n147) );
  XNOR2X4 U214 ( .A(n258), .B(n39), .Y(SUM[10]) );
  AND2X1 U215 ( .A(n245), .B(n250), .Y(n39) );
  OAI2BB1X2 U216 ( .A0N(n105), .A1N(n106), .B0(n107), .Y(n93) );
  NOR2BX2 U217 ( .AN(n204), .B(n225), .Y(n218) );
  NOR2X2 U218 ( .A(n225), .B(n233), .Y(n213) );
  INVX1 U219 ( .A(n75), .Y(n81) );
  NAND2X2 U220 ( .A(n40), .B(n255), .Y(n254) );
  AND2X1 U221 ( .A(n250), .B(n251), .Y(n40) );
  INVX1 U222 ( .A(n154), .Y(n146) );
  INVX1 U223 ( .A(n177), .Y(n193) );
  INVX4 U224 ( .A(n264), .Y(n90) );
  BUFX3 U225 ( .A(n74), .Y(n50) );
  INVX1 U226 ( .A(B[7]), .Y(n51) );
  NOR2X4 U227 ( .A(A[19]), .B(B[19]), .Y(n43) );
  NAND2X2 U228 ( .A(B[8]), .B(A[8]), .Y(n63) );
  NAND2X2 U229 ( .A(B[9]), .B(A[9]), .Y(n58) );
  NAND2X1 U230 ( .A(B[10]), .B(A[10]), .Y(n245) );
  NAND2XL U231 ( .A(B[15]), .B(A[15]), .Y(n221) );
  NAND2XL U232 ( .A(B[14]), .B(A[14]), .Y(n223) );
  NAND2XL U233 ( .A(B[14]), .B(A[14]), .Y(n230) );
  OR2X2 U234 ( .A(A[26]), .B(B[26]), .Y(n129) );
  OR2X2 U235 ( .A(A[25]), .B(B[25]), .Y(n136) );
  NAND2X1 U236 ( .A(B[26]), .B(A[26]), .Y(n121) );
  NOR2X1 U237 ( .A(A[29]), .B(B[29]), .Y(n47) );
  NAND2X1 U238 ( .A(B[29]), .B(A[29]), .Y(n102) );
  OR2X2 U239 ( .A(A[28]), .B(B[28]), .Y(n112) );
  OR2X2 U240 ( .A(A[30]), .B(B[30]), .Y(n98) );
  XOR3X2 U241 ( .A(B[31]), .B(A[31]), .C(n94), .Y(SUM[31]) );
  NAND2X1 U242 ( .A(n95), .B(n96), .Y(n94) );
  NAND3BX4 U243 ( .AN(n261), .B(n89), .C(n217), .Y(n72) );
  NAND3X4 U244 ( .A(n196), .B(n197), .C(n195), .Y(n169) );
  NOR2X2 U245 ( .A(B[14]), .B(A[14]), .Y(n225) );
  BUFX4 U246 ( .A(n275), .Y(SUM[16]) );
  AOI21X2 U247 ( .A0(n191), .A1(n169), .B0(n193), .Y(n192) );
  NAND2X1 U248 ( .A(B[11]), .B(A[11]), .Y(n247) );
  AOI21X2 U249 ( .A0(n61), .A1(n62), .B0(n15), .Y(n241) );
  INVXL U250 ( .A(B[3]), .Y(n54) );
  NAND3BX4 U251 ( .AN(n55), .B(n70), .C(n18), .Y(n273) );
  NAND2X2 U252 ( .A(B[6]), .B(A[6]), .Y(n69) );
  CLKINVX8 U253 ( .A(n70), .Y(n78) );
  INVX3 U254 ( .A(n69), .Y(n271) );
  XOR2X1 U255 ( .A(n169), .B(n194), .Y(n275) );
  XOR2X4 U256 ( .A(n56), .B(n57), .Y(SUM[9]) );
  XNOR2X4 U257 ( .A(n59), .B(n60), .Y(SUM[8]) );
  XOR2X4 U258 ( .A(n65), .B(n66), .Y(SUM[7]) );
  XOR2X4 U259 ( .A(n87), .B(n88), .Y(SUM[3]) );
  NOR2BX4 U260 ( .AN(n89), .B(n53), .Y(n88) );
  XOR2X4 U261 ( .A(n131), .B(n132), .Y(SUM[27]) );
  OAI21X4 U262 ( .A0(n133), .A1(n123), .B0(n121), .Y(n131) );
  NAND2X4 U263 ( .A(n115), .B(n126), .Y(n137) );
  NAND2X4 U264 ( .A(n139), .B(n140), .Y(n115) );
  OAI21X4 U265 ( .A0(n143), .A1(n144), .B0(n145), .Y(n139) );
  XOR2X4 U266 ( .A(n158), .B(n159), .Y(SUM[23]) );
  OR2X4 U267 ( .A(A[23]), .B(B[23]), .Y(n157) );
  XOR2X4 U268 ( .A(n161), .B(n162), .Y(SUM[22]) );
  NAND2X4 U269 ( .A(n167), .B(n168), .Y(n165) );
  XOR2X4 U270 ( .A(n183), .B(n184), .Y(SUM[19]) );
  OAI21X4 U271 ( .A0(n185), .A1(n42), .B0(n175), .Y(n183) );
  XOR2X4 U272 ( .A(n186), .B(n187), .Y(SUM[18]) );
  NAND2X4 U273 ( .A(n204), .B(n205), .Y(n203) );
  NOR2X4 U274 ( .A(n207), .B(n208), .Y(n198) );
  AOI31X2 U275 ( .A0(n89), .A1(n216), .A2(n217), .B0(n11), .Y(n212) );
  XOR2X4 U276 ( .A(n226), .B(n227), .Y(SUM[15]) );
  OR2X4 U277 ( .A(A[15]), .B(B[15]), .Y(n204) );
  XOR2X4 U278 ( .A(n228), .B(n231), .Y(SUM[14]) );
  OR2X4 U279 ( .A(B[14]), .B(A[14]), .Y(n209) );
  OAI21X4 U280 ( .A0(n232), .A1(n233), .B0(n222), .Y(n228) );
  XOR2X4 U281 ( .A(n17), .B(n235), .Y(SUM[13]) );
  NOR2BX4 U282 ( .AN(n222), .B(n233), .Y(n235) );
  CLKINVX3 U283 ( .A(n205), .Y(n233) );
  OR2X4 U284 ( .A(A[13]), .B(B[13]), .Y(n205) );
  OAI2BB1X4 U285 ( .A0N(n236), .A1N(n237), .B0(n238), .Y(n234) );
  OAI2BB1X4 U286 ( .A0N(n242), .A1N(n243), .B0(n244), .Y(n201) );
  AOI2BB1X4 U287 ( .A0N(n16), .A1N(n245), .B0(n246), .Y(n244) );
  OR2X4 U288 ( .A(A[12]), .B(B[12]), .Y(n206) );
  OR2X4 U289 ( .A(A[11]), .B(B[11]), .Y(n249) );
  NAND2BX4 U290 ( .AN(n253), .B(n254), .Y(n252) );
  AOI21X4 U291 ( .A0(n251), .A1(n56), .B0(n259), .Y(n258) );
  NAND3X4 U292 ( .A(n256), .B(n63), .C(n257), .Y(n56) );
  NAND2X4 U293 ( .A(n262), .B(n263), .Y(n217) );
  OR2X4 U294 ( .A(A[1]), .B(B[1]), .Y(n105) );
  NAND2BX4 U295 ( .AN(n92), .B(n264), .Y(n216) );
  OR2X4 U296 ( .A(A[3]), .B(B[3]), .Y(n264) );
  NAND2X4 U297 ( .A(B[2]), .B(A[2]), .Y(n92) );
  NOR2X4 U298 ( .A(A[7]), .B(B[7]), .Y(n265) );
  NAND2BX4 U299 ( .AN(n266), .B(n199), .Y(n256) );
  NAND2BX4 U300 ( .AN(n267), .B(n268), .Y(n199) );
  AOI21X4 U301 ( .A0(n269), .A1(n270), .B0(n271), .Y(n268) );
  NOR2X4 U302 ( .A(n78), .B(n272), .Y(n269) );
  OR2X4 U303 ( .A(B[6]), .B(A[6]), .Y(n70) );
  OR2X4 U304 ( .A(B[8]), .B(A[8]), .Y(n64) );
  OR2X4 U305 ( .A(A[10]), .B(B[10]), .Y(n250) );
endmodule


module hash_core ( clk, reset, Wt, inner_busy, first_block_core, output_enable, 
        digest, output_valid );
  input [31:0] Wt;
  output [3:0] digest;
  input clk, reset, inner_busy, first_block_core, output_enable;
  output output_valid;
  wire   N177, N178, N179, N180, N181, N182, N183, N851, N852, N853, N854,
         N855, N856, N857, N858, N859, N860, N861, N862, N863, N864, N865,
         N866, N867, N868, N869, N870, N871, N872, N873, N874, N875, N876,
         N877, N878, N879, N880, N881, N882, N883, N884, N885, N886, N887,
         N888, N889, N890, N891, N892, N893, N894, N895, N896, N897, N898,
         N899, N900, N901, N902, N903, N904, N905, N906, N907, N908, N909,
         N910, N911, N912, N913, N914, N915, N916, N917, N918, N919, N920,
         N921, N922, N923, N924, N925, N926, N927, N928, N929, N930, N931,
         N932, N933, N934, N935, N936, N937, N938, N939, N940, N941, N942,
         N943, N944, N945, N946, N947, N948, N949, N950, N951, N952, N953,
         N954, N955, N956, N957, N958, N959, N960, N961, N962, N963, N964,
         N965, N966, N967, N968, N969, N970, N971, N972, N973, N974, N975,
         N976, N977, N978, N979, N980, N981, N982, N983, N984, N985, N986,
         N987, N988, N989, N990, N991, N992, N993, N994, N995, N996, N997,
         N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006, N1007,
         N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1017,
         N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027,
         N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036, N1037,
         N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046, N1047,
         N1048, N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056, N1057,
         N1058, N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066, N1067,
         N1068, N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076, N1077,
         N1078, N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086, N1087,
         N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096, N1097,
         N1098, N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106, N3002,
         N3003, N3004, N3005, N3006, N3007, N3008, N3009, N3010, N3011, N3012,
         N3013, N3014, N3015, N3016, N3017, N3018, N3019, N3020, N3021, N3022,
         N3023, N3024, N3025, N3026, N3027, N3028, N3029, N3030, N3031, N3032,
         N3033, N3433, N3434, N3435, N3444, N3445, N3446, N3447, N3448, N3449,
         N3450, N3451, N3452, N3453, n1337, n1371, n1384, n1389, n1397, n1434,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1456, n1457,
         n1458, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1487, n1488, n1489, n1490,
         n1491, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1611, n1612, n1615, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1631, n1632, n1633,
         n1635, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1720,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1755,
         n1756, n1757, n1758, n1759, n1760, n1763, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1785, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1849, n1859, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1878, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2179, n2180, n2181,
         n2183, n2184, n2185, n2186, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2239, n2240, n2241, n2242, n2244, n2245, n2247,
         n2248, n2249, n2250, n2251, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, T2_32_9_,
         T2_32_8_, T2_32_7_, T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_, T2_32_31_,
         T2_32_30_, T2_32_2_, T2_32_29_, T2_32_28_, T2_32_27_, T2_32_26_,
         T2_32_25_, T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_, T2_32_20_,
         T2_32_1_, T2_32_19_, T2_32_18_, T2_32_17_, T2_32_16_, T2_32_15_,
         T2_32_14_, T2_32_13_, T2_32_12_, T2_32_11_, T2_32_10_, T2_32_0_, N99,
         N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85,
         N84, N83, N82, N81, N80, N175, N174, N173, N172, N171, N170, N169,
         N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158,
         N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147,
         N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136,
         N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125,
         N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114,
         N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103,
         N102, N101, N100, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n112, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950;
  wire   [31:0] f1_EFG_32;
  wire   [31:0] f2_ABC_32;
  wire   [31:0] f3_A_32;
  wire   [31:0] f4_E_32;
  wire   [31:0] Kt;
  wire   [31:0] T1_32;
  wire   [31:0] next_E;
  wire   [31:0] next_A;
  wire   [255:0] SHA256_result;
  wire   [6:0] round;
  wire   [31:0] H0;
  wire   [31:1] H1;
  wire   [31:0] H2;
  wire   [31:1] H3;
  wire   [31:0] H4;
  wire   [31:0] H5;
  wire   [31:2] H6;
  wire   [31:0] H7;
  wire   [5:0] read_counter;

  DFFHQX4 B_reg_0_ ( .D(n2954), .CK(clk), .Q(SHA256_result[192]) );
  DFFHQX4 E_reg_0_ ( .D(n2857), .CK(clk), .Q(SHA256_result[96]) );
  DFFHQX4 E_reg_1_ ( .D(n2856), .CK(clk), .Q(SHA256_result[97]) );
  DFFHQX4 E_reg_2_ ( .D(n2855), .CK(clk), .Q(SHA256_result[98]) );
  DFFHQX4 E_reg_4_ ( .D(n2853), .CK(clk), .Q(SHA256_result[100]) );
  DFFHQX4 E_reg_7_ ( .D(n2850), .CK(clk), .Q(SHA256_result[103]) );
  DFFHQX4 E_reg_11_ ( .D(n2846), .CK(clk), .Q(SHA256_result[107]) );
  DFFHQX4 E_reg_13_ ( .D(n2844), .CK(clk), .Q(SHA256_result[109]) );
  DFFHQX4 F_reg_2_ ( .D(n2823), .CK(clk), .Q(SHA256_result[66]) );
  DFFHQX4 F_reg_3_ ( .D(n2822), .CK(clk), .Q(SHA256_result[67]) );
  DFFHQX4 G_reg_1_ ( .D(n2633), .CK(clk), .Q(SHA256_result[33]) );
  DFFHQX4 G_reg_3_ ( .D(n2631), .CK(clk), .Q(SHA256_result[35]) );
  DFFHQX4 Kt_reg_8_ ( .D(N3010), .CK(clk), .Q(Kt[8]) );
  DFFHQX4 Kt_reg_3_ ( .D(N3005), .CK(clk), .Q(Kt[3]) );
  DFFHQX4 Kt_reg_2_ ( .D(N3004), .CK(clk), .Q(Kt[2]) );
  DFFHQX4 Kt_reg_1_ ( .D(N3003), .CK(clk), .Q(Kt[1]) );
  DFFHQX4 Kt_reg_0_ ( .D(N3002), .CK(clk), .Q(Kt[0]) );
  AND2X2 U1332 ( .A(n2177), .B(n51), .Y(n1989) );
  AND2X2 U1333 ( .A(n2179), .B(n51), .Y(n1988) );
  AND2X2 U1335 ( .A(n2180), .B(n51), .Y(n1991) );
  AND2X2 U1336 ( .A(n2181), .B(n51), .Y(n1990) );
  AND2X2 U1338 ( .A(n2177), .B(n50), .Y(n1993) );
  AND2X2 U1339 ( .A(n2179), .B(n50), .Y(n1992) );
  AND2X2 U1341 ( .A(n2180), .B(n50), .Y(n1995) );
  AND2X2 U1342 ( .A(n2181), .B(n50), .Y(n1994) );
  AND2X2 U1345 ( .A(n2177), .B(n48), .Y(n2001) );
  AND2X2 U1346 ( .A(n2179), .B(n48), .Y(n2000) );
  AND2X2 U1348 ( .A(n2180), .B(n48), .Y(n2003) );
  AND2X2 U1349 ( .A(n2181), .B(n48), .Y(n2002) );
  AND2X2 U1351 ( .A(n2177), .B(n49), .Y(n2005) );
  AND2X2 U1352 ( .A(n2189), .B(n2190), .Y(n2177) );
  AND2X2 U1353 ( .A(n2179), .B(n49), .Y(n2004) );
  AND2X2 U1354 ( .A(n2189), .B(n2191), .Y(n2179) );
  AND2X2 U1356 ( .A(n2180), .B(n49), .Y(n2007) );
  AND2X2 U1357 ( .A(n2192), .B(n2190), .Y(n2180) );
  AND2X2 U1358 ( .A(n2181), .B(n49), .Y(n2006) );
  AND2X2 U1359 ( .A(n2192), .B(n2191), .Y(n2181) );
  AND2X2 U1362 ( .A(n51), .B(n2197), .Y(n2013) );
  AND2X2 U1363 ( .A(n51), .B(n2198), .Y(n2012) );
  AND2X2 U1365 ( .A(n51), .B(n2199), .Y(n2015) );
  AND2X2 U1366 ( .A(n51), .B(n2200), .Y(n2014) );
  AND2X2 U1368 ( .A(n50), .B(n2197), .Y(n2017) );
  AND2X2 U1369 ( .A(n50), .B(n2198), .Y(n2016) );
  AND2X2 U1371 ( .A(n50), .B(n2199), .Y(n2019) );
  AND2X2 U1372 ( .A(n50), .B(n2200), .Y(n2018) );
  AND2X2 U1375 ( .A(n2197), .B(n48), .Y(n2024) );
  AND2X2 U1376 ( .A(n48), .B(n2198), .Y(n1977) );
  AND2X2 U1378 ( .A(n2199), .B(n48), .Y(n2026) );
  AND2X2 U1379 ( .A(n2200), .B(n48), .Y(n2025) );
  AND2X2 U1381 ( .A(n49), .B(n2197), .Y(n2028) );
  AND2X2 U1382 ( .A(n2190), .B(n2205), .Y(n2197) );
  AND2X2 U1383 ( .A(n49), .B(n2198), .Y(n2027) );
  AND2X2 U1384 ( .A(n2191), .B(n2205), .Y(n2198) );
  AND2X2 U1386 ( .A(n49), .B(n2199), .Y(n2030) );
  AND2X2 U1387 ( .A(n2206), .B(n2190), .Y(n2199) );
  AND2X2 U1388 ( .A(read_counter[0]), .B(n950), .Y(n2190) );
  AND2X2 U1389 ( .A(n49), .B(n2200), .Y(n2029) );
  AND2X2 U1390 ( .A(n2206), .B(n2191), .Y(n2200) );
  AND2X2 U1395 ( .A(n2215), .B(n51), .Y(n2040) );
  AND2X2 U1396 ( .A(n2216), .B(n51), .Y(n2039) );
  AND2X2 U1398 ( .A(n2217), .B(n51), .Y(n2042) );
  AND2X2 U1399 ( .A(n2218), .B(n51), .Y(n2041) );
  AND2X2 U1401 ( .A(n2215), .B(n50), .Y(n2044) );
  AND2X2 U1402 ( .A(n2216), .B(n50), .Y(n2043) );
  AND2X2 U1404 ( .A(n2217), .B(n50), .Y(n2046) );
  AND2X2 U1405 ( .A(n2218), .B(n50), .Y(n2045) );
  AND2X2 U1408 ( .A(n2215), .B(n48), .Y(n2052) );
  AND2X2 U1409 ( .A(n2216), .B(n48), .Y(n2051) );
  AND2X2 U1411 ( .A(n2217), .B(n48), .Y(n2054) );
  AND2X2 U1412 ( .A(n2218), .B(n48), .Y(n2053) );
  AND2X2 U1414 ( .A(n2215), .B(n49), .Y(n2056) );
  AND2X2 U1415 ( .A(n2223), .B(n2189), .Y(n2215) );
  AND2X2 U1416 ( .A(n2216), .B(n49), .Y(n2055) );
  AND2X2 U1417 ( .A(n2224), .B(n2189), .Y(n2216) );
  AND2X2 U1418 ( .A(read_counter[4]), .B(n948), .Y(n2189) );
  AND2X2 U1420 ( .A(n2217), .B(n49), .Y(n2058) );
  AND2X2 U1421 ( .A(n2223), .B(n2192), .Y(n2217) );
  AND2X2 U1422 ( .A(n2218), .B(n49), .Y(n2057) );
  AND2X2 U1423 ( .A(n2224), .B(n2192), .Y(n2218) );
  AND2X2 U1424 ( .A(read_counter[4]), .B(read_counter[1]), .Y(n2192) );
  AND2X2 U1427 ( .A(n2229), .B(n51), .Y(n2064) );
  AND2X2 U1428 ( .A(n2230), .B(n51), .Y(n2063) );
  AND2X2 U1430 ( .A(n2231), .B(n51), .Y(n2066) );
  AND2X2 U1431 ( .A(n2232), .B(n51), .Y(n2065) );
  AND2X2 U1434 ( .A(n2229), .B(n50), .Y(n2068) );
  AND2X2 U1435 ( .A(n2230), .B(n50), .Y(n2067) );
  AND2X2 U1437 ( .A(n2231), .B(n50), .Y(n2070) );
  AND2X2 U1438 ( .A(n2232), .B(n50), .Y(n2069) );
  AND2X2 U1442 ( .A(n2229), .B(n48), .Y(n2076) );
  AND2X2 U1443 ( .A(n2230), .B(n48), .Y(n2075) );
  AND2X2 U1445 ( .A(n2231), .B(n48), .Y(n2078) );
  AND2X2 U1446 ( .A(n2232), .B(n48), .Y(n2077) );
  AND2X2 U1449 ( .A(n2229), .B(n49), .Y(n2080) );
  AND2X2 U1450 ( .A(n2223), .B(n2205), .Y(n2229) );
  AND2X2 U1451 ( .A(n2230), .B(n49), .Y(n2079) );
  AND2X2 U1452 ( .A(n2224), .B(n2205), .Y(n2230) );
  AND2X2 U1455 ( .A(n2231), .B(n49), .Y(n2082) );
  AND2X2 U1456 ( .A(n2223), .B(n2206), .Y(n2231) );
  AND2X2 U1457 ( .A(read_counter[0]), .B(read_counter[5]), .Y(n2223) );
  AND2X2 U1458 ( .A(n2232), .B(n49), .Y(n2081) );
  AND2X2 U1460 ( .A(n2224), .B(n2206), .Y(n2232) );
  AND2X2 U1523 ( .A(n2355), .B(n330), .Y(n2294) );
  CLKINVX4 U2120 ( .A(reset), .Y(n1434) );
  hash_core_DW01_add_0 add_318 ( .A({SHA256_result[63:33], n95}), .B({H7[31:2], 
        n109, H7[0]}), .SUM({N1106, N1105, N1104, N1103, N1102, N1101, N1100, 
        N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, 
        N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, 
        N1079, N1078, N1077, N1076, N1075}) );
  hash_core_DW01_add_1 add_317 ( .A({SHA256_result[95:66], n115, n107}), .B({
        H6, n110, n114}), .SUM({N1074, N1073, N1072, N1071, N1070, N1069, 
        N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, 
        N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, 
        N1048, N1047, N1046, N1045, N1044, N1043}) );
  hash_core_DW01_add_2 add_316 ( .A({SHA256_result[127], n145, 
        SHA256_result[125:124], n73, SHA256_result[122:118], n146, 
        SHA256_result[116], n147, SHA256_result[114], n148, SHA256_result[112], 
        n149, SHA256_result[110:109], n150, SHA256_result[107], n151, n152, 
        n153, SHA256_result[103], n154, SHA256_result[101:98], n74, n76}), .B(
        H5), .SUM({N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, 
        N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, 
        N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, 
        N1014, N1013, N1012, N1011}) );
  hash_core_DW01_add_4 add_314 ( .A({SHA256_result[191:162], n86, n89}), .B({
        H3, n112}), .SUM({N978, N977, N976, N975, N974, N973, N972, N971, N970, 
        N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, 
        N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947}) );
  hash_core_DW01_add_5 add_313 ( .A(SHA256_result[223:192]), .B(H2), .SUM({
        N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, 
        N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, 
        N922, N921, N920, N919, N918, N917, N916, N915}) );
  hash_core_DW01_add_6 add_312 ( .A({SHA256_result[255], n155, n156, 
        SHA256_result[252], n157, n158, n159, n160, n161, n37, n162, n163, 
        n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
        n176, n177, n178, n179, n180, n181, n71, n92}), .B({H1, n91}), .SUM({
        N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, 
        N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, 
        N890, N889, N888, N887, N886, N885, N884, N883}) );
  hash_core_DW01_inc_0 add_120 ( .A({round[6], n183, n182, round[3:2], n335, 
        round[0]}), .SUM({N183, N182, N181, N180, N179, N178, N177}) );
  hash_core_DW01_add_15 add_315 ( .A(next_E), .B(H4), .SUM({N1010, N1009, 
        N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, 
        N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, 
        N986, N985, N984, N983, N982, N981, N980, N979}) );
  hash_core_DW01_add_16 add_311 ( .A(next_A), .B(H0), .SUM({N882, N881, N880, 
        N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, 
        N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, 
        N855, N854, N853, N852, N851}) );
  hash_core_DW01_add_20 add_1_root_add_0_root_add_114 ( .A(f2_ABC_32), .B(
        f3_A_32), .SUM({T2_32_31_, T2_32_30_, T2_32_29_, T2_32_28_, T2_32_27_, 
        T2_32_26_, T2_32_25_, T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_, 
        T2_32_20_, T2_32_19_, T2_32_18_, T2_32_17_, T2_32_16_, T2_32_15_, 
        T2_32_14_, T2_32_13_, T2_32_12_, T2_32_11_, T2_32_10_, T2_32_9_, 
        T2_32_8_, T2_32_7_, T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_, T2_32_2_, 
        T2_32_1_, T2_32_0_}) );
  hash_core_DW01_add_19 add_0_root_add_0_root_add_109_4 ( .A({N175, N174, N173, 
        N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, 
        N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, 
        N148, N147, N146, N145, N144}), .B({N143, N142, N141, N140, N139, N138, 
        N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, 
        N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, 
        N113, N112}), .SUM(T1_32) );
  hash_core_DW01_add_26 add_113 ( .A(SHA256_result[159:128]), .B({T1_32[31:27], 
        n55, T1_32[25:23], n56, T1_32[21:0]}), .SUM(next_E) );
  hash_core_DW01_add_27 add_0_root_add_0_root_add_114 ( .A({T2_32_31_, 
        T2_32_30_, T2_32_29_, T2_32_28_, T2_32_27_, T2_32_26_, T2_32_25_, 
        T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_, T2_32_20_, T2_32_19_, 
        T2_32_18_, T2_32_17_, T2_32_16_, T2_32_15_, T2_32_14_, T2_32_13_, 
        T2_32_12_, T2_32_11_, T2_32_10_, T2_32_9_, T2_32_8_, T2_32_7_, 
        T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_, T2_32_2_, T2_32_1_, T2_32_0_}), 
        .B({T1_32[31:27], n55, T1_32[25:23], n56, T1_32[21:0]}), .SUM(next_A)
         );
  hash_core_DW01_add_30 add_2_root_add_0_root_add_109_4 ( .A(
        SHA256_result[31:0]), .B({f1_EFG_32[31:3], n45, f1_EFG_32[1:0]}), 
        .SUM({N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, 
        N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, 
        N152, N151, N150, N149, N148, N147, N146, N145, N144}) );
  hash_core_DW01_add_32 add_3_root_add_0_root_add_109_4 ( .A(Kt), .B(Wt), 
        .SUM({N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, 
        N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, 
        N86, N85, N84, N83, N82, N81, N80}) );
  hash_core_DW01_add_38 add_1_root_add_0_root_add_109_4 ( .A(f4_E_32), .B({
        N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, 
        N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, 
        N85, N84, N83, N82, N81, N80}), .SUM({N143, N142, N141, N140, N139, 
        N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, 
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113, N112}) );
  DFFHQXL A_reg_30_ ( .D(n2988), .CK(clk), .Q(SHA256_result[254]) );
  DFFHQX1 read_counter_reg_3_ ( .D(N3451), .CK(clk), .Q(read_counter[3]) );
  DFFHQX1 read_counter_reg_5_ ( .D(N3453), .CK(clk), .Q(read_counter[5]) );
  DFFHQX1 read_counter_reg_1_ ( .D(N3449), .CK(clk), .Q(read_counter[1]) );
  DFFHQX1 read_counter_reg_2_ ( .D(N3450), .CK(clk), .Q(read_counter[2]) );
  DFFHQX1 read_counter_reg_4_ ( .D(N3452), .CK(clk), .Q(read_counter[4]) );
  DFFHQX1 read_counter_reg_0_ ( .D(N3448), .CK(clk), .Q(read_counter[0]) );
  DFFHQX1 Kt_reg_31_ ( .D(N3033), .CK(clk), .Q(Kt[31]) );
  DFFTRX1 round_reg_6_ ( .D(N183), .RN(n141), .CK(clk), .Q(round[6]), .QN(
        n1337) );
  DFFHQX1 Kt_reg_30_ ( .D(N3032), .CK(clk), .Q(Kt[30]) );
  DFFHQX1 Kt_reg_29_ ( .D(N3031), .CK(clk), .Q(Kt[29]) );
  DFFHQX1 Kt_reg_28_ ( .D(N3030), .CK(clk), .Q(Kt[28]) );
  DFFHQX1 Kt_reg_27_ ( .D(N3029), .CK(clk), .Q(Kt[27]) );
  DFFHQX1 Kt_reg_26_ ( .D(N3028), .CK(clk), .Q(Kt[26]) );
  DFFHQX1 Kt_reg_25_ ( .D(N3027), .CK(clk), .Q(Kt[25]) );
  DFFHQX1 Kt_reg_24_ ( .D(N3026), .CK(clk), .Q(Kt[24]) );
  DFFHQX1 Kt_reg_23_ ( .D(N3025), .CK(clk), .Q(Kt[23]) );
  DFFHQX1 G_reg_21_ ( .D(n2613), .CK(clk), .Q(SHA256_result[53]) );
  DFFHQX1 D_reg_1_ ( .D(n2888), .CK(clk), .Q(SHA256_result[129]) );
  DFFHQX1 H_reg_16_ ( .D(n2586), .CK(clk), .Q(SHA256_result[16]) );
  DFFHQX1 C_reg_12_ ( .D(n2909), .CK(clk), .Q(SHA256_result[172]) );
  DFFHQX1 C_reg_13_ ( .D(n2908), .CK(clk), .Q(SHA256_result[173]) );
  DFFHQX1 C_reg_10_ ( .D(n2911), .CK(clk), .Q(SHA256_result[170]) );
  DFFHQX1 F_reg_20_ ( .D(n2805), .CK(clk), .Q(SHA256_result[84]) );
  DFFHQX1 F_reg_21_ ( .D(n2804), .CK(clk), .Q(SHA256_result[85]) );
  DFFHQX1 B_reg_12_ ( .D(n2942), .CK(clk), .Q(SHA256_result[204]) );
  DFFHQX1 B_reg_13_ ( .D(n2941), .CK(clk), .Q(SHA256_result[205]) );
  DFFHQX1 B_reg_14_ ( .D(n2940), .CK(clk), .Q(SHA256_result[206]) );
  DFFHQX1 G_reg_20_ ( .D(n2614), .CK(clk), .Q(SHA256_result[52]) );
  DFFHQX1 C_reg_11_ ( .D(n2910), .CK(clk), .Q(SHA256_result[171]) );
  DFFHQX1 A_reg_6_ ( .D(n3012), .CK(clk), .Q(SHA256_result[230]) );
  DFFHQX1 A_reg_23_ ( .D(n2995), .CK(clk), .Q(SHA256_result[247]) );
  DFFHQX1 A_reg_24_ ( .D(n2994), .CK(clk), .Q(SHA256_result[248]) );
  DFFHQXL A_reg_25_ ( .D(n2993), .CK(clk), .Q(SHA256_result[249]) );
  DFFHQXL A_reg_26_ ( .D(n2992), .CK(clk), .Q(SHA256_result[250]) );
  DFFHQXL A_reg_27_ ( .D(n2991), .CK(clk), .Q(SHA256_result[251]) );
  DFFHQXL A_reg_29_ ( .D(n2989), .CK(clk), .Q(SHA256_result[253]) );
  DFFHQX1 Kt_reg_22_ ( .D(N3024), .CK(clk), .Q(Kt[22]) );
  DFFHQX1 Kt_reg_21_ ( .D(N3023), .CK(clk), .Q(Kt[21]) );
  DFFHQX1 Kt_reg_20_ ( .D(N3022), .CK(clk), .Q(Kt[20]) );
  DFFHQX1 Kt_reg_19_ ( .D(N3021), .CK(clk), .Q(Kt[19]) );
  DFFHQX1 H6_reg_4_ ( .D(n2661), .CK(clk), .Q(H6[4]) );
  DFFHQX1 F_reg_14_ ( .D(n2811), .CK(clk), .Q(SHA256_result[78]) );
  DFFHQX1 F_reg_15_ ( .D(n2810), .CK(clk), .Q(SHA256_result[79]) );
  DFFHQX1 F_reg_16_ ( .D(n2809), .CK(clk), .Q(SHA256_result[80]) );
  DFFHQX1 F_reg_17_ ( .D(n2808), .CK(clk), .Q(SHA256_result[81]) );
  DFFHQX1 G_reg_15_ ( .D(n2619), .CK(clk), .Q(SHA256_result[47]) );
  DFFHQX1 H_reg_15_ ( .D(n2587), .CK(clk), .Q(SHA256_result[15]) );
  DFFHQX1 H_reg_17_ ( .D(n2585), .CK(clk), .Q(SHA256_result[17]) );
  DFFHQX1 C_reg_5_ ( .D(n2916), .CK(clk), .Q(SHA256_result[165]) );
  DFFHQX1 C_reg_8_ ( .D(n2913), .CK(clk), .Q(SHA256_result[168]) );
  DFFHQX1 B_reg_5_ ( .D(n2949), .CK(clk), .Q(SHA256_result[197]) );
  DFFHQX1 B_reg_6_ ( .D(n2948), .CK(clk), .Q(SHA256_result[198]) );
  DFFHQX1 F_reg_18_ ( .D(n2807), .CK(clk), .Q(SHA256_result[82]) );
  DFFHQX1 B_reg_8_ ( .D(n2946), .CK(clk), .Q(SHA256_result[200]) );
  DFFHQX1 B_reg_9_ ( .D(n2945), .CK(clk), .Q(SHA256_result[201]) );
  DFFHQX1 G_reg_16_ ( .D(n2618), .CK(clk), .Q(SHA256_result[48]) );
  DFFHQX1 G_reg_17_ ( .D(n2617), .CK(clk), .Q(SHA256_result[49]) );
  DFFHQX1 B_reg_11_ ( .D(n2943), .CK(clk), .Q(SHA256_result[203]) );
  DFFHQX1 A_reg_3_ ( .D(n3015), .CK(clk), .Q(SHA256_result[227]) );
  DFFHQX1 A_reg_4_ ( .D(n3014), .CK(clk), .Q(SHA256_result[228]) );
  DFFHQX1 A_reg_5_ ( .D(n3013), .CK(clk), .Q(SHA256_result[229]) );
  DFFHQX1 E_reg_10_ ( .D(n2847), .CK(clk), .Q(SHA256_result[106]) );
  DFFHQX1 E_reg_19_ ( .D(n2838), .CK(clk), .Q(SHA256_result[115]) );
  DFFHQXL E_reg_30_ ( .D(n2827), .CK(clk), .Q(SHA256_result[126]) );
  DFFHQX1 Kt_reg_18_ ( .D(N3020), .CK(clk), .Q(Kt[18]) );
  DFFHQX1 Kt_reg_17_ ( .D(N3019), .CK(clk), .Q(Kt[17]) );
  DFFHQX1 Kt_reg_16_ ( .D(N3018), .CK(clk), .Q(Kt[16]) );
  DFFHQX1 H3_reg_2_ ( .D(n2727), .CK(clk), .Q(H3[2]) );
  DFFHQX1 H7_reg_2_ ( .D(n2568), .CK(clk), .Q(H7[2]) );
  DFFHQX1 H2_reg_2_ ( .D(n2696), .CK(clk), .Q(H2[2]) );
  DFFHQX1 H_reg_3_ ( .D(n2599), .CK(clk), .Q(SHA256_result[3]) );
  DFFHQX1 H_reg_11_ ( .D(n2591), .CK(clk), .Q(SHA256_result[11]) );
  DFFHQX1 C_reg_4_ ( .D(n2917), .CK(clk), .Q(SHA256_result[164]) );
  DFFHQX1 B_reg_4_ ( .D(n2950), .CK(clk), .Q(SHA256_result[196]) );
  DFFHQX1 E_reg_23_ ( .D(n2834), .CK(clk), .Q(SHA256_result[119]) );
  DFFTRX1 output_valid_reg ( .D(output_enable), .RN(n1434), .CK(clk), .Q(
        output_valid) );
  DFFHQX1 digest_reg_3_ ( .D(N3447), .CK(clk), .Q(digest[3]) );
  DFFHQX1 digest_reg_2_ ( .D(N3446), .CK(clk), .Q(digest[2]) );
  DFFHQX1 digest_reg_1_ ( .D(N3445), .CK(clk), .Q(digest[1]) );
  DFFHQX1 digest_reg_0_ ( .D(N3444), .CK(clk), .Q(digest[0]) );
  DFFHQXL H2_reg_11_ ( .D(n2687), .CK(clk), .Q(H2[11]) );
  DFFHQXL H3_reg_11_ ( .D(n2718), .CK(clk), .Q(H3[11]) );
  DFFHQXL H5_reg_10_ ( .D(n2783), .CK(clk), .Q(H5[10]) );
  DFFHQXL H2_reg_10_ ( .D(n2688), .CK(clk), .Q(H2[10]) );
  DFFHQXL H3_reg_10_ ( .D(n2719), .CK(clk), .Q(H3[10]) );
  DFFHQXL H_reg_23_ ( .D(n2579), .CK(clk), .Q(SHA256_result[23]) );
  DFFHQXL H_reg_21_ ( .D(n2581), .CK(clk), .Q(SHA256_result[21]) );
  DFFHQXL E_reg_21_ ( .D(n2836), .CK(clk), .Q(SHA256_result[117]) );
  DFFHQXL A_reg_21_ ( .D(n2997), .CK(clk), .Q(SHA256_result[245]) );
  DFFHQXL A_reg_10_ ( .D(n3008), .CK(clk), .Q(SHA256_result[234]) );
  DFFHQXL A_reg_12_ ( .D(n3006), .CK(clk), .Q(SHA256_result[236]) );
  DFFHQXL A_reg_11_ ( .D(n3007), .CK(clk), .Q(SHA256_result[235]) );
  DFFHQXL E_reg_17_ ( .D(n2840), .CK(clk), .Q(SHA256_result[113]) );
  DFFHQXL H3_reg_9_ ( .D(n2720), .CK(clk), .Q(H3[9]) );
  DFFHQXL H1_reg_8_ ( .D(n2978), .CK(clk), .Q(H1[8]) );
  DFFHQXL H2_reg_7_ ( .D(n2691), .CK(clk), .Q(H2[7]) );
  DFFHQXL H3_reg_7_ ( .D(n2722), .CK(clk), .Q(H3[7]) );
  DFFHQXL D_reg_0_ ( .D(n2889), .CK(clk), .Q(SHA256_result[128]) );
  DFFHQXL A_reg_9_ ( .D(n3009), .CK(clk), .Q(SHA256_result[233]) );
  DFFHQXL A_reg_18_ ( .D(n3000), .CK(clk), .Q(SHA256_result[242]) );
  DFFHQXL A_reg_20_ ( .D(n2998), .CK(clk), .Q(SHA256_result[244]) );
  DFFHQXL A_reg_16_ ( .D(n3002), .CK(clk), .Q(SHA256_result[240]) );
  DFFHQXL A_reg_17_ ( .D(n3001), .CK(clk), .Q(SHA256_result[241]) );
  DFFHQXL A_reg_8_ ( .D(n3010), .CK(clk), .Q(SHA256_result[232]) );
  DFFHQXL A_reg_19_ ( .D(n2999), .CK(clk), .Q(SHA256_result[243]) );
  DFFHQXL A_reg_15_ ( .D(n3003), .CK(clk), .Q(SHA256_result[239]) );
  DFFHQXL H5_reg_6_ ( .D(n2787), .CK(clk), .Q(H5[6]) );
  DFFHQXL H1_reg_6_ ( .D(n2980), .CK(clk), .Q(H1[6]) );
  DFFHQXL H2_reg_5_ ( .D(n2693), .CK(clk), .Q(H2[5]) );
  DFFHQXL H3_reg_5_ ( .D(n2724), .CK(clk), .Q(H3[5]) );
  DFFHQXL H5_reg_4_ ( .D(n2789), .CK(clk), .Q(H5[4]) );
  DFFHQXL H7_reg_4_ ( .D(n2566), .CK(clk), .Q(H7[4]) );
  DFFHQXL A_reg_13_ ( .D(n3005), .CK(clk), .Q(SHA256_result[237]) );
  DFFHQXL A_reg_14_ ( .D(n3004), .CK(clk), .Q(SHA256_result[238]) );
  DFFHQXL E_reg_15_ ( .D(n2842), .CK(clk), .Q(SHA256_result[111]) );
  DFFHQXL H2_reg_3_ ( .D(n2695), .CK(clk), .Q(H2[3]) );
  DFFHQXL H3_reg_3_ ( .D(n2726), .CK(clk), .Q(H3[3]) );
  DFFHQX1 H_reg_18_ ( .D(n2584), .CK(clk), .Q(SHA256_result[18]) );
  DFFHQX1 H_reg_19_ ( .D(n2583), .CK(clk), .Q(SHA256_result[19]) );
  DFFHQX1 H2_reg_6_ ( .D(n2692), .CK(clk), .Q(H2[6]) );
  DFFHQX1 H5_reg_5_ ( .D(n2788), .CK(clk), .Q(H5[5]) );
  DFFHQX1 H6_reg_5_ ( .D(n2660), .CK(clk), .Q(H6[5]) );
  DFFHQX1 H_reg_7_ ( .D(n2595), .CK(clk), .Q(SHA256_result[7]) );
  DFFHQX1 H_reg_5_ ( .D(n2597), .CK(clk), .Q(SHA256_result[5]) );
  DFFHQX1 C_reg_7_ ( .D(n2914), .CK(clk), .Q(SHA256_result[167]) );
  DFFHQX1 H1_reg_3_ ( .D(n2983), .CK(clk), .Q(H1[3]) );
  DFFHQX1 H2_reg_4_ ( .D(n2694), .CK(clk), .Q(H2[4]) );
  DFFHQX1 H3_reg_4_ ( .D(n2725), .CK(clk), .Q(H3[4]) );
  DFFHQX1 H5_reg_3_ ( .D(n2790), .CK(clk), .Q(H5[3]) );
  DFFHQX1 B_reg_10_ ( .D(n2944), .CK(clk), .Q(SHA256_result[202]) );
  DFFHQX1 H_reg_14_ ( .D(n2588), .CK(clk), .Q(SHA256_result[14]) );
  DFFHQX1 F_reg_12_ ( .D(n2813), .CK(clk), .Q(SHA256_result[76]) );
  DFFHQX1 C_reg_9_ ( .D(n2912), .CK(clk), .Q(SHA256_result[169]) );
  DFFHQX1 G_reg_11_ ( .D(n2623), .CK(clk), .Q(SHA256_result[43]) );
  DFFHQXL D_reg_31_ ( .D(n2858), .CK(clk), .Q(SHA256_result[159]) );
  DFFHQXL B_reg_30_ ( .D(n2924), .CK(clk), .Q(SHA256_result[222]) );
  DFFHQXL C_reg_30_ ( .D(n2891), .CK(clk), .Q(SHA256_result[190]) );
  DFFHQXL H_reg_31_ ( .D(n2571), .CK(clk), .Q(SHA256_result[31]) );
  DFFHQX1 H3_reg_19_ ( .D(n2710), .CK(clk), .Q(H3[19]) );
  DFFHQX1 H6_reg_23_ ( .D(n2642), .CK(clk), .Q(H6[23]) );
  DFFHQX1 G_reg_31_ ( .D(n2603), .CK(clk), .Q(SHA256_result[63]) );
  DFFHQX1 F_reg_23_ ( .D(n2802), .CK(clk), .Q(SHA256_result[87]) );
  DFFHQX1 C_reg_19_ ( .D(n2902), .CK(clk), .Q(SHA256_result[179]) );
  DFFHQXL H0_reg_31_ ( .D(n3019), .CK(clk), .Q(H0[31]) );
  DFFHQXL H1_reg_30_ ( .D(n2956), .CK(clk), .Q(H1[30]) );
  DFFHQXL H5_reg_30_ ( .D(n2763), .CK(clk), .Q(H5[30]) );
  DFFHQXL H6_reg_30_ ( .D(n2635), .CK(clk), .Q(H6[30]) );
  DFFHQXL H2_reg_30_ ( .D(n2668), .CK(clk), .Q(H2[30]) );
  DFFHQXL H4_reg_31_ ( .D(n2730), .CK(clk), .Q(H4[31]) );
  DFFHQXL H7_reg_30_ ( .D(n2540), .CK(clk), .Q(H7[30]) );
  DFFHQXL H3_reg_30_ ( .D(n2699), .CK(clk), .Q(H3[30]) );
  DFFHQXL H2_reg_31_ ( .D(n2667), .CK(clk), .Q(H2[31]) );
  DFFHQXL H6_reg_31_ ( .D(n2634), .CK(clk), .Q(H6[31]) );
  DFFHQXL H7_reg_31_ ( .D(n2539), .CK(clk), .Q(H7[31]) );
  DFFHQXL H1_reg_31_ ( .D(n2955), .CK(clk), .Q(H1[31]) );
  DFFHQXL H5_reg_31_ ( .D(n2762), .CK(clk), .Q(H5[31]) );
  DFFHQXL H3_reg_31_ ( .D(n2698), .CK(clk), .Q(H3[31]) );
  DFFHQXL H0_reg_28_ ( .D(n3022), .CK(clk), .Q(H0[28]) );
  DFFHQXL H4_reg_28_ ( .D(n2733), .CK(clk), .Q(H4[28]) );
  DFFHQXL H0_reg_29_ ( .D(n3021), .CK(clk), .Q(H0[29]) );
  DFFHQXL H4_reg_29_ ( .D(n2732), .CK(clk), .Q(H4[29]) );
  DFFHQXL H0_reg_30_ ( .D(n3020), .CK(clk), .Q(H0[30]) );
  DFFHQXL H4_reg_30_ ( .D(n2731), .CK(clk), .Q(H4[30]) );
  DFFHQXL H3_reg_27_ ( .D(n2702), .CK(clk), .Q(H3[27]) );
  DFFHQXL H1_reg_27_ ( .D(n2959), .CK(clk), .Q(H1[27]) );
  DFFHQXL H1_reg_28_ ( .D(n2958), .CK(clk), .Q(H1[28]) );
  DFFHQXL H2_reg_28_ ( .D(n2670), .CK(clk), .Q(H2[28]) );
  DFFHQXL H3_reg_29_ ( .D(n2700), .CK(clk), .Q(H3[29]) );
  DFFHQXL H5_reg_27_ ( .D(n2766), .CK(clk), .Q(H5[27]) );
  DFFHQXL H5_reg_28_ ( .D(n2765), .CK(clk), .Q(H5[28]) );
  DFFHQXL H6_reg_28_ ( .D(n2637), .CK(clk), .Q(H6[28]) );
  DFFHQXL H7_reg_27_ ( .D(n2543), .CK(clk), .Q(H7[27]) );
  DFFHQXL H7_reg_28_ ( .D(n2542), .CK(clk), .Q(H7[28]) );
  DFFHQXL H3_reg_28_ ( .D(n2701), .CK(clk), .Q(H3[28]) );
  DFFHQXL H5_reg_29_ ( .D(n2764), .CK(clk), .Q(H5[29]) );
  DFFHQXL H6_reg_29_ ( .D(n2636), .CK(clk), .Q(H6[29]) );
  DFFHQXL H7_reg_29_ ( .D(n2541), .CK(clk), .Q(H7[29]) );
  DFFHQXL H1_reg_29_ ( .D(n2957), .CK(clk), .Q(H1[29]) );
  DFFHQXL H2_reg_27_ ( .D(n2671), .CK(clk), .Q(H2[27]) );
  DFFHQXL H2_reg_29_ ( .D(n2669), .CK(clk), .Q(H2[29]) );
  DFFHQXL H4_reg_21_ ( .D(n2740), .CK(clk), .Q(H4[21]) );
  DFFHQXL H0_reg_21_ ( .D(n3029), .CK(clk), .Q(H0[21]) );
  DFFHQXL H4_reg_23_ ( .D(n2738), .CK(clk), .Q(H4[23]) );
  DFFHQXL H0_reg_22_ ( .D(n3028), .CK(clk), .Q(H0[22]) );
  DFFHQXL H0_reg_23_ ( .D(n3027), .CK(clk), .Q(H0[23]) );
  DFFHQXL H4_reg_26_ ( .D(n2735), .CK(clk), .Q(H4[26]) );
  DFFHQXL H4_reg_27_ ( .D(n2734), .CK(clk), .Q(H4[27]) );
  DFFHQXL H0_reg_27_ ( .D(n3023), .CK(clk), .Q(H0[27]) );
  DFFHQXL H0_reg_20_ ( .D(n3030), .CK(clk), .Q(H0[20]) );
  DFFHQXL H4_reg_20_ ( .D(n2741), .CK(clk), .Q(H4[20]) );
  DFFHQXL D_reg_30_ ( .D(n2859), .CK(clk), .Q(SHA256_result[158]) );
  DFFHQXL H4_reg_22_ ( .D(n2739), .CK(clk), .Q(H4[22]) );
  DFFHQXL H0_reg_26_ ( .D(n3024), .CK(clk), .Q(H0[26]) );
  DFFHQXL H0_reg_25_ ( .D(n3025), .CK(clk), .Q(H0[25]) );
  DFFHQXL H0_reg_24_ ( .D(n3026), .CK(clk), .Q(H0[24]) );
  DFFHQXL H4_reg_25_ ( .D(n2736), .CK(clk), .Q(H4[25]) );
  DFFHQXL H4_reg_24_ ( .D(n2737), .CK(clk), .Q(H4[24]) );
  DFFHQXL H2_reg_24_ ( .D(n2674), .CK(clk), .Q(H2[24]) );
  DFFHQXL H5_reg_26_ ( .D(n2767), .CK(clk), .Q(H5[26]) );
  DFFHQXL H1_reg_25_ ( .D(n2961), .CK(clk), .Q(H1[25]) );
  DFFHQXL H2_reg_26_ ( .D(n2672), .CK(clk), .Q(H2[26]) );
  DFFHQXL H3_reg_24_ ( .D(n2705), .CK(clk), .Q(H3[24]) );
  DFFHQXL H3_reg_26_ ( .D(n2703), .CK(clk), .Q(H3[26]) );
  DFFHQXL H5_reg_24_ ( .D(n2769), .CK(clk), .Q(H5[24]) );
  DFFHQXL H6_reg_26_ ( .D(n2639), .CK(clk), .Q(H6[26]) );
  DFFHQXL H7_reg_25_ ( .D(n2545), .CK(clk), .Q(H7[25]) );
  DFFHQXL H6_reg_24_ ( .D(n2641), .CK(clk), .Q(H6[24]) );
  DFFHQXL H1_reg_26_ ( .D(n2960), .CK(clk), .Q(H1[26]) );
  DFFHQXL H2_reg_25_ ( .D(n2673), .CK(clk), .Q(H2[25]) );
  DFFHQXL H7_reg_26_ ( .D(n2544), .CK(clk), .Q(H7[26]) );
  DFFHQXL H7_reg_24_ ( .D(n2546), .CK(clk), .Q(H7[24]) );
  DFFHQXL H6_reg_25_ ( .D(n2640), .CK(clk), .Q(H6[25]) );
  DFFHQXL H4_reg_15_ ( .D(n2746), .CK(clk), .Q(H4[15]) );
  DFFHQXL H0_reg_18_ ( .D(n3032), .CK(clk), .Q(H0[18]) );
  DFFHQXL H0_reg_11_ ( .D(n3039), .CK(clk), .Q(H0[11]) );
  DFFHQXL H0_reg_17_ ( .D(n3033), .CK(clk), .Q(H0[17]) );
  DFFHQXL H0_reg_12_ ( .D(n3038), .CK(clk), .Q(H0[12]) );
  DFFHQXL H0_reg_15_ ( .D(n3035), .CK(clk), .Q(H0[15]) );
  DFFHQXL H0_reg_19_ ( .D(n3031), .CK(clk), .Q(H0[19]) );
  DFFHQXL H4_reg_13_ ( .D(n2748), .CK(clk), .Q(H4[13]) );
  DFFHQXL H4_reg_16_ ( .D(n2745), .CK(clk), .Q(H4[16]) );
  DFFHQXL H0_reg_14_ ( .D(n3036), .CK(clk), .Q(H0[14]) );
  DFFHQXL H4_reg_17_ ( .D(n2744), .CK(clk), .Q(H4[17]) );
  DFFHQXL H4_reg_19_ ( .D(n2742), .CK(clk), .Q(H4[19]) );
  DFFHQXL H4_reg_12_ ( .D(n2749), .CK(clk), .Q(H4[12]) );
  DFFHQXL H4_reg_11_ ( .D(n2750), .CK(clk), .Q(H4[11]) );
  DFFHQXL H4_reg_14_ ( .D(n2747), .CK(clk), .Q(H4[14]) );
  DFFHQXL H4_reg_18_ ( .D(n2743), .CK(clk), .Q(H4[18]) );
  DFFHQXL H0_reg_13_ ( .D(n3037), .CK(clk), .Q(H0[13]) );
  DFFHQXL H0_reg_10_ ( .D(n3040), .CK(clk), .Q(H0[10]) );
  DFFHQXL H4_reg_10_ ( .D(n2751), .CK(clk), .Q(H4[10]) );
  DFFHQXL H0_reg_16_ ( .D(n3034), .CK(clk), .Q(H0[16]) );
  DFFHQXL D_reg_29_ ( .D(n2860), .CK(clk), .Q(SHA256_result[157]) );
  DFFHQXL D_reg_28_ ( .D(n2861), .CK(clk), .Q(SHA256_result[156]) );
  DFFHQXL H5_reg_23_ ( .D(n2770), .CK(clk), .Q(H5[23]) );
  DFFHQXL H5_reg_22_ ( .D(n2771), .CK(clk), .Q(H5[22]) );
  DFFHQXL H1_reg_24_ ( .D(n2962), .CK(clk), .Q(H1[24]) );
  DFFHQXL H2_reg_22_ ( .D(n2676), .CK(clk), .Q(H2[22]) );
  DFFHQXL H3_reg_22_ ( .D(n2707), .CK(clk), .Q(H3[22]) );
  DFFHQXL H1_reg_22_ ( .D(n2964), .CK(clk), .Q(H1[22]) );
  DFFHQXL H1_reg_23_ ( .D(n2963), .CK(clk), .Q(H1[23]) );
  DFFHQXL H3_reg_23_ ( .D(n2706), .CK(clk), .Q(H3[23]) );
  DFFHQXL H0_reg_8_ ( .D(n3042), .CK(clk), .Q(H0[8]) );
  DFFHQXL H0_reg_4_ ( .D(n3046), .CK(clk), .Q(H0[4]) );
  DFFHQXL H0_reg_3_ ( .D(n3047), .CK(clk), .Q(H0[3]) );
  DFFHQXL H4_reg_8_ ( .D(n2753), .CK(clk), .Q(H4[8]) );
  DFFHQXL H0_reg_6_ ( .D(n3044), .CK(clk), .Q(H0[6]) );
  DFFHQXL H0_reg_7_ ( .D(n3043), .CK(clk), .Q(H0[7]) );
  DFFHQXL H0_reg_2_ ( .D(n3048), .CK(clk), .Q(H0[2]) );
  DFFHQXL H0_reg_9_ ( .D(n3041), .CK(clk), .Q(H0[9]) );
  DFFHQXL D_reg_25_ ( .D(n2864), .CK(clk), .Q(SHA256_result[153]) );
  DFFHQXL D_reg_24_ ( .D(n2865), .CK(clk), .Q(SHA256_result[152]) );
  DFFHQXL D_reg_26_ ( .D(n2863), .CK(clk), .Q(SHA256_result[154]) );
  DFFHQXL D_reg_27_ ( .D(n2862), .CK(clk), .Q(SHA256_result[155]) );
  DFFHQXL H1_reg_20_ ( .D(n2966), .CK(clk), .Q(H1[20]) );
  DFFHQXL H5_reg_20_ ( .D(n2773), .CK(clk), .Q(H5[20]) );
  DFFHQXL H6_reg_20_ ( .D(n2645), .CK(clk), .Q(H6[20]) );
  DFFHQXL H7_reg_20_ ( .D(n2550), .CK(clk), .Q(H7[20]) );
  DFFHQXL H3_reg_20_ ( .D(n2709), .CK(clk), .Q(H3[20]) );
  DFFHQXL H6_reg_22_ ( .D(n2643), .CK(clk), .Q(H6[22]) );
  DFFHQXL H2_reg_21_ ( .D(n2677), .CK(clk), .Q(H2[21]) );
  DFFHQXL H7_reg_22_ ( .D(n2548), .CK(clk), .Q(H7[22]) );
  DFFHQXL H2_reg_19_ ( .D(n2679), .CK(clk), .Q(H2[19]) );
  DFFHQXL H1_reg_19_ ( .D(n2967), .CK(clk), .Q(H1[19]) );
  DFFHQXL H2_reg_20_ ( .D(n2678), .CK(clk), .Q(H2[20]) );
  DFFHQXL H3_reg_21_ ( .D(n2708), .CK(clk), .Q(H3[21]) );
  DFFHQXL H5_reg_19_ ( .D(n2774), .CK(clk), .Q(H5[19]) );
  DFFHQXL H5_reg_21_ ( .D(n2772), .CK(clk), .Q(H5[21]) );
  DFFHQXL H6_reg_21_ ( .D(n2644), .CK(clk), .Q(H6[21]) );
  DFFHQXL H7_reg_21_ ( .D(n2549), .CK(clk), .Q(H7[21]) );
  DFFHQXL H0_reg_0_ ( .D(n3050), .CK(clk), .Q(H0[0]) );
  DFFHQXL H4_reg_4_ ( .D(n2757), .CK(clk), .Q(H4[4]) );
  DFFHQXL H4_reg_0_ ( .D(n2761), .CK(clk), .Q(H4[0]) );
  DFFHQXL H4_reg_1_ ( .D(n2760), .CK(clk), .Q(H4[1]) );
  DFFHQXL H4_reg_3_ ( .D(n2758), .CK(clk), .Q(H4[3]) );
  DFFHQXL H4_reg_7_ ( .D(n2754), .CK(clk), .Q(H4[7]) );
  DFFHQXL H4_reg_2_ ( .D(n2759), .CK(clk), .Q(H4[2]) );
  DFFHQXL H4_reg_5_ ( .D(n2756), .CK(clk), .Q(H4[5]) );
  DFFHQXL H_reg_30_ ( .D(n2572), .CK(clk), .Q(SHA256_result[30]) );
  DFFHQXL D_reg_23_ ( .D(n2866), .CK(clk), .Q(SHA256_result[151]) );
  DFFHQXL C_reg_29_ ( .D(n2892), .CK(clk), .Q(SHA256_result[189]) );
  DFFHQXL D_reg_18_ ( .D(n2871), .CK(clk), .Q(SHA256_result[146]) );
  DFFHQXL D_reg_19_ ( .D(n2870), .CK(clk), .Q(SHA256_result[147]) );
  DFFHQXL D_reg_16_ ( .D(n2873), .CK(clk), .Q(SHA256_result[144]) );
  DFFHQXL B_reg_29_ ( .D(n2925), .CK(clk), .Q(SHA256_result[221]) );
  DFFHQXL D_reg_22_ ( .D(n2867), .CK(clk), .Q(SHA256_result[150]) );
  DFFHQXL B_reg_28_ ( .D(n2926), .CK(clk), .Q(SHA256_result[220]) );
  DFFHQXL C_reg_28_ ( .D(n2893), .CK(clk), .Q(SHA256_result[188]) );
  DFFHQXL D_reg_21_ ( .D(n2868), .CK(clk), .Q(SHA256_result[149]) );
  DFFHQXL D_reg_20_ ( .D(n2869), .CK(clk), .Q(SHA256_result[148]) );
  DFFHQXL H6_reg_18_ ( .D(n2647), .CK(clk), .Q(H6[18]) );
  DFFHQXL H7_reg_17_ ( .D(n2553), .CK(clk), .Q(H7[17]) );
  DFFHQXL H7_reg_18_ ( .D(n2552), .CK(clk), .Q(H7[18]) );
  DFFHQXL H1_reg_18_ ( .D(n2968), .CK(clk), .Q(H1[18]) );
  DFFHQXL H6_reg_17_ ( .D(n2648), .CK(clk), .Q(H6[17]) );
  DFFHQXL H2_reg_17_ ( .D(n2681), .CK(clk), .Q(H2[17]) );
  DFFHQXL H5_reg_18_ ( .D(n2775), .CK(clk), .Q(H5[18]) );
  DFFHQXL H3_reg_18_ ( .D(n2711), .CK(clk), .Q(H3[18]) );
  DFFHQXL H5_reg_17_ ( .D(n2776), .CK(clk), .Q(H5[17]) );
  DFFHQXL H_reg_28_ ( .D(n2574), .CK(clk), .Q(SHA256_result[28]) );
  DFFHQXL H_reg_29_ ( .D(n2573), .CK(clk), .Q(SHA256_result[29]) );
  DFFHQXL D_reg_17_ ( .D(n2872), .CK(clk), .Q(SHA256_result[145]) );
  DFFHQXL G_reg_28_ ( .D(n2606), .CK(clk), .Q(SHA256_result[60]) );
  DFFHQXL G_reg_30_ ( .D(n2604), .CK(clk), .Q(SHA256_result[62]) );
  DFFHQXL C_reg_26_ ( .D(n2895), .CK(clk), .Q(SHA256_result[186]) );
  DFFHQXL C_reg_24_ ( .D(n2897), .CK(clk), .Q(SHA256_result[184]) );
  DFFHQXL D_reg_14_ ( .D(n2875), .CK(clk), .Q(SHA256_result[142]) );
  DFFHQXL D_reg_12_ ( .D(n2877), .CK(clk), .Q(SHA256_result[140]) );
  DFFHQXL D_reg_10_ ( .D(n2879), .CK(clk), .Q(SHA256_result[138]) );
  DFFHQXL D_reg_11_ ( .D(n2878), .CK(clk), .Q(SHA256_result[139]) );
  DFFHQXL D_reg_13_ ( .D(n2876), .CK(clk), .Q(SHA256_result[141]) );
  DFFHQXL B_reg_27_ ( .D(n2927), .CK(clk), .Q(SHA256_result[219]) );
  DFFHQXL B_reg_26_ ( .D(n2928), .CK(clk), .Q(SHA256_result[218]) );
  DFFHQXL D_reg_15_ ( .D(n2874), .CK(clk), .Q(SHA256_result[143]) );
  DFFHQXL F_reg_29_ ( .D(n2796), .CK(clk), .Q(SHA256_result[93]) );
  DFFHQXL G_reg_29_ ( .D(n2605), .CK(clk), .Q(SHA256_result[61]) );
  DFFHQXL F_reg_30_ ( .D(n2795), .CK(clk), .Q(SHA256_result[94]) );
  DFFHQXL C_reg_27_ ( .D(n2894), .CK(clk), .Q(SHA256_result[187]) );
  DFFHQXL B_reg_24_ ( .D(n2930), .CK(clk), .Q(SHA256_result[216]) );
  DFFHQXL H7_reg_16_ ( .D(n2554), .CK(clk), .Q(H7[16]) );
  DFFHQXL H1_reg_15_ ( .D(n2971), .CK(clk), .Q(H1[15]) );
  DFFHQXL H1_reg_16_ ( .D(n2970), .CK(clk), .Q(H1[16]) );
  DFFHQXL H5_reg_14_ ( .D(n2779), .CK(clk), .Q(H5[14]) );
  DFFHQXL H5_reg_16_ ( .D(n2777), .CK(clk), .Q(H5[16]) );
  DFFHQXL H6_reg_15_ ( .D(n2650), .CK(clk), .Q(H6[15]) );
  DFFHQXL H6_reg_16_ ( .D(n2649), .CK(clk), .Q(H6[16]) );
  DFFHQXL H7_reg_15_ ( .D(n2555), .CK(clk), .Q(H7[15]) );
  DFFHQXL H2_reg_15_ ( .D(n2683), .CK(clk), .Q(H2[15]) );
  DFFHQXL H3_reg_16_ ( .D(n2713), .CK(clk), .Q(H3[16]) );
  DFFHQXL H1_reg_14_ ( .D(n2972), .CK(clk), .Q(H1[14]) );
  DFFHQXL H2_reg_16_ ( .D(n2682), .CK(clk), .Q(H2[16]) );
  DFFHQXL H5_reg_15_ ( .D(n2778), .CK(clk), .Q(H5[15]) );
  DFFHQXL D_reg_3_ ( .D(n2886), .CK(clk), .Q(SHA256_result[131]) );
  DFFHQXL D_reg_4_ ( .D(n2885), .CK(clk), .Q(SHA256_result[132]) );
  DFFHQXL H_reg_24_ ( .D(n2578), .CK(clk), .Q(SHA256_result[24]) );
  DFFHQXL H_reg_25_ ( .D(n2577), .CK(clk), .Q(SHA256_result[25]) );
  DFFHQXL H_reg_26_ ( .D(n2576), .CK(clk), .Q(SHA256_result[26]) );
  DFFHQXL H_reg_27_ ( .D(n2575), .CK(clk), .Q(SHA256_result[27]) );
  DFFHQXL D_reg_9_ ( .D(n2880), .CK(clk), .Q(SHA256_result[137]) );
  DFFHQXL D_reg_7_ ( .D(n2882), .CK(clk), .Q(SHA256_result[135]) );
  DFFHQXL D_reg_6_ ( .D(n2883), .CK(clk), .Q(SHA256_result[134]) );
  DFFHQXL C_reg_22_ ( .D(n2899), .CK(clk), .Q(SHA256_result[182]) );
  DFFHQXL D_reg_8_ ( .D(n2881), .CK(clk), .Q(SHA256_result[136]) );
  DFFHQXL G_reg_27_ ( .D(n2607), .CK(clk), .Q(SHA256_result[59]) );
  DFFHQXL D_reg_5_ ( .D(n2884), .CK(clk), .Q(SHA256_result[133]) );
  DFFHQXL B_reg_21_ ( .D(n2933), .CK(clk), .Q(SHA256_result[213]) );
  DFFHQXL B_reg_22_ ( .D(n2932), .CK(clk), .Q(SHA256_result[214]) );
  DFFHQXL C_reg_21_ ( .D(n2900), .CK(clk), .Q(SHA256_result[181]) );
  DFFHQXL C_reg_23_ ( .D(n2898), .CK(clk), .Q(SHA256_result[183]) );
  DFFHQXL C_reg_20_ ( .D(n2901), .CK(clk), .Q(SHA256_result[180]) );
  DFFHQXL F_reg_28_ ( .D(n2797), .CK(clk), .Q(SHA256_result[92]) );
  DFFHQXL B_reg_20_ ( .D(n2934), .CK(clk), .Q(SHA256_result[212]) );
  DFFHQXL B_reg_25_ ( .D(n2929), .CK(clk), .Q(SHA256_result[217]) );
  DFFHQXL H5_reg_12_ ( .D(n2781), .CK(clk), .Q(H5[12]) );
  DFFHQXL H6_reg_13_ ( .D(n2652), .CK(clk), .Q(H6[13]) );
  DFFHQXL H7_reg_12_ ( .D(n2558), .CK(clk), .Q(H7[12]) );
  DFFHQXL H7_reg_13_ ( .D(n2557), .CK(clk), .Q(H7[13]) );
  DFFHQXL H5_reg_11_ ( .D(n2782), .CK(clk), .Q(H5[11]) );
  DFFHQXL H1_reg_11_ ( .D(n2975), .CK(clk), .Q(H1[11]) );
  DFFHQXL H1_reg_13_ ( .D(n2973), .CK(clk), .Q(H1[13]) );
  DFFHQXL H6_reg_12_ ( .D(n2653), .CK(clk), .Q(H6[12]) );
  DFFHQXL H6_reg_14_ ( .D(n2651), .CK(clk), .Q(H6[14]) );
  DFFHQXL H2_reg_13_ ( .D(n2685), .CK(clk), .Q(H2[13]) );
  DFFHQXL H2_reg_14_ ( .D(n2684), .CK(clk), .Q(H2[14]) );
  DFFHQXL H3_reg_14_ ( .D(n2715), .CK(clk), .Q(H3[14]) );
  DFFHQXL H2_reg_12_ ( .D(n2686), .CK(clk), .Q(H2[12]) );
  DFFHQXL H3_reg_12_ ( .D(n2717), .CK(clk), .Q(H3[12]) );
  DFFHQXL H1_reg_12_ ( .D(n2974), .CK(clk), .Q(H1[12]) );
  DFFHQXL H5_reg_13_ ( .D(n2780), .CK(clk), .Q(H5[13]) );
  DFFHQXL D_reg_2_ ( .D(n2887), .CK(clk), .Q(SHA256_result[130]) );
  DFFHQXL H_reg_20_ ( .D(n2582), .CK(clk), .Q(SHA256_result[20]) );
  DFFHQXL C_reg_18_ ( .D(n2903), .CK(clk), .Q(SHA256_result[178]) );
  DFFHQXL H_reg_22_ ( .D(n2580), .CK(clk), .Q(SHA256_result[22]) );
  DFFHQXL G_reg_24_ ( .D(n2610), .CK(clk), .Q(SHA256_result[56]) );
  DFFHQXL F_reg_26_ ( .D(n2799), .CK(clk), .Q(SHA256_result[90]) );
  DFFHQXL F_reg_24_ ( .D(n2801), .CK(clk), .Q(SHA256_result[88]) );
  DFFHQXL G_reg_25_ ( .D(n2609), .CK(clk), .Q(SHA256_result[57]) );
  DFFHQXL B_reg_19_ ( .D(n2935), .CK(clk), .Q(SHA256_result[211]) );
  DFFHQXL F_reg_25_ ( .D(n2800), .CK(clk), .Q(SHA256_result[89]) );
  DFFHQXL G_reg_26_ ( .D(n2608), .CK(clk), .Q(SHA256_result[58]) );
  DFFHQXL H4_reg_6_ ( .D(n2755), .CK(clk), .Q(H4[6]) );
  DFFHQXL H4_reg_9_ ( .D(n2752), .CK(clk), .Q(H4[9]) );
  DFFHQXL H0_reg_5_ ( .D(n3045), .CK(clk), .Q(H0[5]) );
  DFFHQXL H0_reg_1_ ( .D(n3049), .CK(clk), .Q(H0[1]) );
  DFFHQX1 H6_reg_6_ ( .D(n2659), .CK(clk), .Q(H6[6]) );
  DFFHQX1 H7_reg_5_ ( .D(n2565), .CK(clk), .Q(H7[5]) );
  DFFHQX1 H_reg_12_ ( .D(n2590), .CK(clk), .Q(SHA256_result[12]) );
  DFFHQX1 H_reg_4_ ( .D(n2598), .CK(clk), .Q(SHA256_result[4]) );
  DFFHQX1 B_reg_7_ ( .D(n2947), .CK(clk), .Q(SHA256_result[199]) );
  DFFX4 F_reg_1_ ( .D(n2824), .CK(clk), .Q(n115), .QN(n116) );
  DFFHQXL C_reg_31_ ( .D(n2890), .CK(clk), .Q(SHA256_result[191]) );
  DFFHQX4 H7_reg_0_ ( .D(n2570), .CK(clk), .Q(H7[0]) );
  DFFHQX1 H7_reg_23_ ( .D(n2547), .CK(clk), .Q(H7[23]) );
  DFFHQX1 H7_reg_3_ ( .D(n2567), .CK(clk), .Q(H7[3]) );
  DFFHQX1 H2_reg_18_ ( .D(n2680), .CK(clk), .Q(H2[18]) );
  DFFHQX1 G_reg_23_ ( .D(n2611), .CK(clk), .Q(SHA256_result[55]) );
  DFFHQX1 B_reg_18_ ( .D(n2936), .CK(clk), .Q(SHA256_result[210]) );
  DFFHQXL H3_reg_13_ ( .D(n2716), .CK(clk), .Q(H3[13]) );
  DFFHQXL C_reg_16_ ( .D(n2905), .CK(clk), .Q(SHA256_result[176]) );
  DFFHQXL G_reg_22_ ( .D(n2612), .CK(clk), .Q(SHA256_result[54]) );
  DFFHQXL B_reg_15_ ( .D(n2939), .CK(clk), .Q(SHA256_result[207]) );
  DFFHQXL B_reg_17_ ( .D(n2937), .CK(clk), .Q(SHA256_result[209]) );
  DFFHQXL F_reg_22_ ( .D(n2803), .CK(clk), .Q(SHA256_result[86]) );
  DFFHQXL B_reg_16_ ( .D(n2938), .CK(clk), .Q(SHA256_result[208]) );
  DFFHQX1 H_reg_2_ ( .D(n2600), .CK(clk), .Q(SHA256_result[2]) );
  DFFHQX1 C_reg_14_ ( .D(n2907), .CK(clk), .Q(SHA256_result[174]) );
  DFFHQXL H6_reg_11_ ( .D(n2654), .CK(clk), .Q(H6[11]) );
  DFFHQX1 H_reg_1_ ( .D(n2601), .CK(clk), .Q(SHA256_result[1]) );
  DFFX4 H6_reg_0_ ( .D(n2665), .CK(clk), .Q(n114) );
  DFFHQX1 H3_reg_17_ ( .D(n2712), .CK(clk), .Q(H3[17]) );
  DFFHQX1 C_reg_17_ ( .D(n2904), .CK(clk), .Q(SHA256_result[177]) );
  DFFHQXL H7_reg_11_ ( .D(n2559), .CK(clk), .Q(H7[11]) );
  DFFX4 H3_reg_0_ ( .D(n2729), .CK(clk), .Q(n112) );
  DFFX4 H6_reg_1_ ( .D(n2664), .CK(clk), .Q(n110) );
  DFFHQX4 B_reg_1_ ( .D(n2953), .CK(clk), .Q(SHA256_result[193]) );
  DFFHQX1 H6_reg_27_ ( .D(n2638), .CK(clk), .Q(H6[27]) );
  DFFHQX1 F_reg_27_ ( .D(n2798), .CK(clk), .Q(SHA256_result[91]) );
  DFFX4 F_reg_0_ ( .D(n2825), .CK(clk), .Q(n107), .QN(n106) );
  DFFHQX1 H3_reg_15_ ( .D(n2714), .CK(clk), .Q(H3[15]) );
  DFFHQX4 H3_reg_1_ ( .D(n2728), .CK(clk), .Q(H3[1]) );
  DFFHQXL F_reg_31_ ( .D(n2794), .CK(clk), .Q(SHA256_result[95]) );
  DFFHQXL B_reg_31_ ( .D(n2923), .CK(clk), .Q(SHA256_result[223]) );
  DFFX4 A_reg_1_ ( .D(n3017), .CK(clk), .Q(n101), .QN(n102) );
  DFFHQX1 H5_reg_25_ ( .D(n2768), .CK(clk), .Q(H5[25]) );
  DFFTRX1 round_reg_5_ ( .D(N182), .RN(n141), .CK(clk), .Q(round[5]), .QN(
        n1371) );
  DFFHQX1 H5_reg_8_ ( .D(n2785), .CK(clk), .Q(H5[8]) );
  DFFHQX1 H5_reg_9_ ( .D(n2784), .CK(clk), .Q(H5[9]) );
  DFFHQX1 H6_reg_9_ ( .D(n2656), .CK(clk), .Q(H6[9]) );
  DFFHQX1 H6_reg_10_ ( .D(n2655), .CK(clk), .Q(H6[10]) );
  DFFHQX1 H7_reg_9_ ( .D(n2561), .CK(clk), .Q(H7[9]) );
  DFFHQX1 H1_reg_9_ ( .D(n2977), .CK(clk), .Q(H1[9]) );
  DFFHQX1 H2_reg_8_ ( .D(n2690), .CK(clk), .Q(H2[8]) );
  DFFHQX1 H2_reg_9_ ( .D(n2689), .CK(clk), .Q(H2[9]) );
  DFFHQX1 H3_reg_8_ ( .D(n2721), .CK(clk), .Q(H3[8]) );
  DFFHQX1 H6_reg_8_ ( .D(n2657), .CK(clk), .Q(H6[8]) );
  DFFHQX1 H7_reg_8_ ( .D(n2562), .CK(clk), .Q(H7[8]) );
  DFFHQX1 H7_reg_10_ ( .D(n2560), .CK(clk), .Q(H7[10]) );
  DFFHQX1 G_reg_18_ ( .D(n2616), .CK(clk), .Q(SHA256_result[50]) );
  DFFHQX1 E_reg_24_ ( .D(n2833), .CK(clk), .Q(SHA256_result[120]) );
  DFFHQX1 H1_reg_5_ ( .D(n2981), .CK(clk), .Q(H1[5]) );
  DFFHQX1 H3_reg_6_ ( .D(n2723), .CK(clk), .Q(H3[6]) );
  DFFHQX1 H7_reg_6_ ( .D(n2564), .CK(clk), .Q(H7[6]) );
  DFFHQX1 H7_reg_7_ ( .D(n2563), .CK(clk), .Q(H7[7]) );
  DFFHQX1 H1_reg_7_ ( .D(n2979), .CK(clk), .Q(H1[7]) );
  DFFHQX1 H5_reg_7_ ( .D(n2786), .CK(clk), .Q(H5[7]) );
  DFFHQX1 H6_reg_7_ ( .D(n2658), .CK(clk), .Q(H6[7]) );
  DFFHQX1 H_reg_6_ ( .D(n2596), .CK(clk), .Q(SHA256_result[6]) );
  DFFHQX1 H_reg_9_ ( .D(n2593), .CK(clk), .Q(SHA256_result[9]) );
  DFFHQX1 H_reg_13_ ( .D(n2589), .CK(clk), .Q(SHA256_result[13]) );
  DFFHQX1 F_reg_7_ ( .D(n2818), .CK(clk), .Q(SHA256_result[71]) );
  DFFHQX1 C_reg_15_ ( .D(n2906), .CK(clk), .Q(SHA256_result[175]) );
  DFFHQX1 E_reg_6_ ( .D(n2851), .CK(clk), .Q(SHA256_result[102]) );
  DFFHQX1 E_reg_12_ ( .D(n2845), .CK(clk), .Q(SHA256_result[108]) );
  DFFHQX1 E_reg_8_ ( .D(n2849), .CK(clk), .Q(SHA256_result[104]) );
  DFFHQX1 E_reg_9_ ( .D(n2848), .CK(clk), .Q(SHA256_result[105]) );
  DFFHQX1 H_reg_8_ ( .D(n2594), .CK(clk), .Q(SHA256_result[8]) );
  DFFHQX1 H_reg_10_ ( .D(n2592), .CK(clk), .Q(SHA256_result[10]) );
  DFFHQX1 C_reg_6_ ( .D(n2915), .CK(clk), .Q(SHA256_result[166]) );
  DFFHQX1 F_reg_13_ ( .D(n2812), .CK(clk), .Q(SHA256_result[77]) );
  DFFHQX1 G_reg_12_ ( .D(n2622), .CK(clk), .Q(SHA256_result[44]) );
  DFFHQX1 E_reg_22_ ( .D(n2835), .CK(clk), .Q(SHA256_result[118]) );
  DFFX4 G_reg_0_ ( .D(n2666), .CK(clk), .Q(n95), .QN(n94) );
  DFFHQX4 H5_reg_0_ ( .D(n2793), .CK(clk), .Q(H5[0]) );
  DFFHQX4 H2_reg_0_ ( .D(n2922), .CK(clk), .Q(H2[0]) );
  DFFX4 C_reg_0_ ( .D(n2921), .CK(clk), .Q(n89), .QN(n88) );
  DFFX4 C_reg_1_ ( .D(n2920), .CK(clk), .Q(n86), .QN(n85) );
  DFFHQX2 H2_reg_1_ ( .D(n2697), .CK(clk), .Q(H2[1]) );
  DFFHQX4 H5_reg_1_ ( .D(n2792), .CK(clk), .Q(H5[1]) );
  DFFHQX2 G_reg_13_ ( .D(n2621), .CK(clk), .Q(SHA256_result[45]) );
  DFFHQXL E_reg_27_ ( .D(n2830), .CK(clk), .Q(SHA256_result[123]) );
  DFFHQX4 A_reg_28_ ( .D(n2990), .CK(clk), .Q(SHA256_result[252]) );
  DFFHQX4 E_reg_31_ ( .D(n2826), .CK(clk), .Q(SHA256_result[127]) );
  DFFHQX4 E_reg_29_ ( .D(n2828), .CK(clk), .Q(SHA256_result[125]) );
  DFFHQXL A_reg_7_ ( .D(n3011), .CK(clk), .Q(SHA256_result[231]) );
  DFFHQX2 G_reg_10_ ( .D(n2624), .CK(clk), .Q(SHA256_result[42]) );
  DFFHQX4 A_reg_31_ ( .D(n2987), .CK(clk), .Q(SHA256_result[255]) );
  DFFTRX1 round_reg_4_ ( .D(N181), .RN(n141), .CK(clk), .Q(n334), .QN(n332) );
  DFFTRX1 round_reg_1_ ( .D(N178), .RN(n141), .CK(clk), .Q(n331), .QN(n336) );
  DFFTRX2 round_reg_3_ ( .D(N180), .RN(n141), .CK(clk), .Q(round[3]), .QN(
        n1384) );
  DFFTRX2 round_reg_2_ ( .D(N179), .RN(n141), .CK(clk), .Q(round[2]), .QN(
        n1389) );
  DFFHQX2 B_reg_2_ ( .D(n2952), .CK(clk), .Q(SHA256_result[194]) );
  DFFTRX2 round_reg_0_ ( .D(N177), .RN(n141), .CK(clk), .Q(round[0]), .QN(
        n1397) );
  DFFHQX2 F_reg_8_ ( .D(n2817), .CK(clk), .Q(SHA256_result[72]) );
  DFFHQX2 E_reg_16_ ( .D(n2841), .CK(clk), .Q(SHA256_result[112]) );
  DFFHQX2 E_reg_26_ ( .D(n2831), .CK(clk), .Q(SHA256_result[122]) );
  DFFHQX2 E_reg_28_ ( .D(n2829), .CK(clk), .Q(SHA256_result[124]) );
  DFFHQX2 F_reg_5_ ( .D(n2820), .CK(clk), .Q(SHA256_result[69]) );
  DFFHQX2 G_reg_5_ ( .D(n2629), .CK(clk), .Q(SHA256_result[37]) );
  DFFHQX2 Kt_reg_15_ ( .D(N3017), .CK(clk), .Q(Kt[15]) );
  DFFHQX2 Kt_reg_14_ ( .D(N3016), .CK(clk), .Q(Kt[14]) );
  DFFHQX2 Kt_reg_12_ ( .D(N3014), .CK(clk), .Q(Kt[12]) );
  DFFHQX2 Kt_reg_11_ ( .D(N3013), .CK(clk), .Q(Kt[11]) );
  DFFHQX2 Kt_reg_10_ ( .D(N3012), .CK(clk), .Q(Kt[10]) );
  DFFHQX2 Kt_reg_9_ ( .D(N3011), .CK(clk), .Q(Kt[9]) );
  DFFHQX2 Kt_reg_7_ ( .D(N3009), .CK(clk), .Q(Kt[7]) );
  DFFHQX2 Kt_reg_6_ ( .D(N3008), .CK(clk), .Q(Kt[6]) );
  DFFHQX2 Kt_reg_5_ ( .D(N3007), .CK(clk), .Q(Kt[5]) );
  DFFHQX2 Kt_reg_4_ ( .D(N3006), .CK(clk), .Q(Kt[4]) );
  DFFHQX1 H_reg_0_ ( .D(n2602), .CK(clk), .Q(SHA256_result[0]) );
  DFFHQX1 H6_reg_19_ ( .D(n2646), .CK(clk), .Q(H6[19]) );
  DFFHQX1 F_reg_19_ ( .D(n2806), .CK(clk), .Q(SHA256_result[83]) );
  DFFX2 H1_reg_0_ ( .D(n2986), .CK(clk), .Q(n91) );
  DFFHQX1 H1_reg_17_ ( .D(n2969), .CK(clk), .Q(H1[17]) );
  DFFHQX1 H6_reg_3_ ( .D(n2662), .CK(clk), .Q(H6[3]) );
  DFFHQX1 H5_reg_2_ ( .D(n2791), .CK(clk), .Q(H5[2]) );
  DFFHQX1 H7_reg_19_ ( .D(n2551), .CK(clk), .Q(H7[19]) );
  DFFHQX1 G_reg_19_ ( .D(n2615), .CK(clk), .Q(SHA256_result[51]) );
  DFFHQX1 H1_reg_10_ ( .D(n2976), .CK(clk), .Q(H1[10]) );
  DFFHQX2 F_reg_10_ ( .D(n2815), .CK(clk), .Q(SHA256_result[74]) );
  DFFHQX2 F_reg_9_ ( .D(n2816), .CK(clk), .Q(SHA256_result[73]) );
  DFFHQX2 G_reg_9_ ( .D(n2625), .CK(clk), .Q(SHA256_result[41]) );
  DFFHQX1 H1_reg_2_ ( .D(n2984), .CK(clk), .Q(H1[2]) );
  DFFHQX1 A_reg_2_ ( .D(n3016), .CK(clk), .Q(SHA256_result[226]) );
  DFFHQX1 G_reg_7_ ( .D(n2627), .CK(clk), .Q(SHA256_result[39]) );
  DFFHQX1 H3_reg_25_ ( .D(n2704), .CK(clk), .Q(H3[25]) );
  DFFHQX1 C_reg_25_ ( .D(n2896), .CK(clk), .Q(SHA256_result[185]) );
  DFFHQX1 H1_reg_4_ ( .D(n2982), .CK(clk), .Q(H1[4]) );
  DFFHQX1 H1_reg_21_ ( .D(n2965), .CK(clk), .Q(H1[21]) );
  DFFHQX1 H2_reg_23_ ( .D(n2675), .CK(clk), .Q(H2[23]) );
  DFFHQX1 B_reg_23_ ( .D(n2931), .CK(clk), .Q(SHA256_result[215]) );
  DFFHQX1 H7_reg_14_ ( .D(n2556), .CK(clk), .Q(H7[14]) );
  DFFHQX1 G_reg_14_ ( .D(n2620), .CK(clk), .Q(SHA256_result[46]) );
  DFFHQX2 H6_reg_2_ ( .D(n2663), .CK(clk), .Q(H6[2]) );
  DFFHQX2 G_reg_8_ ( .D(n2626), .CK(clk), .Q(SHA256_result[40]) );
  DFFHQX1 E_reg_18_ ( .D(n2839), .CK(clk), .Q(SHA256_result[114]) );
  DFFHQX1 E_reg_20_ ( .D(n2837), .CK(clk), .Q(SHA256_result[116]) );
  DFFHQX2 H1_reg_1_ ( .D(n2985), .CK(clk), .Q(H1[1]) );
  DFFX4 A_reg_0_ ( .D(n3018), .CK(clk), .Q(n92), .QN(n93) );
  DFFX4 H7_reg_1_ ( .D(n2569), .CK(clk), .Q(n109) );
  DFFHQX4 E_reg_5_ ( .D(n2852), .CK(clk), .Q(SHA256_result[101]) );
  DFFHQX4 G_reg_6_ ( .D(n2628), .CK(clk), .Q(SHA256_result[38]) );
  DFFHQX2 F_reg_11_ ( .D(n2814), .CK(clk), .Q(SHA256_result[75]) );
  DFFHQX2 F_reg_6_ ( .D(n2819), .CK(clk), .Q(SHA256_result[70]) );
  DFFHQXL A_reg_22_ ( .D(n2996), .CK(clk), .Q(SHA256_result[246]) );
  DFFHQX2 C_reg_3_ ( .D(n2918), .CK(clk), .Q(SHA256_result[163]) );
  DFFHQX4 E_reg_3_ ( .D(n2854), .CK(clk), .Q(SHA256_result[99]) );
  DFFHQX4 E_reg_14_ ( .D(n2843), .CK(clk), .Q(SHA256_result[110]) );
  DFFHQX2 B_reg_3_ ( .D(n2951), .CK(clk), .Q(SHA256_result[195]) );
  DFFHQX4 E_reg_25_ ( .D(n2832), .CK(clk), .Q(SHA256_result[121]) );
  DFFHQX4 G_reg_2_ ( .D(n2632), .CK(clk), .Q(SHA256_result[34]) );
  DFFHQX2 Kt_reg_13_ ( .D(N3015), .CK(clk), .Q(Kt[13]) );
  DFFHQX4 G_reg_4_ ( .D(n2630), .CK(clk), .Q(SHA256_result[36]) );
  DFFHQX4 F_reg_4_ ( .D(n2821), .CK(clk), .Q(SHA256_result[68]) );
  DFFHQX4 C_reg_2_ ( .D(n2919), .CK(clk), .Q(SHA256_result[162]) );
  INVX1 U3 ( .A(n1437), .Y(n315) );
  OAI21XL U4 ( .A0(n181), .A1(SHA256_result[194]), .B0(SHA256_result[162]), 
        .Y(n572) );
  INVX12 U5 ( .A(n41), .Y(n327) );
  NOR2XL U15 ( .A(first_block_core), .B(n324), .Y(n41) );
  OAI2BB1X4 U16 ( .A0N(N1005), .A1N(n238), .B0(n424), .Y(n2831) );
  OAI211X4 U17 ( .A0(n26), .A1(n399), .B0(n358), .C0(n357), .Y(n2630) );
  OAI211X4 U18 ( .A0(n324), .A1(n402), .B0(n61), .C0(n1539), .Y(n2662) );
  INVX1 U19 ( .A(SHA256_result[35]), .Y(n402) );
  MX2X2 U20 ( .A(SHA256_result[49]), .B(SHA256_result[81]), .S0(n148), .Y(
        f1_EFG_32[17]) );
  OAI211XL U21 ( .A0(n324), .A1(n401), .B0(n58), .C0(n1608), .Y(n2790) );
  INVX1 U22 ( .A(SHA256_result[67]), .Y(n401) );
  NAND2XL U23 ( .A(n403), .B(SHA256_result[98]), .Y(n80) );
  CLKINVX3 U24 ( .A(SHA256_result[66]), .Y(n403) );
  XOR3X4 U25 ( .A(n77), .B(SHA256_result[109]), .C(SHA256_result[114]), .Y(
        f4_E_32[7]) );
  INVX12 U26 ( .A(n75), .Y(n77) );
  NAND2X4 U27 ( .A(n42), .B(n577), .Y(n2988) );
  NAND2X4 U28 ( .A(N881), .B(n248), .Y(n577) );
  INVX12 U29 ( .A(n1456), .Y(n10) );
  INVX12 U30 ( .A(n1456), .Y(n11) );
  INVX1 U31 ( .A(n284), .Y(n12) );
  INVX1 U32 ( .A(n285), .Y(n13) );
  INVX1 U33 ( .A(n286), .Y(n14) );
  INVX1 U34 ( .A(n287), .Y(n15) );
  INVX1 U35 ( .A(n312), .Y(n16) );
  CLKINVX2 U36 ( .A(n313), .Y(n17) );
  INVX1 U37 ( .A(n314), .Y(n18) );
  INVX1 U38 ( .A(n303), .Y(n19) );
  INVX1 U39 ( .A(n302), .Y(n20) );
  INVX1 U40 ( .A(n310), .Y(n21) );
  INVX1 U41 ( .A(n311), .Y(n22) );
  INVX1 U42 ( .A(n308), .Y(n23) );
  INVX1 U43 ( .A(n307), .Y(n24) );
  INVX1 U44 ( .A(n309), .Y(n25) );
  INVX1 U45 ( .A(n306), .Y(n26) );
  INVX1 U46 ( .A(n305), .Y(n27) );
  INVX1 U47 ( .A(n304), .Y(n28) );
  CLKINVX8 U48 ( .A(n289), .Y(n29) );
  CLKINVX4 U49 ( .A(n290), .Y(n30) );
  INVX1 U50 ( .A(n293), .Y(n31) );
  CLKINVX3 U51 ( .A(n295), .Y(n32) );
  INVX1 U52 ( .A(n291), .Y(n33) );
  CLKINVX3 U53 ( .A(n288), .Y(n34) );
  CLKINVX3 U54 ( .A(n294), .Y(n35) );
  CLKINVX8 U55 ( .A(n292), .Y(n36) );
  INVX1 U56 ( .A(n298), .Y(n289) );
  INVX1 U57 ( .A(n298), .Y(n290) );
  OR3X1 U58 ( .A(n1849), .B(n341), .C(n340), .Y(n1456) );
  INVX1 U59 ( .A(n312), .Y(n299) );
  NAND2X4 U60 ( .A(n117), .B(n1454), .Y(n2571) );
  OAI211X4 U61 ( .A0(n324), .A1(n94), .B0(n61), .C0(n1541), .Y(n2665) );
  BUFX4 U62 ( .A(SHA256_result[249]), .Y(n159) );
  MX2X4 U63 ( .A(SHA256_result[46]), .B(SHA256_result[78]), .S0(
        SHA256_result[110]), .Y(f1_EFG_32[14]) );
  XOR3X4 U64 ( .A(n180), .B(n169), .C(n161), .Y(f3_A_32[1]) );
  BUFX8 U65 ( .A(SHA256_result[238]), .Y(n169) );
  BUFX4 U66 ( .A(SHA256_result[240]), .Y(n167) );
  MXI2X4 U67 ( .A(n402), .B(n401), .S0(SHA256_result[99]), .Y(f1_EFG_32[3]) );
  OAI21X1 U68 ( .A0(n180), .A1(SHA256_result[195]), .B0(SHA256_result[163]), 
        .Y(n571) );
  XOR3X4 U69 ( .A(n178), .B(n167), .C(n159), .Y(f3_A_32[3]) );
  OAI21X2 U70 ( .A0(SHA256_result[197]), .A1(n178), .B0(SHA256_result[165]), 
        .Y(n569) );
  OAI2BB1X4 U71 ( .A0N(SHA256_result[197]), .A1N(n178), .B0(n569), .Y(
        f2_ABC_32[5]) );
  BUFX4 U72 ( .A(SHA256_result[229]), .Y(n178) );
  CLKBUFX8 U73 ( .A(SHA256_result[246]), .Y(n37) );
  OAI211XL U74 ( .A0(n26), .A1(n397), .B0(n355), .C0(n354), .Y(n2629) );
  CLKINVX3 U75 ( .A(SHA256_result[69]), .Y(n397) );
  INVX1 U76 ( .A(SHA256_result[37]), .Y(n398) );
  MXI2X2 U77 ( .A(n405), .B(n116), .S0(n74), .Y(f1_EFG_32[1]) );
  MX2X4 U78 ( .A(SHA256_result[43]), .B(SHA256_result[75]), .S0(
        SHA256_result[107]), .Y(f1_EFG_32[11]) );
  MX2X4 U79 ( .A(SHA256_result[38]), .B(SHA256_result[70]), .S0(n154), .Y(
        f1_EFG_32[6]) );
  MXI2X4 U80 ( .A(n400), .B(n399), .S0(SHA256_result[100]), .Y(f1_EFG_32[4])
         );
  CLKINVX3 U81 ( .A(SHA256_result[68]), .Y(n399) );
  MXI2X4 U82 ( .A(n398), .B(n397), .S0(SHA256_result[101]), .Y(f1_EFG_32[5])
         );
  OAI21X2 U83 ( .A0(n187), .A1(n761), .B0(n1785), .Y(n2953) );
  OAI2BB1X4 U84 ( .A0N(n197), .A1N(SHA256_result[191]), .B0(n1723), .Y(n2890)
         );
  AND2X4 U85 ( .A(n121), .B(n122), .Y(n1724) );
  NAND2X4 U86 ( .A(N945), .B(n238), .Y(n121) );
  CLKINVX8 U87 ( .A(N978), .Y(n125) );
  INVX4 U88 ( .A(n92), .Y(n69) );
  OAI2BB2XL U89 ( .B0(n327), .B1(n761), .A0N(H1[1]), .A1N(n261), .Y(n2985) );
  OAI2BB1X4 U90 ( .A0N(SHA256_result[194]), .A1N(n181), .B0(n572), .Y(
        f2_ABC_32[2]) );
  BUFX12 U91 ( .A(SHA256_result[226]), .Y(n181) );
  XOR3X2 U92 ( .A(n152), .B(SHA256_result[110]), .C(SHA256_result[124]), .Y(
        f4_E_32[3]) );
  XOR3X2 U93 ( .A(n153), .B(SHA256_result[109]), .C(n73), .Y(f4_E_32[2]) );
  XOR3X2 U94 ( .A(SHA256_result[107]), .B(SHA256_result[112]), .C(n145), .Y(
        f4_E_32[5]) );
  INVXL U95 ( .A(n283), .Y(n313) );
  CLKINVX3 U96 ( .A(n1491), .Y(n340) );
  INVX1 U97 ( .A(n200), .Y(n199) );
  CLKBUFX8 U98 ( .A(SHA256_result[254]), .Y(n155) );
  BUFX4 U99 ( .A(SHA256_result[115]), .Y(n147) );
  BUFX3 U100 ( .A(SHA256_result[253]), .Y(n156) );
  INVX1 U101 ( .A(n297), .Y(n292) );
  NOR2X1 U102 ( .A(n54), .B(n46), .Y(n53) );
  XOR3X2 U103 ( .A(SHA256_result[103]), .B(n150), .C(SHA256_result[122]), .Y(
        f4_E_32[1]) );
  MX2X1 U104 ( .A(SHA256_result[51]), .B(SHA256_result[83]), .S0(n147), .Y(
        f1_EFG_32[19]) );
  MX2X2 U105 ( .A(SHA256_result[39]), .B(SHA256_result[71]), .S0(
        SHA256_result[103]), .Y(f1_EFG_32[7]) );
  OAI2BB1X1 U106 ( .A0N(SHA256_result[195]), .A1N(n180), .B0(n571), .Y(
        f2_ABC_32[3]) );
  XOR3X2 U107 ( .A(n181), .B(n170), .C(n37), .Y(f3_A_32[0]) );
  NAND2X1 U108 ( .A(n1859), .B(n1337), .Y(n341) );
  INVX1 U109 ( .A(n185), .Y(n184) );
  BUFX3 U110 ( .A(SHA256_result[123]), .Y(n73) );
  NAND2BX1 U111 ( .AN(n1859), .B(round[6]), .Y(n339) );
  BUFX3 U112 ( .A(SHA256_result[251]), .Y(n157) );
  CLKINVX3 U113 ( .A(SHA256_result[96]), .Y(n75) );
  BUFX3 U114 ( .A(SHA256_result[247]), .Y(n161) );
  INVX4 U115 ( .A(n75), .Y(n76) );
  BUFX3 U116 ( .A(n101), .Y(n71) );
  CLKBUFX8 U117 ( .A(SHA256_result[105]), .Y(n152) );
  CLKBUFX8 U118 ( .A(SHA256_result[102]), .Y(n154) );
  BUFX3 U119 ( .A(SHA256_result[250]), .Y(n158) );
  CLKBUFX8 U120 ( .A(SHA256_result[104]), .Y(n153) );
  BUFX4 U121 ( .A(SHA256_result[108]), .Y(n150) );
  INVX12 U122 ( .A(n267), .Y(n261) );
  BUFX3 U123 ( .A(SHA256_result[237]), .Y(n170) );
  BUFX3 U124 ( .A(SHA256_result[243]), .Y(n164) );
  CLKBUFX8 U125 ( .A(SHA256_result[241]), .Y(n166) );
  BUFX3 U126 ( .A(SHA256_result[244]), .Y(n163) );
  BUFX3 U127 ( .A(SHA256_result[242]), .Y(n165) );
  BUFX3 U128 ( .A(SHA256_result[233]), .Y(n174) );
  BUFX3 U129 ( .A(SHA256_result[235]), .Y(n172) );
  BUFX3 U130 ( .A(SHA256_result[234]), .Y(n173) );
  BUFX3 U131 ( .A(SHA256_result[245]), .Y(n162) );
  OAI222XL U132 ( .A0(n749), .A1(n715), .B0(n717), .B1(n2269), .C0(n753), .C1(
        n1397), .Y(n2396) );
  BUFX3 U133 ( .A(SHA256_result[126]), .Y(n145) );
  BUFX3 U134 ( .A(SHA256_result[232]), .Y(n175) );
  BUFX3 U135 ( .A(SHA256_result[113]), .Y(n148) );
  BUFX3 U136 ( .A(SHA256_result[111]), .Y(n149) );
  CLKINVX3 U137 ( .A(SHA256_result[36]), .Y(n400) );
  BUFX3 U138 ( .A(SHA256_result[230]), .Y(n177) );
  BUFX3 U139 ( .A(SHA256_result[236]), .Y(n171) );
  INVX1 U140 ( .A(n300), .Y(n288) );
  BUFX3 U141 ( .A(SHA256_result[117]), .Y(n146) );
  NOR2X1 U142 ( .A(n753), .B(round[0]), .Y(n1878) );
  NOR2X1 U143 ( .A(n758), .B(n183), .Y(n2271) );
  BUFX3 U144 ( .A(round[5]), .Y(n183) );
  OAI221XL U145 ( .A0(n28), .A1(n647), .B0(n675), .B1(n646), .C0(n645), .Y(
        n3011) );
  OAI211X1 U146 ( .A0(n324), .A1(n405), .B0(n68), .C0(n1540), .Y(n2664) );
  OAI21XL U147 ( .A0(n186), .A1(n914), .B0(n1494), .Y(n2604) );
  NAND3X1 U148 ( .A(n99), .B(n100), .C(n1458), .Y(n2572) );
  OR2X2 U149 ( .A(n16), .B(n914), .Y(n99) );
  OR2X2 U150 ( .A(n1457), .B(n947), .Y(n100) );
  AND2X2 U151 ( .A(n105), .B(n270), .Y(n1458) );
  OAI2BB1X1 U152 ( .A0N(n198), .A1N(SHA256_result[158]), .B0(n1692), .Y(n2859)
         );
  AND2X2 U153 ( .A(n83), .B(n84), .Y(n1692) );
  NAND2X1 U154 ( .A(N977), .B(n237), .Y(n83) );
  NAND3X2 U155 ( .A(n1691), .B(n124), .C(n123), .Y(n2858) );
  NAND2X1 U156 ( .A(N866), .B(n248), .Y(n622) );
  OAI211X1 U157 ( .A0(n442), .A1(n22), .B0(n441), .C0(n440), .Y(n2838) );
  NAND3X2 U158 ( .A(n582), .B(n581), .C(n580), .Y(n2989) );
  NAND2X2 U159 ( .A(N880), .B(n248), .Y(n580) );
  OAI2BB1X1 U160 ( .A0N(N875), .A1N(n239), .B0(n599), .Y(n2994) );
  NAND3X1 U161 ( .A(n416), .B(n415), .C(n414), .Y(n2829) );
  OAI2BB1X1 U162 ( .A0N(N995), .A1N(n239), .B0(n450), .Y(n2841) );
  MX2X2 U163 ( .A(SHA256_result[40]), .B(SHA256_result[72]), .S0(n153), .Y(
        f1_EFG_32[8]) );
  AOI21XL U164 ( .A0(N971), .A1(n237), .B0(n275), .Y(n1698) );
  NOR2X4 U165 ( .A(n125), .B(n126), .Y(n127) );
  NAND2X4 U166 ( .A(n120), .B(n53), .Y(n2603) );
  AOI22X2 U167 ( .A0(N1073), .A1(n235), .B0(SHA256_result[94]), .B1(n11), .Y(
        n1494) );
  NAND2X1 U168 ( .A(n404), .B(n78), .Y(n79) );
  CLKINVX3 U169 ( .A(SHA256_result[98]), .Y(n78) );
  CLKINVX3 U170 ( .A(n69), .Y(n70) );
  AOI222X4 U171 ( .A0(n2408), .A1(n330), .B0(n2409), .B1(n333), .C0(n2410), 
        .C1(n1397), .Y(n2401) );
  CLKINVX3 U172 ( .A(n1437), .Y(n59) );
  INVX2 U173 ( .A(n675), .Y(n678) );
  INVX1 U174 ( .A(n59), .Y(n63) );
  INVX1 U175 ( .A(n59), .Y(n62) );
  INVX1 U176 ( .A(n210), .Y(n204) );
  INVXL U177 ( .A(n679), .Y(n266) );
  INVXL U178 ( .A(n137), .Y(n316) );
  INVX1 U179 ( .A(n316), .Y(n325) );
  INVX2 U180 ( .A(n60), .Y(n68) );
  INVXL U181 ( .A(n60), .Y(n57) );
  INVX1 U182 ( .A(n60), .Y(n67) );
  INVX1 U183 ( .A(n60), .Y(n64) );
  INVX1 U184 ( .A(n138), .Y(n636) );
  NOR2BX1 U185 ( .AN(first_block_core), .B(n1490), .Y(n138) );
  NOR3X1 U186 ( .A(n1849), .B(round[6]), .C(n261), .Y(n137) );
  INVX4 U187 ( .A(n1437), .Y(n60) );
  INVX1 U188 ( .A(n130), .Y(n730) );
  CLKINVX3 U189 ( .A(n59), .Y(n61) );
  CLKINVX3 U190 ( .A(n60), .Y(n66) );
  CLKINVX3 U191 ( .A(n60), .Y(n65) );
  CLKINVX3 U192 ( .A(n1456), .Y(n284) );
  CLKINVX3 U193 ( .A(n675), .Y(n237) );
  NOR2X1 U194 ( .A(n1371), .B(n332), .Y(n40) );
  AND2X2 U195 ( .A(n578), .B(n579), .Y(n42) );
  AND2X2 U196 ( .A(n586), .B(n587), .Y(n43) );
  AND2X2 U197 ( .A(n104), .B(n103), .Y(n44) );
  AND2X2 U198 ( .A(n79), .B(n80), .Y(n45) );
  NOR2X1 U199 ( .A(n186), .B(n915), .Y(n46) );
  INVX1 U200 ( .A(n316), .Y(n326) );
  NOR2X1 U201 ( .A(n1371), .B(n182), .Y(n47) );
  NOR2X2 U202 ( .A(read_counter[3]), .B(read_counter[2]), .Y(n48) );
  NOR2X2 U203 ( .A(n949), .B(read_counter[3]), .Y(n49) );
  AND2X2 U204 ( .A(read_counter[3]), .B(read_counter[2]), .Y(n50) );
  AND2X2 U205 ( .A(read_counter[3]), .B(n949), .Y(n51) );
  INVX1 U206 ( .A(n85), .Y(n87) );
  INVX1 U207 ( .A(n88), .Y(n90) );
  INVX1 U208 ( .A(n94), .Y(n96) );
  NOR2X1 U209 ( .A(n1384), .B(round[2]), .Y(n136) );
  NOR2XL U210 ( .A(n1384), .B(n1389), .Y(n2349) );
  AOI21X1 U211 ( .A0(n213), .A1(n155), .B0(n272), .Y(n579) );
  BUFX16 U212 ( .A(T1_32[26]), .Y(n55) );
  DLY1X1 U213 ( .A(next_E[23]), .Y(n52) );
  AND2X1 U214 ( .A(SHA256_result[95]), .B(n10), .Y(n54) );
  BUFX16 U215 ( .A(T1_32[22]), .Y(n56) );
  NAND2X4 U216 ( .A(N1042), .B(n246), .Y(n394) );
  NAND2BX1 U217 ( .AN(n324), .B(first_block_core), .Y(n1437) );
  OAI211X1 U218 ( .A0(n324), .A1(n413), .B0(n61), .C0(n1582), .Y(n2733) );
  OAI211X1 U219 ( .A0(n324), .A1(n487), .B0(n66), .C0(n1591), .Y(n2756) );
  OAI211X1 U220 ( .A0(n324), .A1(n491), .B0(n58), .C0(n1592), .Y(n2757) );
  CLKINVX3 U221 ( .A(n137), .Y(n324) );
  XOR3X2 U222 ( .A(n151), .B(n149), .C(SHA256_result[125]), .Y(f4_E_32[4]) );
  NAND2BX2 U223 ( .AN(n1849), .B(output_enable), .Y(n1491) );
  NAND2BX1 U224 ( .AN(n343), .B(n1491), .Y(n1490) );
  AOI21X1 U225 ( .A0(N1024), .A1(n240), .B0(n275), .Y(n1628) );
  OAI2BB1X4 U226 ( .A0N(N879), .A1N(n239), .B0(n584), .Y(n2990) );
  NAND2X2 U227 ( .A(n43), .B(n585), .Y(n2991) );
  NAND2X4 U228 ( .A(N1009), .B(n246), .Y(n406) );
  NAND2X1 U229 ( .A(N998), .B(n246), .Y(n440) );
  NAND2XL U230 ( .A(N1011), .B(n246), .Y(n392) );
  NAND2XL U231 ( .A(N1003), .B(n246), .Y(n429) );
  NAND2XL U232 ( .A(N986), .B(n246), .Y(n480) );
  NAND2XL U233 ( .A(N993), .B(n246), .Y(n453) );
  NAND2XL U234 ( .A(N989), .B(n246), .Y(n466) );
  NAND2XL U235 ( .A(N1007), .B(n246), .Y(n414) );
  NAND3X2 U236 ( .A(n406), .B(n407), .C(n408), .Y(n2827) );
  OAI2BB1X4 U237 ( .A0N(n238), .A1N(N1010), .B0(n513), .Y(n2826) );
  OAI2BB1X4 U238 ( .A0N(n235), .A1N(N882), .B0(n576), .Y(n2987) );
  OAI2BB1X4 U239 ( .A0N(N1006), .A1N(n248), .B0(n420), .Y(n2830) );
  BUFX12 U240 ( .A(SHA256_result[228]), .Y(n179) );
  INVXL U241 ( .A(next_A[5]), .Y(n654) );
  AOI22XL U242 ( .A0(n2039), .A1(n70), .B0(n2040), .B1(n179), .Y(n2214) );
  INVX1 U243 ( .A(n315), .Y(n58) );
  CLKBUFX2 U244 ( .A(n101), .Y(n72) );
  AOI22X1 U245 ( .A0(N1052), .A1(n235), .B0(SHA256_result[73]), .B1(n10), .Y(
        n1515) );
  NAND2XL U246 ( .A(H7[0]), .B(n258), .Y(n1453) );
  NAND2X1 U247 ( .A(N1105), .B(n244), .Y(n105) );
  MX2X4 U248 ( .A(n96), .B(n108), .S0(n77), .Y(f1_EFG_32[0]) );
  MX2X4 U249 ( .A(SHA256_result[45]), .B(SHA256_result[77]), .S0(
        SHA256_result[109]), .Y(f1_EFG_32[13]) );
  AND2X4 U250 ( .A(n118), .B(n119), .Y(n1454) );
  MX2X4 U251 ( .A(SHA256_result[42]), .B(SHA256_result[74]), .S0(n151), .Y(
        f1_EFG_32[10]) );
  NAND2X4 U252 ( .A(N1041), .B(n246), .Y(n97) );
  BUFX16 U253 ( .A(SHA256_result[97]), .Y(n74) );
  NOR2X1 U254 ( .A(n330), .B(round[0]), .Y(n130) );
  INVXL U255 ( .A(SHA256_result[34]), .Y(n404) );
  OAI2BB1X4 U256 ( .A0N(n198), .A1N(SHA256_result[222]), .B0(n1756), .Y(n2924)
         );
  NAND2X4 U257 ( .A(N913), .B(n237), .Y(n81) );
  NAND2XL U258 ( .A(n155), .B(n10), .Y(n82) );
  AND2X4 U259 ( .A(n81), .B(n82), .Y(n1756) );
  INVXL U260 ( .A(next_A[7]), .Y(n647) );
  NAND2XL U261 ( .A(SHA256_result[190]), .B(n10), .Y(n84) );
  NOR2X4 U262 ( .A(n127), .B(n275), .Y(n1691) );
  NAND2X4 U263 ( .A(n44), .B(n1755), .Y(n2923) );
  AOI21X4 U264 ( .A0(N914), .A1(n241), .B0(n278), .Y(n1755) );
  AOI2BB2X4 U265 ( .B0(N946), .B1(n238), .A0N(n759), .A1N(n34), .Y(n1723) );
  INVX1 U266 ( .A(n350), .Y(n1457) );
  OAI2BB1X1 U267 ( .A0N(n197), .A1N(SHA256_result[94]), .B0(n1611), .Y(n2795)
         );
  AND2X2 U268 ( .A(n97), .B(n98), .Y(n1611) );
  INVX1 U269 ( .A(SHA256_result[62]), .Y(n914) );
  INVX1 U270 ( .A(SHA256_result[30]), .Y(n947) );
  NAND2XL U271 ( .A(n145), .B(n10), .Y(n98) );
  OR2X2 U272 ( .A(n13), .B(n700), .Y(n103) );
  OR2X2 U273 ( .A(n223), .B(n759), .Y(n104) );
  OAI211X2 U274 ( .A0(n14), .A1(n511), .B0(n394), .C0(n395), .Y(n2794) );
  OAI211XL U275 ( .A0(n317), .A1(n821), .B0(n67), .C0(n1580), .Y(n2728) );
  NAND2X4 U276 ( .A(N1106), .B(n237), .Y(n118) );
  INVX1 U277 ( .A(n279), .Y(n273) );
  INVX1 U278 ( .A(n249), .Y(n244) );
  INVX1 U279 ( .A(n106), .Y(n108) );
  NAND2X1 U280 ( .A(SHA256_result[63]), .B(n10), .Y(n119) );
  OAI2BB1X1 U281 ( .A0N(SHA256_result[193]), .A1N(n72), .B0(n573), .Y(
        f2_ABC_32[1]) );
  MX2X4 U282 ( .A(SHA256_result[41]), .B(SHA256_result[73]), .S0(n152), .Y(
        f1_EFG_32[9]) );
  OAI2BB2XL U283 ( .B0(n327), .B1(n820), .A0N(n112), .A1N(n265), .Y(n2729) );
  OAI21XL U284 ( .A0(SHA256_result[193]), .A1(n72), .B0(n87), .Y(n573) );
  OAI211X1 U285 ( .A0(n26), .A1(n401), .B0(n360), .C0(n359), .Y(n2631) );
  OAI2BB2XL U286 ( .B0(n327), .B1(n918), .A0N(n109), .A1N(n264), .Y(n2569) );
  CLKINVX2 U287 ( .A(n675), .Y(n235) );
  INVX1 U288 ( .A(n675), .Y(n238) );
  INVX1 U289 ( .A(SHA256_result[191]), .Y(n818) );
  OAI211XL U290 ( .A0(n318), .A1(n917), .B0(n68), .C0(n1453), .Y(n2570) );
  NAND2X4 U291 ( .A(N1074), .B(n235), .Y(n120) );
  INVX1 U292 ( .A(n216), .Y(n213) );
  INVX1 U293 ( .A(n296), .Y(n295) );
  INVX1 U294 ( .A(n297), .Y(n294) );
  INVX1 U295 ( .A(n299), .Y(n293) );
  INVX1 U296 ( .A(n270), .Y(n278) );
  INVX1 U297 ( .A(n279), .Y(n275) );
  CLKINVX3 U298 ( .A(n326), .Y(n317) );
  NOR2XL U299 ( .A(n191), .B(n597), .Y(n598) );
  NOR2XL U300 ( .A(n130), .B(n2261), .Y(n2519) );
  NAND2X1 U301 ( .A(N870), .B(n248), .Y(n612) );
  OAI211X1 U302 ( .A0(n614), .A1(n34), .B0(n613), .C0(n612), .Y(n2999) );
  NAND2X1 U303 ( .A(N865), .B(n247), .Y(n625) );
  NAND2X1 U304 ( .A(N864), .B(n248), .Y(n628) );
  NAND2X1 U305 ( .A(N860), .B(n248), .Y(n640) );
  NAND2X1 U306 ( .A(N863), .B(n248), .Y(n631) );
  NAND2XL U307 ( .A(n193), .B(n171), .Y(n632) );
  NAND2XL U308 ( .A(N853), .B(n248), .Y(n668) );
  NAND2XL U309 ( .A(N856), .B(n678), .Y(n653) );
  NAND2XL U310 ( .A(N855), .B(n248), .Y(n657) );
  INVXL U311 ( .A(n136), .Y(n754) );
  AOI211XL U312 ( .A0(n722), .A1(round[2]), .B0(n2337), .C0(n2338), .Y(n2336)
         );
  AOI221XL U313 ( .A0(n2267), .A1(n335), .B0(n130), .B1(n40), .C0(n2338), .Y(
        n2383) );
  AOI211XL U314 ( .A0(n722), .A1(n136), .B0(n2286), .C0(n2287), .Y(n2276) );
  AOI21XL U315 ( .A0(n136), .A1(n2473), .B0(n2274), .Y(n2279) );
  XOR3X4 U316 ( .A(n154), .B(SHA256_result[107]), .C(SHA256_result[121]), .Y(
        f4_E_32[0]) );
  INVXL U317 ( .A(SHA256_result[33]), .Y(n405) );
  AOI22X1 U318 ( .A0(N938), .A1(n238), .B0(SHA256_result[215]), .B1(n10), .Y(
        n1731) );
  BUFX4 U319 ( .A(SHA256_result[231]), .Y(n176) );
  BUFX8 U320 ( .A(SHA256_result[248]), .Y(n160) );
  NAND2XL U321 ( .A(N1044), .B(n245), .Y(n365) );
  NAND2XL U322 ( .A(N979), .B(n247), .Y(n508) );
  NAND2XL U323 ( .A(N1014), .B(n247), .Y(n385) );
  NAND2XL U324 ( .A(N1013), .B(n245), .Y(n387) );
  NAND2XL U325 ( .A(N1016), .B(n245), .Y(n379) );
  MX2X1 U326 ( .A(SHA256_result[53]), .B(SHA256_result[85]), .S0(n146), .Y(
        f1_EFG_32[21]) );
  AOI222XL U327 ( .A0(n130), .A1(n2245), .B0(n2318), .B1(n336), .C0(n2427), 
        .C1(n1397), .Y(n2480) );
  AOI211XL U328 ( .A0(n2520), .A1(n136), .B0(n2446), .C0(n2448), .Y(n2515) );
  INVX1 U329 ( .A(n237), .Y(n126) );
  OAI2BB1X1 U330 ( .A0N(n194), .A1N(SHA256_result[190]), .B0(n1724), .Y(n2891)
         );
  NAND2X1 U331 ( .A(SHA256_result[222]), .B(n11), .Y(n122) );
  OR2X2 U332 ( .A(n705), .B(n916), .Y(n117) );
  OR2X2 U333 ( .A(n14), .B(n818), .Y(n123) );
  OR2X2 U334 ( .A(n233), .B(n819), .Y(n124) );
  INVXL U335 ( .A(n200), .Y(n198) );
  INVXL U336 ( .A(n201), .Y(n196) );
  OAI2BB1X2 U337 ( .A0N(N874), .A1N(n236), .B0(n603), .Y(n2995) );
  NAND2XL U338 ( .A(n343), .B(n1491), .Y(n674) );
  NAND2XL U339 ( .A(n1490), .B(n1491), .Y(n350) );
  INVXL U340 ( .A(n1456), .Y(n285) );
  INVXL U341 ( .A(n1456), .Y(n286) );
  INVXL U342 ( .A(n261), .Y(n251) );
  INVXL U343 ( .A(n1456), .Y(n287) );
  AOI222XL U344 ( .A0(n2427), .A1(n2258), .B0(n2409), .B1(n2428), .C0(n2429), 
        .C1(n333), .Y(n2421) );
  NAND2XL U345 ( .A(n130), .B(n2501), .Y(n2307) );
  AOI21XL U346 ( .A0(n213), .A1(n168), .B0(n272), .Y(n623) );
  AOI21XL U347 ( .A0(n213), .A1(n169), .B0(n272), .Y(n626) );
  AOI21XL U348 ( .A0(n213), .A1(n170), .B0(n273), .Y(n629) );
  AOI21XL U349 ( .A0(n213), .A1(n164), .B0(n272), .Y(n613) );
  AOI21XL U350 ( .A0(n213), .A1(n147), .B0(n278), .Y(n441) );
  NAND2XL U351 ( .A(next_A[30]), .B(n11), .Y(n578) );
  AOI21XL U352 ( .A0(n145), .A1(n212), .B0(n277), .Y(n408) );
  NAND2X2 U353 ( .A(N878), .B(n248), .Y(n585) );
  AOI21XL U354 ( .A0(n214), .A1(n157), .B0(n272), .Y(n587) );
  AOI21XL U355 ( .A0(n213), .A1(n156), .B0(n272), .Y(n582) );
  AOI21XL U356 ( .A0(n159), .A1(n211), .B0(n272), .Y(n595) );
  NOR2XL U357 ( .A(n191), .B(n605), .Y(n606) );
  NOR2XL U358 ( .A(n191), .B(n426), .Y(n427) );
  OAI2BB1X2 U359 ( .A0N(N1002), .A1N(n235), .B0(n433), .Y(n2834) );
  OAI2BB1X2 U360 ( .A0N(N1008), .A1N(n236), .B0(n412), .Y(n2828) );
  AOI21XL U361 ( .A0(next_A[31]), .A1(n11), .B0(n575), .Y(n576) );
  AOI21XL U362 ( .A0(next_E[31]), .A1(n11), .B0(n512), .Y(n513) );
  NOR2XL U363 ( .A(n191), .B(n422), .Y(n423) );
  INVXL U364 ( .A(next_E[10]), .Y(n468) );
  AOI21XL U365 ( .A0(n212), .A1(n148), .B0(n273), .Y(n447) );
  NAND2XL U366 ( .A(N996), .B(n246), .Y(n446) );
  INVXL U367 ( .A(next_E[9]), .Y(n472) );
  NAND2XL U368 ( .A(N988), .B(n246), .Y(n471) );
  AOI21XL U369 ( .A0(n152), .A1(n212), .B0(n277), .Y(n470) );
  AOI21XL U370 ( .A0(n214), .A1(n174), .B0(n273), .Y(n639) );
  AOI21XL U371 ( .A0(n212), .A1(n150), .B0(n273), .Y(n458) );
  AOI22XL U372 ( .A0(next_E[12]), .A1(n10), .B0(N991), .B1(n239), .Y(n459) );
  INVXL U373 ( .A(next_A[8]), .Y(n644) );
  INVXL U374 ( .A(next_E[8]), .Y(n477) );
  NAND2XL U375 ( .A(N987), .B(n246), .Y(n475) );
  OR2X2 U376 ( .A(n340), .B(n128), .Y(n675) );
  OR2XL U377 ( .A(n1849), .B(n339), .Y(n128) );
  AOI21XL U378 ( .A0(N1098), .A1(n244), .B0(n275), .Y(n1466) );
  AOI21XL U379 ( .A0(N1097), .A1(n244), .B0(n273), .Y(n1467) );
  AOI21XL U380 ( .A0(N1096), .A1(n244), .B0(n277), .Y(n1468) );
  AOI21XL U381 ( .A0(N1089), .A1(n244), .B0(n277), .Y(n1475) );
  AOI21XL U382 ( .A0(N1085), .A1(n243), .B0(n274), .Y(n1479) );
  AOI21XL U383 ( .A0(N1083), .A1(n243), .B0(n271), .Y(n1481) );
  AOI21XL U384 ( .A0(N901), .A1(n241), .B0(n278), .Y(n1768) );
  AOI21XL U385 ( .A0(N900), .A1(n241), .B0(n278), .Y(n1769) );
  AOI21XL U386 ( .A0(N898), .A1(n242), .B0(n278), .Y(n1771) );
  AOI21XL U387 ( .A0(N933), .A1(n237), .B0(n277), .Y(n1736) );
  AOI21XL U388 ( .A0(N932), .A1(n240), .B0(n277), .Y(n1737) );
  AOI21XL U389 ( .A0(N934), .A1(n240), .B0(n277), .Y(n1735) );
  AOI21XL U390 ( .A0(N1051), .A1(n242), .B0(n274), .Y(n1516) );
  AOI21XL U391 ( .A0(N1054), .A1(n243), .B0(n274), .Y(n1513) );
  AOI21XL U392 ( .A0(N930), .A1(n240), .B0(n277), .Y(n1739) );
  AOI21XL U393 ( .A0(N929), .A1(n240), .B0(n277), .Y(n1740) );
  AOI21XL U394 ( .A0(N1066), .A1(n243), .B0(n274), .Y(n1501) );
  AOI21XL U395 ( .A0(N899), .A1(n242), .B0(n278), .Y(n1770) );
  AOI21XL U396 ( .A0(N893), .A1(n242), .B0(n273), .Y(n1776) );
  AOI21XL U397 ( .A0(N890), .A1(n242), .B0(n272), .Y(n1779) );
  AOI21XL U398 ( .A0(N1050), .A1(n242), .B0(n274), .Y(n1517) );
  AOI21XL U399 ( .A0(N924), .A1(n241), .B0(n277), .Y(n1745) );
  AOI21XL U400 ( .A0(N921), .A1(n240), .B0(n277), .Y(n1748) );
  AOI21XL U401 ( .A0(N1055), .A1(n243), .B0(n274), .Y(n1512) );
  AOI22XL U402 ( .A0(N906), .A1(n238), .B0(n161), .B1(n10), .Y(n1763) );
  AOI22XL U403 ( .A0(N1026), .A1(n236), .B0(n149), .B1(n10), .Y(n1626) );
  AOI22XL U404 ( .A0(N1023), .A1(n236), .B0(n150), .B1(n11), .Y(n1629) );
  AOI22XL U405 ( .A0(N1021), .A1(n236), .B0(n151), .B1(n10), .Y(n1631) );
  AOI22XL U406 ( .A0(N1020), .A1(n236), .B0(n152), .B1(n11), .Y(n1632) );
  AOI22XL U407 ( .A0(N1019), .A1(n237), .B0(n153), .B1(n11), .Y(n1633) );
  AOI22XL U408 ( .A0(N902), .A1(n237), .B0(n164), .B1(n11), .Y(n1767) );
  AOI22XL U409 ( .A0(N1017), .A1(n237), .B0(n154), .B1(n10), .Y(n1635) );
  AOI22XL U410 ( .A0(N887), .A1(n238), .B0(n179), .B1(n11), .Y(n1782) );
  AOI22XL U411 ( .A0(N884), .A1(n238), .B0(n72), .B1(n11), .Y(n1785) );
  AOI22XL U412 ( .A0(N888), .A1(n239), .B0(n178), .B1(n11), .Y(n1781) );
  AOI22XL U413 ( .A0(N886), .A1(n242), .B0(n180), .B1(n10), .Y(n1783) );
  INVXL U414 ( .A(next_A[6]), .Y(n650) );
  AOI21XL U415 ( .A0(n214), .A1(n177), .B0(n273), .Y(n648) );
  AOI21XL U416 ( .A0(n178), .A1(n211), .B0(n273), .Y(n652) );
  AOI21XL U417 ( .A0(n181), .A1(n211), .B0(n273), .Y(n667) );
  INVXL U418 ( .A(next_A[1]), .Y(n673) );
  NAND2XL U419 ( .A(N852), .B(n244), .Y(n672) );
  AOI21XL U420 ( .A0(n72), .A1(n211), .B0(n273), .Y(n671) );
  INVXL U421 ( .A(next_E[6]), .Y(n486) );
  NAND2XL U422 ( .A(N985), .B(n246), .Y(n485) );
  AOI21XL U423 ( .A0(n154), .A1(n212), .B0(n271), .Y(n484) );
  INVXL U424 ( .A(next_A[4]), .Y(n659) );
  AOI2BB2XL U425 ( .B0(N950), .B1(n239), .A0N(n26), .A1N(n519), .Y(n514) );
  AOI2BB2XL U426 ( .B0(N948), .B1(n239), .A0N(n29), .A1N(n85), .Y(n516) );
  AOI2BB2XL U427 ( .B0(N905), .B1(n239), .A0N(n25), .A1N(n605), .Y(n537) );
  AOI2BB2XL U428 ( .B0(N885), .B1(n239), .A0N(n16), .A1N(n666), .Y(n539) );
  AOI22XL U429 ( .A0(next_A[0]), .A1(n10), .B0(n70), .B1(n211), .Y(n677) );
  AOI21XL U430 ( .A0(N851), .A1(n248), .B0(n273), .Y(n676) );
  INVX1 U431 ( .A(n331), .Y(n330) );
  INVXL U432 ( .A(next_A[3]), .Y(n665) );
  INVX1 U433 ( .A(n144), .Y(n268) );
  AOI222XL U434 ( .A0(n2399), .A1(n1397), .B0(n2308), .B1(n131), .C0(n2400), 
        .C1(n333), .Y(n2393) );
  AOI31XL U435 ( .A0(n742), .A1(n336), .A2(n2349), .B0(n1878), .Y(n2334) );
  AOI22XL U436 ( .A0(n2325), .A1(n129), .B0(n2261), .B1(n2271), .Y(n2327) );
  AOI211XL U437 ( .A0(n2465), .A1(n333), .B0(n2496), .C0(n2537), .Y(n2534) );
  AOI22XL U438 ( .A0(n136), .A1(n2375), .B0(n2486), .B1(n329), .Y(n2528) );
  AOI222XL U439 ( .A0(n2479), .A1(n333), .B0(n2310), .B1(n47), .C0(n2299), 
        .C1(n129), .Y(n2511) );
  AOI222XL U440 ( .A0(n2313), .A1(round[2]), .B0(n2308), .B1(n333), .C0(n2312), 
        .C1(n708), .Y(n2505) );
  AOI211XL U441 ( .A0(n2391), .A1(n136), .B0(n2406), .C0(n2471), .Y(n2467) );
  AOI222XL U442 ( .A0(n2344), .A1(n131), .B0(n2447), .B1(n130), .C0(n2438), 
        .C1(n47), .Y(n2440) );
  AOI222XL U443 ( .A0(n743), .A1(n329), .B0(n2438), .B1(n333), .C0(n2370), 
        .C1(n183), .Y(n2430) );
  AOI222XL U444 ( .A0(n2427), .A1(n330), .B0(n2410), .B1(n129), .C0(n2437), 
        .C1(n2391), .Y(n2431) );
  NOR2X1 U445 ( .A(round[0]), .B(n335), .Y(n129) );
  NOR2XL U446 ( .A(n330), .B(n328), .Y(n2258) );
  OAI32XL U447 ( .A0(n742), .A1(n335), .A2(n758), .B0(round[2]), .B1(n2367), 
        .Y(n2366) );
  AOI31XL U448 ( .A0(n756), .A1(n714), .A2(n723), .B0(n333), .Y(n2463) );
  AOI21XL U449 ( .A0(round[2]), .A1(n130), .B0(n2247), .Y(n2241) );
  AOI31XL U450 ( .A0(n183), .A1(round[2]), .A2(n130), .B0(n2527), .Y(n2526) );
  NOR2X1 U451 ( .A(n332), .B(n183), .Y(n131) );
  NOR2XL U452 ( .A(n328), .B(n758), .Y(n2310) );
  AOI21XL U453 ( .A0(n753), .A1(n2296), .B0(n330), .Y(n2426) );
  NAND2XL U454 ( .A(n136), .B(n183), .Y(n2269) );
  NOR2XL U455 ( .A(n330), .B(n183), .Y(n2391) );
  OAI2BB1X4 U456 ( .A0N(n338), .A1N(n337), .B0(n1434), .Y(n1849) );
  OAI211XL U457 ( .A0(n317), .A1(n928), .B0(n65), .C0(n1448), .Y(n2559) );
  NAND2XL U458 ( .A(H7[11]), .B(n260), .Y(n1448) );
  OAI211XL U459 ( .A0(n318), .A1(n927), .B0(n68), .C0(n1449), .Y(n2560) );
  NAND2XL U460 ( .A(H7[10]), .B(n260), .Y(n1449) );
  OAI211XL U461 ( .A0(n318), .A1(n925), .B0(n64), .C0(n1450), .Y(n2562) );
  NAND2XL U462 ( .A(H7[8]), .B(n260), .Y(n1450) );
  OAI211XL U463 ( .A0(n318), .A1(n921), .B0(n66), .C0(n1451), .Y(n2566) );
  OAI211XL U464 ( .A0(n318), .A1(n920), .B0(n62), .C0(n1452), .Y(n2567) );
  OAI211XL U465 ( .A0(n319), .A1(n895), .B0(n61), .C0(n1535), .Y(n2654) );
  NAND2XL U466 ( .A(H6[11]), .B(n259), .Y(n1535) );
  OAI211XL U467 ( .A0(n319), .A1(n892), .B0(n63), .C0(n1536), .Y(n2657) );
  NAND2XL U468 ( .A(H6[8]), .B(n259), .Y(n1536) );
  OAI211XL U469 ( .A0(n319), .A1(n891), .B0(n64), .C0(n1537), .Y(n2658) );
  NAND2XL U470 ( .A(H6[7]), .B(n259), .Y(n1537) );
  OAI211XL U471 ( .A0(n321), .A1(n870), .B0(n68), .C0(n1606), .Y(n2782) );
  NAND2XL U472 ( .A(H5[11]), .B(n254), .Y(n1606) );
  OAI211XL U473 ( .A0(n321), .A1(n866), .B0(n64), .C0(n1607), .Y(n2786) );
  NAND2XL U474 ( .A(H5[7]), .B(n254), .Y(n1607) );
  INVXL U475 ( .A(n150), .Y(n851) );
  OAI211XL U476 ( .A0(n317), .A1(n830), .B0(n61), .C0(n1575), .Y(n2719) );
  OAI211XL U477 ( .A0(n317), .A1(n828), .B0(n68), .C0(n1576), .Y(n2721) );
  NAND2XL U478 ( .A(H3[8]), .B(n256), .Y(n1576) );
  OAI211XL U479 ( .A0(n317), .A1(n825), .B0(n62), .C0(n1577), .Y(n2724) );
  OAI211XL U480 ( .A0(n317), .A1(n824), .B0(n62), .C0(n1578), .Y(n2725) );
  NAND2XL U481 ( .A(H3[4]), .B(n256), .Y(n1578) );
  OAI211XL U482 ( .A0(n317), .A1(n823), .B0(n64), .C0(n1579), .Y(n2726) );
  NAND2XL U483 ( .A(H3[1]), .B(n256), .Y(n1580) );
  OAI211XL U484 ( .A0(n320), .A1(n796), .B0(n68), .C0(n1556), .Y(n2689) );
  NAND2XL U485 ( .A(H2[9]), .B(n257), .Y(n1556) );
  OAI211XL U486 ( .A0(n320), .A1(n795), .B0(n63), .C0(n1557), .Y(n2690) );
  NAND2XL U487 ( .A(H2[8]), .B(n257), .Y(n1557) );
  OAI211XL U488 ( .A0(n320), .A1(n793), .B0(n61), .C0(n1558), .Y(n2692) );
  NAND2XL U489 ( .A(H2[6]), .B(n257), .Y(n1558) );
  OAI211XL U490 ( .A0(n320), .A1(n792), .B0(n66), .C0(n1559), .Y(n2693) );
  OAI211XL U491 ( .A0(n320), .A1(n791), .B0(n67), .C0(n1560), .Y(n2694) );
  NAND2XL U492 ( .A(H2[4]), .B(n257), .Y(n1560) );
  NAND2XL U493 ( .A(H2[1]), .B(n257), .Y(n1561) );
  OAI211XL U494 ( .A0(n322), .A1(n771), .B0(n63), .C0(n1800), .Y(n2975) );
  NAND2XL U495 ( .A(H1[11]), .B(n253), .Y(n1800) );
  OAI211XL U496 ( .A0(n322), .A1(n770), .B0(n65), .C0(n1801), .Y(n2976) );
  OAI211XL U497 ( .A0(n322), .A1(n769), .B0(n65), .C0(n1802), .Y(n2977) );
  NAND2XL U498 ( .A(H1[9]), .B(n253), .Y(n1802) );
  OAI211XL U499 ( .A0(n322), .A1(n767), .B0(n66), .C0(n1803), .Y(n2979) );
  NAND2XL U500 ( .A(H1[7]), .B(n253), .Y(n1803) );
  OAI211XL U501 ( .A0(n322), .A1(n762), .B0(n66), .C0(n1804), .Y(n2984) );
  OAI211XL U502 ( .A0(n317), .A1(n941), .B0(n65), .C0(n1442), .Y(n2546) );
  NAND2XL U503 ( .A(H7[24]), .B(n261), .Y(n1442) );
  OAI211XL U504 ( .A0(n317), .A1(n940), .B0(n62), .C0(n1443), .Y(n2547) );
  NAND2XL U505 ( .A(H7[23]), .B(n261), .Y(n1443) );
  OAI211XL U506 ( .A0(n317), .A1(n939), .B0(n66), .C0(n1444), .Y(n2548) );
  NAND2XL U507 ( .A(H7[22]), .B(n261), .Y(n1444) );
  OAI211XL U508 ( .A0(n317), .A1(n938), .B0(n67), .C0(n1445), .Y(n2549) );
  NAND2XL U509 ( .A(H7[21]), .B(n261), .Y(n1445) );
  OAI211XL U510 ( .A0(n317), .A1(n398), .B0(n61), .C0(n1538), .Y(n2660) );
  NAND2XL U511 ( .A(H6[5]), .B(n259), .Y(n1538) );
  AOI21XL U512 ( .A0(n212), .A1(SHA256_result[114]), .B0(n273), .Y(n444) );
  NAND2XL U513 ( .A(N997), .B(n246), .Y(n443) );
  AOI2BB2XL U514 ( .B0(n196), .B1(SHA256_result[109]), .A0N(n25), .A1N(n456), 
        .Y(n457) );
  AOI21XL U515 ( .A0(n213), .A1(SHA256_result[95]), .B0(n271), .Y(n395) );
  BUFX8 U516 ( .A(SHA256_result[227]), .Y(n180) );
  CLKBUFX8 U517 ( .A(SHA256_result[106]), .Y(n151) );
  INVXL U518 ( .A(SHA256_result[162]), .Y(n523) );
  NAND2XL U519 ( .A(H2[2]), .B(n257), .Y(n522) );
  NAND2XL U520 ( .A(H2[0]), .B(n260), .Y(n530) );
  INVXL U521 ( .A(n179), .Y(n656) );
  INVXL U522 ( .A(n180), .Y(n661) );
  NAND2XL U523 ( .A(H5[4]), .B(n258), .Y(n381) );
  NAND2XL U524 ( .A(H5[1]), .B(n260), .Y(n388) );
  NAND2XL U525 ( .A(H5[0]), .B(n258), .Y(n391) );
  INVXL U526 ( .A(n151), .Y(n465) );
  INVXL U527 ( .A(n153), .Y(n474) );
  NAND2XL U528 ( .A(H2[3]), .B(n259), .Y(n518) );
  AOI22XL U529 ( .A0(N1040), .A1(n239), .B0(SHA256_result[125]), .B1(n11), .Y(
        n1612) );
  NAND2XL U530 ( .A(H6[3]), .B(n259), .Y(n1539) );
  NAND2XL U531 ( .A(n110), .B(n259), .Y(n1540) );
  NAND2XL U532 ( .A(n114), .B(n257), .Y(n1541) );
  NAND2XL U533 ( .A(H5[3]), .B(n254), .Y(n1608) );
  OAI211XL U534 ( .A0(n324), .A1(n403), .B0(n63), .C0(n1609), .Y(n2791) );
  NAND2XL U535 ( .A(H5[2]), .B(n254), .Y(n1609) );
  NAND3XL U536 ( .A(n132), .B(n64), .C(n1581), .Y(n2731) );
  OR2XL U537 ( .A(n317), .B(n396), .Y(n132) );
  NAND3XL U538 ( .A(n133), .B(n67), .C(n1589), .Y(n2752) );
  OR2XL U539 ( .A(n317), .B(n469), .Y(n133) );
  NAND3XL U540 ( .A(n134), .B(n61), .C(n1590), .Y(n2755) );
  OR2XL U541 ( .A(n317), .B(n483), .Y(n134) );
  NAND3XL U542 ( .A(n135), .B(n65), .C(n1873), .Y(n3045) );
  OR2XL U543 ( .A(n317), .B(n651), .Y(n135) );
  NAND3BXL U544 ( .AN(n670), .B(n66), .C(n1875), .Y(n3049) );
  OAI2BB2XL U545 ( .B0(n327), .B1(n926), .A0N(H7[9]), .A1N(n264), .Y(n2561) );
  OAI2BB2XL U546 ( .B0(n327), .B1(n924), .A0N(H7[7]), .A1N(n264), .Y(n2563) );
  OAI2BB2XL U547 ( .B0(n327), .B1(n923), .A0N(H7[6]), .A1N(n264), .Y(n2564) );
  OAI2BB2XL U548 ( .B0(n327), .B1(n922), .A0N(H7[5]), .A1N(n264), .Y(n2565) );
  OAI2BB2XL U549 ( .B0(n327), .B1(n894), .A0N(H6[10]), .A1N(n265), .Y(n2655)
         );
  OAI2BB2XL U550 ( .B0(n327), .B1(n893), .A0N(H6[9]), .A1N(n265), .Y(n2656) );
  OAI2BB2XL U551 ( .B0(n327), .B1(n890), .A0N(H6[6]), .A1N(n262), .Y(n2659) );
  OAI2BB2XL U552 ( .B0(n327), .B1(n869), .A0N(H5[10]), .A1N(n263), .Y(n2783)
         );
  OAI2BB2XL U553 ( .B0(n327), .B1(n868), .A0N(H5[9]), .A1N(n263), .Y(n2784) );
  OAI2BB2XL U554 ( .B0(n327), .B1(n867), .A0N(H5[8]), .A1N(n263), .Y(n2785) );
  OAI2BB2XL U555 ( .B0(n327), .B1(n865), .A0N(H5[6]), .A1N(n262), .Y(n2787) );
  INVXL U556 ( .A(n149), .Y(n854) );
  OAI2BB2XL U557 ( .B0(n327), .B1(n831), .A0N(H3[11]), .A1N(n263), .Y(n2718)
         );
  OAI2BB2XL U558 ( .B0(n327), .B1(n829), .A0N(H3[9]), .A1N(n265), .Y(n2720) );
  OAI2BB2XL U559 ( .B0(n327), .B1(n827), .A0N(H3[7]), .A1N(n265), .Y(n2722) );
  OAI2BB2XL U560 ( .B0(n327), .B1(n826), .A0N(H3[6]), .A1N(n265), .Y(n2723) );
  OAI2BB2XL U561 ( .B0(n327), .B1(n798), .A0N(H2[11]), .A1N(n264), .Y(n2687)
         );
  OAI2BB2XL U562 ( .B0(n327), .B1(n797), .A0N(H2[10]), .A1N(n265), .Y(n2688)
         );
  OAI2BB2XL U563 ( .B0(n327), .B1(n794), .A0N(H2[7]), .A1N(n262), .Y(n2691) );
  OAI2BB2XL U564 ( .B0(n327), .B1(n768), .A0N(H1[8]), .A1N(n262), .Y(n2978) );
  OAI2BB2XL U565 ( .B0(n327), .B1(n766), .A0N(H1[6]), .A1N(n262), .Y(n2980) );
  OAI2BB2XL U566 ( .B0(n327), .B1(n764), .A0N(H1[4]), .A1N(n262), .Y(n2982) );
  OAI2BB2XL U567 ( .B0(n327), .B1(n691), .A0N(H0[17]), .A1N(n262), .Y(n3033)
         );
  OAI2BB2XL U568 ( .B0(n327), .B1(n685), .A0N(H0[11]), .A1N(n262), .Y(n3039)
         );
  OAI2BB2XL U569 ( .B0(n327), .B1(n682), .A0N(H0[8]), .A1N(n262), .Y(n3042) );
  INVXL U570 ( .A(next_E[16]), .Y(n449) );
  AOI21XL U571 ( .A0(n212), .A1(SHA256_result[120]), .B0(n276), .Y(n431) );
  CLKBUFX8 U572 ( .A(SHA256_result[239]), .Y(n168) );
  NAND2XL U573 ( .A(H6[4]), .B(n258), .Y(n356) );
  NAND2XL U574 ( .A(H5[5]), .B(n258), .Y(n378) );
  NAND2XL U575 ( .A(H6[2]), .B(n258), .Y(n361) );
  AOI21XL U576 ( .A0(n214), .A1(SHA256_result[91]), .B0(n271), .Y(n371) );
  AOI22XL U577 ( .A0(N1033), .A1(n235), .B0(SHA256_result[118]), .B1(n10), .Y(
        n1619) );
  AOI22XL U578 ( .A0(N926), .A1(n237), .B0(SHA256_result[203]), .B1(n10), .Y(
        n1743) );
  AOI22XL U579 ( .A0(N925), .A1(n237), .B0(SHA256_result[202]), .B1(n10), .Y(
        n1744) );
  AOI22XL U580 ( .A0(N922), .A1(n237), .B0(SHA256_result[199]), .B1(n11), .Y(
        n1747) );
  AOI22XL U581 ( .A0(N958), .A1(n237), .B0(SHA256_result[171]), .B1(n11), .Y(
        n1711) );
  AOI22XL U582 ( .A0(N954), .A1(n238), .B0(SHA256_result[167]), .B1(n11), .Y(
        n1715) );
  AOI22XL U583 ( .A0(N947), .A1(n238), .B0(n90), .B1(n10), .Y(n1722) );
  AOI22XL U584 ( .A0(N931), .A1(n238), .B0(SHA256_result[208]), .B1(n10), .Y(
        n1738) );
  AOI22XL U585 ( .A0(N956), .A1(n238), .B0(SHA256_result[169]), .B1(n10), .Y(
        n1713) );
  AOI22XL U586 ( .A0(N953), .A1(n238), .B0(SHA256_result[166]), .B1(n11), .Y(
        n1716) );
  AOI22XL U587 ( .A0(N1034), .A1(n243), .B0(SHA256_result[119]), .B1(n10), .Y(
        n1618) );
  AOI22XL U588 ( .A0(N1065), .A1(n240), .B0(SHA256_result[86]), .B1(n11), .Y(
        n1502) );
  AOI22XL U589 ( .A0(N1061), .A1(n237), .B0(SHA256_result[82]), .B1(n11), .Y(
        n1506) );
  AOI22XL U590 ( .A0(N1056), .A1(n236), .B0(SHA256_result[77]), .B1(n11), .Y(
        n1511) );
  AOI22XL U591 ( .A0(N1053), .A1(n244), .B0(SHA256_result[74]), .B1(n10), .Y(
        n1514) );
  AOI22XL U592 ( .A0(N1049), .A1(n235), .B0(SHA256_result[70]), .B1(n10), .Y(
        n1518) );
  AOI21XL U593 ( .A0(SHA256_result[33]), .A1(n212), .B0(n271), .Y(n364) );
  AOI22XL U594 ( .A0(N1077), .A1(n235), .B0(SHA256_result[34]), .B1(n10), .Y(
        n1487) );
  AOI22XL U595 ( .A0(N1076), .A1(n235), .B0(SHA256_result[33]), .B1(n11), .Y(
        n1488) );
  AOI22XL U596 ( .A0(N1080), .A1(n235), .B0(SHA256_result[37]), .B1(n11), .Y(
        n1484) );
  AOI22XL U597 ( .A0(N1092), .A1(n236), .B0(SHA256_result[49]), .B1(n11), .Y(
        n1472) );
  AOI22XL U598 ( .A0(N1091), .A1(n236), .B0(SHA256_result[48]), .B1(n11), .Y(
        n1473) );
  AOI22XL U599 ( .A0(N1088), .A1(n236), .B0(SHA256_result[45]), .B1(n10), .Y(
        n1476) );
  AOI22XL U600 ( .A0(N1087), .A1(n236), .B0(SHA256_result[44]), .B1(n10), .Y(
        n1477) );
  AOI22XL U601 ( .A0(N1082), .A1(n235), .B0(SHA256_result[39]), .B1(n10), .Y(
        n1482) );
  AOI22XL U602 ( .A0(N1095), .A1(n236), .B0(SHA256_result[52]), .B1(n11), .Y(
        n1469) );
  AOI22XL U603 ( .A0(N1094), .A1(n236), .B0(SHA256_result[51]), .B1(n11), .Y(
        n1470) );
  AOI22XL U604 ( .A0(N1093), .A1(n236), .B0(SHA256_result[50]), .B1(n11), .Y(
        n1471) );
  AOI22XL U605 ( .A0(N1084), .A1(n236), .B0(SHA256_result[41]), .B1(n10), .Y(
        n1480) );
  AOI22XL U606 ( .A0(N1081), .A1(n235), .B0(SHA256_result[38]), .B1(n10), .Y(
        n1483) );
  NAND2XL U607 ( .A(n108), .B(n196), .Y(n393) );
  AOI21XL U608 ( .A0(SHA256_result[37]), .A1(n212), .B0(n271), .Y(n354) );
  INVXL U609 ( .A(next_E[7]), .Y(n482) );
  INVXL U610 ( .A(next_E[3]), .Y(n498) );
  INVXL U611 ( .A(next_E[2]), .Y(n501) );
  INVXL U612 ( .A(next_E[1]), .Y(n505) );
  INVXL U613 ( .A(next_E[5]), .Y(n490) );
  AOI21XL U614 ( .A0(SHA256_result[101]), .A1(n211), .B0(n272), .Y(n488) );
  INVXL U615 ( .A(next_E[4]), .Y(n494) );
  AOI21XL U616 ( .A0(SHA256_result[100]), .A1(n211), .B0(n274), .Y(n492) );
  AOI21XL U617 ( .A0(n77), .A1(n211), .B0(n272), .Y(n507) );
  AOI21XL U618 ( .A0(SHA256_result[35]), .A1(n211), .B0(n271), .Y(n359) );
  OAI211XL U619 ( .A0(n23), .A1(n106), .B0(n367), .C0(n366), .Y(n2666) );
  AOI21XL U620 ( .A0(n96), .A1(n212), .B0(n271), .Y(n366) );
  AOI21XL U621 ( .A0(SHA256_result[67]), .A1(n212), .B0(n271), .Y(n384) );
  AOI21XL U622 ( .A0(SHA256_result[66]), .A1(n212), .B0(n271), .Y(n386) );
  NAND2XL U623 ( .A(SHA256_result[69]), .B(n196), .Y(n380) );
  NAND2XL U624 ( .A(n90), .B(n197), .Y(n529) );
  NAND2XL U625 ( .A(N916), .B(n247), .Y(n527) );
  AOI21XL U626 ( .A0(n87), .A1(n211), .B0(n272), .Y(n526) );
  NAND2XL U627 ( .A(SHA256_result[36]), .B(n195), .Y(n358) );
  NAND2XL U628 ( .A(N1047), .B(n244), .Y(n357) );
  NAND2XL U629 ( .A(N1022), .B(n245), .Y(n375) );
  AOI21XL U630 ( .A0(n213), .A1(SHA256_result[75]), .B0(n271), .Y(n374) );
  NAND2XL U631 ( .A(N1018), .B(n245), .Y(n377) );
  AOI21XL U632 ( .A0(n213), .A1(SHA256_result[71]), .B0(n271), .Y(n376) );
  NAND2XL U633 ( .A(SHA256_result[68]), .B(n194), .Y(n383) );
  NAND2XL U634 ( .A(N1015), .B(n245), .Y(n382) );
  NAND2XL U635 ( .A(n115), .B(n197), .Y(n390) );
  NAND2XL U636 ( .A(N1012), .B(n245), .Y(n389) );
  NAND2XL U637 ( .A(SHA256_result[163]), .B(n195), .Y(n521) );
  NAND2XL U638 ( .A(N918), .B(n247), .Y(n520) );
  NAND2XL U639 ( .A(SHA256_result[162]), .B(n196), .Y(n525) );
  NAND2XL U640 ( .A(N917), .B(n247), .Y(n524) );
  AOI2BB2XL U641 ( .B0(N883), .B1(n239), .A0N(n13), .A1N(n93), .Y(n541) );
  NOR3XL U642 ( .A(output_enable), .B(round[6]), .C(n1849), .Y(n141) );
  NAND2XL U643 ( .A(output_enable), .B(n1434), .Y(n1975) );
  AOI31XL U644 ( .A0(n329), .A1(n1389), .A2(n2357), .B0(n2407), .Y(n2402) );
  AOI22XL U645 ( .A0(n2260), .A1(n330), .B0(n2382), .B1(n1371), .Y(n2376) );
  AOI221XL U646 ( .A0(n722), .A1(n1384), .B0(n2308), .B1(n183), .C0(n2309), 
        .Y(n2302) );
  AOI2BB2XL U647 ( .B0(n2300), .B1(round[2]), .A0N(n2289), .A1N(n1397), .Y(
        n2290) );
  AOI31XL U648 ( .A0(n2349), .A1(n333), .A2(n2261), .B0(n2313), .Y(n2522) );
  NOR3XL U649 ( .A(n2496), .B(n2271), .C(n2313), .Y(n2488) );
  AOI211XL U650 ( .A0(n2425), .A1(n333), .B0(n2462), .C0(n2463), .Y(n2461) );
  AND3X1 U651 ( .A(n1434), .B(n1337), .C(inner_busy), .Y(n144) );
  NOR3XL U652 ( .A(n1371), .B(round[2]), .C(n140), .Y(n2446) );
  NOR3XL U653 ( .A(n742), .B(n1384), .C(n330), .Y(n2357) );
  NOR3XL U654 ( .A(n1384), .B(n183), .C(n717), .Y(n2263) );
  INVX1 U655 ( .A(n329), .Y(n328) );
  OAI22XL U656 ( .A0(round[3]), .A1(n2304), .B0(n2518), .B1(n1371), .Y(n2517)
         );
  NOR2XL U657 ( .A(n1389), .B(round[3]), .Y(n2262) );
  NOR2XL U658 ( .A(n1371), .B(round[3]), .Y(n2329) );
  AOI222XL U659 ( .A0(n2473), .A1(n1384), .B0(n2425), .B1(n1371), .C0(n2429), 
        .C1(n183), .Y(n2513) );
  AOI22XL U660 ( .A0(n2053), .A1(SHA256_result[200]), .B0(n2054), .B1(
        SHA256_result[204]), .Y(n2221) );
  AOI22XL U661 ( .A0(n2055), .A1(SHA256_result[208]), .B0(n2056), .B1(
        SHA256_result[212]), .Y(n2220) );
  AOI22XL U662 ( .A0(n2063), .A1(SHA256_result[162]), .B0(n2064), .B1(
        SHA256_result[166]), .Y(n2120) );
  AOI22XL U663 ( .A0(n2051), .A1(SHA256_result[194]), .B0(n2052), .B1(
        SHA256_result[198]), .Y(n2116) );
  AOI22XL U664 ( .A0(n2051), .A1(SHA256_result[195]), .B0(n2052), .B1(
        SHA256_result[199]), .Y(n2050) );
  AOI22XL U665 ( .A0(n2053), .A1(SHA256_result[203]), .B0(n2054), .B1(
        SHA256_result[207]), .Y(n2049) );
  AOI22XL U666 ( .A0(n2055), .A1(SHA256_result[211]), .B0(n2056), .B1(
        SHA256_result[215]), .Y(n2048) );
  AOI22XL U667 ( .A0(n2014), .A1(SHA256_result[41]), .B0(n2015), .B1(
        SHA256_result[45]), .Y(n2141) );
  AOI22XL U668 ( .A0(n2053), .A1(SHA256_result[201]), .B0(n2054), .B1(
        SHA256_result[205]), .Y(n2157) );
  AOI22XL U669 ( .A0(n2055), .A1(SHA256_result[209]), .B0(n2056), .B1(
        SHA256_result[213]), .Y(n2156) );
  AOI22XL U670 ( .A0(n2053), .A1(SHA256_result[202]), .B0(n2054), .B1(
        SHA256_result[206]), .Y(n2115) );
  AOI22XL U671 ( .A0(n2055), .A1(SHA256_result[210]), .B0(n2056), .B1(
        SHA256_result[214]), .Y(n2114) );
  AOI22XL U672 ( .A0(n2014), .A1(SHA256_result[40]), .B0(n2015), .B1(
        SHA256_result[44]), .Y(n2195) );
  AOI22XL U673 ( .A0(n2063), .A1(n87), .B0(n2064), .B1(SHA256_result[165]), 
        .Y(n2162) );
  AOI22XL U674 ( .A0(n2063), .A1(SHA256_result[163]), .B0(n2064), .B1(
        SHA256_result[167]), .Y(n2062) );
  AOI22XL U675 ( .A0(n2000), .A1(SHA256_result[67]), .B0(n2001), .B1(
        SHA256_result[71]), .Y(n1999) );
  AOI22XL U676 ( .A0(n2051), .A1(SHA256_result[193]), .B0(n2052), .B1(
        SHA256_result[197]), .Y(n2158) );
  AOI22XL U677 ( .A0(n2000), .A1(SHA256_result[66]), .B0(n2001), .B1(
        SHA256_result[70]), .Y(n2096) );
  AOI22XL U678 ( .A0(n2051), .A1(SHA256_result[192]), .B0(n2052), .B1(
        SHA256_result[196]), .Y(n2222) );
  AOI22XL U679 ( .A0(n2014), .A1(SHA256_result[42]), .B0(n2015), .B1(
        SHA256_result[46]), .Y(n2099) );
  AOI22XL U680 ( .A0(n2014), .A1(SHA256_result[43]), .B0(n2015), .B1(
        SHA256_result[47]), .Y(n2010) );
  AOI22XL U681 ( .A0(n2027), .A1(SHA256_result[16]), .B0(n2028), .B1(
        SHA256_result[20]), .Y(n2202) );
  AOI22XL U682 ( .A0(n2027), .A1(SHA256_result[17]), .B0(n2028), .B1(
        SHA256_result[21]), .Y(n2144) );
  AOI22XL U683 ( .A0(n2027), .A1(SHA256_result[18]), .B0(n2028), .B1(
        SHA256_result[22]), .Y(n2102) );
  AOI22XL U684 ( .A0(n2027), .A1(SHA256_result[19]), .B0(n2028), .B1(
        SHA256_result[23]), .Y(n2021) );
  AOI22XL U685 ( .A0(n2025), .A1(SHA256_result[11]), .B0(n2026), .B1(
        SHA256_result[15]), .Y(n2022) );
  AOI22XL U686 ( .A0(n1977), .A1(SHA256_result[2]), .B0(n2024), .B1(
        SHA256_result[6]), .Y(n2104) );
  AOI22XL U687 ( .A0(n2025), .A1(SHA256_result[8]), .B0(n2026), .B1(
        SHA256_result[12]), .Y(n2203) );
  AOI22XL U688 ( .A0(n2025), .A1(SHA256_result[9]), .B0(n2026), .B1(
        SHA256_result[13]), .Y(n2145) );
  AOI22XL U689 ( .A0(n2025), .A1(SHA256_result[10]), .B0(n2026), .B1(
        SHA256_result[14]), .Y(n2103) );
  AOI22XL U690 ( .A0(n1977), .A1(SHA256_result[0]), .B0(n2024), .B1(
        SHA256_result[4]), .Y(n2204) );
  AOI22XL U691 ( .A0(n1977), .A1(SHA256_result[1]), .B0(n2024), .B1(
        SHA256_result[5]), .Y(n2146) );
  AOI22XL U692 ( .A0(n2000), .A1(n115), .B0(n2001), .B1(SHA256_result[69]), 
        .Y(n2138) );
  AOI22XL U693 ( .A0(n2075), .A1(SHA256_result[130]), .B0(n2076), .B1(
        SHA256_result[134]), .Y(n2124) );
  AOI22XL U694 ( .A0(n2075), .A1(SHA256_result[128]), .B0(n2076), .B1(
        SHA256_result[132]), .Y(n2236) );
  AOI22XL U695 ( .A0(n1977), .A1(SHA256_result[3]), .B0(n2024), .B1(
        SHA256_result[7]), .Y(n2023) );
  AOI22XL U696 ( .A0(n2075), .A1(SHA256_result[129]), .B0(n2076), .B1(
        SHA256_result[133]), .Y(n2166) );
  AOI22XL U697 ( .A0(n2000), .A1(n108), .B0(n2001), .B1(SHA256_result[68]), 
        .Y(n2186) );
  AOI22XL U698 ( .A0(n2075), .A1(SHA256_result[131]), .B0(n2076), .B1(
        SHA256_result[135]), .Y(n2074) );
  AOI22XL U699 ( .A0(n2063), .A1(n90), .B0(n2064), .B1(SHA256_result[164]), 
        .Y(n2228) );
  AOI22XL U700 ( .A0(n1988), .A1(n77), .B0(n1989), .B1(SHA256_result[100]), 
        .Y(n2176) );
  AOI22XL U701 ( .A0(n2016), .A1(SHA256_result[51]), .B0(n2017), .B1(
        SHA256_result[55]), .Y(n2009) );
  AOI22XL U702 ( .A0(n2012), .A1(SHA256_result[35]), .B0(n2013), .B1(
        SHA256_result[39]), .Y(n2011) );
  AOI22XL U703 ( .A0(n2016), .A1(SHA256_result[50]), .B0(n2017), .B1(
        SHA256_result[54]), .Y(n2098) );
  AOI22XL U704 ( .A0(n2012), .A1(SHA256_result[34]), .B0(n2013), .B1(
        SHA256_result[38]), .Y(n2100) );
  AOI22XL U705 ( .A0(n2067), .A1(SHA256_result[178]), .B0(n2068), .B1(
        SHA256_result[182]), .Y(n2118) );
  AOI22XL U706 ( .A0(n2065), .A1(SHA256_result[170]), .B0(n2066), .B1(
        SHA256_result[174]), .Y(n2119) );
  AOI22XL U707 ( .A0(n2067), .A1(SHA256_result[179]), .B0(n2068), .B1(
        SHA256_result[183]), .Y(n2060) );
  AOI22XL U708 ( .A0(n2065), .A1(SHA256_result[171]), .B0(n2066), .B1(
        SHA256_result[175]), .Y(n2061) );
  AOI22XL U709 ( .A0(n1994), .A1(SHA256_result[120]), .B0(n1995), .B1(
        SHA256_result[124]), .Y(n2173) );
  AOI22XL U710 ( .A0(n1992), .A1(SHA256_result[112]), .B0(n1993), .B1(
        SHA256_result[116]), .Y(n2174) );
  AOI22XL U711 ( .A0(n1990), .A1(n153), .B0(n1991), .B1(n150), .Y(n2175) );
  AOI22XL U712 ( .A0(n2004), .A1(SHA256_result[83]), .B0(n2005), .B1(
        SHA256_result[87]), .Y(n1997) );
  AOI22XL U713 ( .A0(n2002), .A1(SHA256_result[75]), .B0(n2003), .B1(
        SHA256_result[79]), .Y(n1998) );
  AOI22XL U714 ( .A0(n2004), .A1(SHA256_result[82]), .B0(n2005), .B1(
        SHA256_result[86]), .Y(n2094) );
  AOI22XL U715 ( .A0(n2002), .A1(SHA256_result[74]), .B0(n2003), .B1(
        SHA256_result[78]), .Y(n2095) );
  AOI22XL U716 ( .A0(n1994), .A1(SHA256_result[122]), .B0(n1995), .B1(n145), 
        .Y(n2089) );
  AOI22XL U717 ( .A0(n1992), .A1(SHA256_result[114]), .B0(n1993), .B1(
        SHA256_result[118]), .Y(n2090) );
  AOI22XL U718 ( .A0(n1990), .A1(n151), .B0(n1991), .B1(SHA256_result[110]), 
        .Y(n2091) );
  AOI22XL U719 ( .A0(n2016), .A1(SHA256_result[48]), .B0(n2017), .B1(
        SHA256_result[52]), .Y(n2194) );
  AOI22XL U720 ( .A0(n2012), .A1(n96), .B0(n2013), .B1(SHA256_result[36]), .Y(
        n2196) );
  AOI22XL U721 ( .A0(n2067), .A1(SHA256_result[176]), .B0(n2068), .B1(
        SHA256_result[180]), .Y(n2226) );
  AOI22XL U722 ( .A0(n2065), .A1(SHA256_result[168]), .B0(n2066), .B1(
        SHA256_result[172]), .Y(n2227) );
  AOI22XL U723 ( .A0(n2067), .A1(SHA256_result[177]), .B0(n2068), .B1(
        SHA256_result[181]), .Y(n2160) );
  AOI22XL U724 ( .A0(n2065), .A1(SHA256_result[169]), .B0(n2066), .B1(
        SHA256_result[173]), .Y(n2161) );
  AOI22XL U725 ( .A0(n1994), .A1(n73), .B0(n1995), .B1(SHA256_result[127]), 
        .Y(n1984) );
  AOI22XL U726 ( .A0(n1992), .A1(n147), .B0(n1993), .B1(SHA256_result[119]), 
        .Y(n1985) );
  AOI22XL U727 ( .A0(n1990), .A1(SHA256_result[107]), .B0(n1991), .B1(n149), 
        .Y(n1986) );
  AOI22XL U728 ( .A0(n1992), .A1(n148), .B0(n1993), .B1(n146), .Y(n2132) );
  AOI22XL U729 ( .A0(n1990), .A1(n152), .B0(n1991), .B1(SHA256_result[109]), 
        .Y(n2133) );
  AOI22XL U730 ( .A0(n2004), .A1(SHA256_result[80]), .B0(n2005), .B1(
        SHA256_result[84]), .Y(n2184) );
  AOI22XL U731 ( .A0(n2002), .A1(SHA256_result[72]), .B0(n2003), .B1(
        SHA256_result[76]), .Y(n2185) );
  AOI22XL U732 ( .A0(n2045), .A1(n160), .B0(n2046), .B1(SHA256_result[252]), 
        .Y(n2211) );
  AOI22XL U733 ( .A0(n2041), .A1(n175), .B0(n2042), .B1(n171), .Y(n2213) );
  AOI22XL U734 ( .A0(n2043), .A1(n167), .B0(n2044), .B1(n163), .Y(n2212) );
  AOI22XL U735 ( .A0(n2045), .A1(n157), .B0(n2046), .B1(SHA256_result[255]), 
        .Y(n2035) );
  AOI22XL U736 ( .A0(n2041), .A1(n172), .B0(n2042), .B1(n168), .Y(n2037) );
  AOI22XL U737 ( .A0(n2043), .A1(n164), .B0(n2044), .B1(n161), .Y(n2036) );
  AOI22XL U738 ( .A0(n2045), .A1(n158), .B0(n2046), .B1(n155), .Y(n2109) );
  AOI22XL U739 ( .A0(n2041), .A1(n173), .B0(n2042), .B1(n169), .Y(n2111) );
  AOI22XL U740 ( .A0(n2043), .A1(n165), .B0(n2044), .B1(n37), .Y(n2110) );
  AOI22XL U741 ( .A0(n2016), .A1(SHA256_result[49]), .B0(n2017), .B1(
        SHA256_result[53]), .Y(n2140) );
  AOI22XL U742 ( .A0(n2012), .A1(SHA256_result[33]), .B0(n2013), .B1(
        SHA256_result[37]), .Y(n2142) );
  AOI22XL U743 ( .A0(n2004), .A1(SHA256_result[81]), .B0(n2005), .B1(
        SHA256_result[85]), .Y(n2136) );
  AOI22XL U744 ( .A0(n2002), .A1(SHA256_result[73]), .B0(n2003), .B1(
        SHA256_result[77]), .Y(n2137) );
  INVXL U745 ( .A(SHA256_result[252]), .Y(n697) );
  INVXL U746 ( .A(SHA256_result[255]), .Y(n700) );
  INVXL U747 ( .A(n73), .Y(n418) );
  INVXL U748 ( .A(SHA256_result[118]), .Y(n861) );
  INVXL U749 ( .A(SHA256_result[121]), .Y(n426) );
  INVXL U750 ( .A(SHA256_result[127]), .Y(n511) );
  INVXL U751 ( .A(n37), .Y(n605) );
  INVXL U752 ( .A(SHA256_result[193]), .Y(n761) );
  INVXL U753 ( .A(SHA256_result[210]), .Y(n778) );
  INVXL U754 ( .A(SHA256_result[209]), .Y(n777) );
  INVXL U755 ( .A(SHA256_result[201]), .Y(n769) );
  INVXL U756 ( .A(SHA256_result[207]), .Y(n775) );
  INVXL U757 ( .A(SHA256_result[205]), .Y(n773) );
  INVXL U758 ( .A(SHA256_result[211]), .Y(n779) );
  INVXL U759 ( .A(SHA256_result[200]), .Y(n768) );
  INVXL U760 ( .A(SHA256_result[206]), .Y(n774) );
  INVXL U761 ( .A(SHA256_result[204]), .Y(n772) );
  INVXL U762 ( .A(SHA256_result[198]), .Y(n766) );
  INVXL U763 ( .A(SHA256_result[197]), .Y(n765) );
  INVXL U764 ( .A(SHA256_result[196]), .Y(n764) );
  INVXL U765 ( .A(SHA256_result[43]), .Y(n895) );
  INVXL U766 ( .A(SHA256_result[40]), .Y(n892) );
  INVXL U767 ( .A(SHA256_result[80]), .Y(n875) );
  INVXL U768 ( .A(SHA256_result[55]), .Y(n907) );
  INVXL U769 ( .A(SHA256_result[47]), .Y(n899) );
  INVXL U770 ( .A(SHA256_result[46]), .Y(n898) );
  INVXL U771 ( .A(SHA256_result[179]), .Y(n806) );
  INVXL U772 ( .A(SHA256_result[178]), .Y(n805) );
  INVXL U773 ( .A(SHA256_result[177]), .Y(n804) );
  INVXL U774 ( .A(SHA256_result[168]), .Y(n795) );
  INVXL U775 ( .A(SHA256_result[78]), .Y(n873) );
  INVXL U776 ( .A(SHA256_result[175]), .Y(n802) );
  INVXL U777 ( .A(SHA256_result[174]), .Y(n801) );
  INVXL U778 ( .A(SHA256_result[173]), .Y(n800) );
  INVXL U779 ( .A(SHA256_result[172]), .Y(n799) );
  INVXL U780 ( .A(SHA256_result[165]), .Y(n792) );
  INVXL U781 ( .A(SHA256_result[164]), .Y(n791) );
  INVXL U782 ( .A(SHA256_result[42]), .Y(n894) );
  INVXL U783 ( .A(SHA256_result[81]), .Y(n876) );
  INVXL U784 ( .A(SHA256_result[72]), .Y(n867) );
  INVXL U785 ( .A(SHA256_result[54]), .Y(n906) );
  INVXL U786 ( .A(SHA256_result[53]), .Y(n905) );
  INVXL U787 ( .A(SHA256_result[176]), .Y(n803) );
  INVXL U788 ( .A(SHA256_result[170]), .Y(n797) );
  INVXL U789 ( .A(SHA256_result[87]), .Y(n882) );
  INVXL U790 ( .A(SHA256_result[79]), .Y(n874) );
  INVXL U791 ( .A(SHA256_result[76]), .Y(n871) );
  INVXL U792 ( .A(SHA256_result[119]), .Y(n862) );
  INVXL U793 ( .A(SHA256_result[120]), .Y(n863) );
  INVXL U794 ( .A(SHA256_result[114]), .Y(n857) );
  INVXL U795 ( .A(SHA256_result[125]), .Y(n410) );
  INVXL U796 ( .A(SHA256_result[208]), .Y(n776) );
  INVXL U797 ( .A(SHA256_result[203]), .Y(n771) );
  INVXL U798 ( .A(SHA256_result[202]), .Y(n770) );
  INVXL U799 ( .A(SHA256_result[199]), .Y(n767) );
  INVXL U800 ( .A(SHA256_result[194]), .Y(n762) );
  INVXL U801 ( .A(SHA256_result[195]), .Y(n763) );
  INVXL U802 ( .A(SHA256_result[71]), .Y(n866) );
  INVXL U803 ( .A(SHA256_result[39]), .Y(n891) );
  INVXL U804 ( .A(SHA256_result[75]), .Y(n870) );
  INVXL U805 ( .A(SHA256_result[49]), .Y(n901) );
  INVXL U806 ( .A(SHA256_result[48]), .Y(n900) );
  INVXL U807 ( .A(SHA256_result[82]), .Y(n877) );
  INVXL U808 ( .A(SHA256_result[169]), .Y(n796) );
  INVXL U809 ( .A(SHA256_result[44]), .Y(n896) );
  INVXL U810 ( .A(SHA256_result[77]), .Y(n872) );
  INVXL U811 ( .A(SHA256_result[166]), .Y(n793) );
  INVXL U812 ( .A(SHA256_result[51]), .Y(n903) );
  INVXL U813 ( .A(SHA256_result[50]), .Y(n902) );
  INVXL U814 ( .A(SHA256_result[41]), .Y(n893) );
  INVXL U815 ( .A(SHA256_result[83]), .Y(n878) );
  INVXL U816 ( .A(SHA256_result[74]), .Y(n869) );
  INVXL U817 ( .A(SHA256_result[73]), .Y(n868) );
  INVXL U818 ( .A(SHA256_result[171]), .Y(n798) );
  INVXL U819 ( .A(SHA256_result[52]), .Y(n904) );
  INVXL U820 ( .A(SHA256_result[45]), .Y(n897) );
  INVXL U821 ( .A(SHA256_result[38]), .Y(n890) );
  INVXL U822 ( .A(SHA256_result[86]), .Y(n881) );
  INVXL U823 ( .A(SHA256_result[85]), .Y(n880) );
  INVXL U824 ( .A(SHA256_result[84]), .Y(n879) );
  INVXL U825 ( .A(SHA256_result[70]), .Y(n865) );
  INVXL U826 ( .A(SHA256_result[167]), .Y(n794) );
  INVXL U827 ( .A(SHA256_result[2]), .Y(n919) );
  NOR2XL U828 ( .A(n329), .B(n1384), .Y(n2457) );
  INVXL U829 ( .A(SHA256_result[11]), .Y(n928) );
  INVXL U830 ( .A(SHA256_result[131]), .Y(n823) );
  INVXL U831 ( .A(SHA256_result[129]), .Y(n821) );
  INVXL U832 ( .A(SHA256_result[21]), .Y(n938) );
  INVXL U833 ( .A(SHA256_result[1]), .Y(n918) );
  INVXL U834 ( .A(SHA256_result[10]), .Y(n927) );
  INVXL U835 ( .A(SHA256_result[8]), .Y(n925) );
  INVXL U836 ( .A(SHA256_result[23]), .Y(n940) );
  INVXL U837 ( .A(SHA256_result[22]), .Y(n939) );
  INVXL U838 ( .A(SHA256_result[15]), .Y(n932) );
  INVXL U839 ( .A(SHA256_result[14]), .Y(n931) );
  INVXL U840 ( .A(SHA256_result[5]), .Y(n922) );
  INVXL U841 ( .A(SHA256_result[17]), .Y(n934) );
  INVXL U842 ( .A(SHA256_result[16]), .Y(n933) );
  INVXL U843 ( .A(SHA256_result[20]), .Y(n937) );
  INVXL U844 ( .A(SHA256_result[13]), .Y(n930) );
  INVXL U845 ( .A(SHA256_result[12]), .Y(n929) );
  INVXL U846 ( .A(SHA256_result[7]), .Y(n924) );
  INVXL U847 ( .A(SHA256_result[19]), .Y(n936) );
  INVXL U848 ( .A(SHA256_result[18]), .Y(n935) );
  INVXL U849 ( .A(SHA256_result[9]), .Y(n926) );
  INVXL U850 ( .A(SHA256_result[130]), .Y(n822) );
  INVXL U851 ( .A(SHA256_result[128]), .Y(n820) );
  INVXL U852 ( .A(SHA256_result[6]), .Y(n923) );
  INVXL U853 ( .A(SHA256_result[0]), .Y(n917) );
  INVXL U854 ( .A(SHA256_result[3]), .Y(n920) );
  INVXL U855 ( .A(SHA256_result[4]), .Y(n921) );
  INVXL U856 ( .A(SHA256_result[163]), .Y(n519) );
  INVXL U857 ( .A(SHA256_result[122]), .Y(n422) );
  INVXL U858 ( .A(SHA256_result[101]), .Y(n487) );
  INVXL U859 ( .A(SHA256_result[100]), .Y(n491) );
  INVXL U860 ( .A(n77), .Y(n506) );
  INVXL U861 ( .A(SHA256_result[124]), .Y(n413) );
  INVXL U862 ( .A(SHA256_result[110]), .Y(n853) );
  INVXL U863 ( .A(SHA256_result[112]), .Y(n855) );
  INVXL U864 ( .A(SHA256_result[109]), .Y(n852) );
  INVXL U865 ( .A(SHA256_result[107]), .Y(n461) );
  INVXL U866 ( .A(SHA256_result[192]), .Y(n760) );
  AOI22XL U867 ( .A0(n1994), .A1(SHA256_result[121]), .B0(n1995), .B1(
        SHA256_result[125]), .Y(n2131) );
  INVX1 U868 ( .A(n299), .Y(n291) );
  INVX1 U869 ( .A(n217), .Y(n211) );
  INVX1 U870 ( .A(n217), .Y(n212) );
  INVX1 U871 ( .A(n209), .Y(n214) );
  INVX1 U872 ( .A(n199), .Y(n191) );
  INVX1 U873 ( .A(n197), .Y(n186) );
  INVX1 U874 ( .A(n198), .Y(n189) );
  INVX1 U875 ( .A(n198), .Y(n188) );
  INVX1 U876 ( .A(n199), .Y(n190) );
  INVX1 U877 ( .A(n197), .Y(n187) );
  INVX1 U878 ( .A(n279), .Y(n274) );
  INVX1 U879 ( .A(n279), .Y(n276) );
  INVX1 U880 ( .A(n279), .Y(n277) );
  INVX1 U881 ( .A(n270), .Y(n272) );
  INVX1 U882 ( .A(n312), .Y(n300) );
  INVX1 U883 ( .A(n313), .Y(n298) );
  INVX1 U884 ( .A(n313), .Y(n297) );
  INVX1 U885 ( .A(n313), .Y(n296) );
  INVX1 U886 ( .A(n204), .Y(n216) );
  INVX1 U887 ( .A(n204), .Y(n217) );
  INVX1 U888 ( .A(n266), .Y(n255) );
  INVX1 U889 ( .A(n266), .Y(n256) );
  INVX1 U890 ( .A(n251), .Y(n258) );
  INVX1 U891 ( .A(n251), .Y(n257) );
  INVX1 U892 ( .A(n266), .Y(n254) );
  INVX1 U893 ( .A(n266), .Y(n253) );
  INVX1 U894 ( .A(n266), .Y(n259) );
  INVX1 U895 ( .A(n251), .Y(n260) );
  INVX1 U896 ( .A(n266), .Y(n252) );
  INVX1 U897 ( .A(n208), .Y(n233) );
  INVX1 U898 ( .A(n207), .Y(n230) );
  INVX1 U899 ( .A(n207), .Y(n231) );
  INVX1 U900 ( .A(n208), .Y(n232) );
  INVX1 U901 ( .A(n206), .Y(n225) );
  INVX1 U902 ( .A(n206), .Y(n227) );
  INVX1 U903 ( .A(n207), .Y(n228) );
  INVX1 U904 ( .A(n205), .Y(n229) );
  INVX1 U905 ( .A(n205), .Y(n220) );
  INVX1 U906 ( .A(n205), .Y(n221) );
  INVX1 U907 ( .A(n206), .Y(n222) );
  INVX1 U908 ( .A(n206), .Y(n224) );
  INVX1 U909 ( .A(n206), .Y(n226) );
  INVX1 U910 ( .A(n205), .Y(n218) );
  INVX1 U911 ( .A(n207), .Y(n219) );
  INVX1 U912 ( .A(n206), .Y(n223) );
  INVX1 U913 ( .A(n208), .Y(n215) );
  INVX1 U914 ( .A(n675), .Y(n236) );
  INVX1 U915 ( .A(n675), .Y(n239) );
  INVX1 U916 ( .A(n249), .Y(n243) );
  INVX1 U917 ( .A(n250), .Y(n240) );
  INVX1 U918 ( .A(n250), .Y(n242) );
  INVX1 U919 ( .A(n249), .Y(n241) );
  INVX1 U920 ( .A(n675), .Y(n245) );
  INVX1 U921 ( .A(n675), .Y(n247) );
  INVX1 U922 ( .A(n675), .Y(n248) );
  INVX1 U923 ( .A(n675), .Y(n246) );
  INVX1 U924 ( .A(n326), .Y(n318) );
  INVX1 U925 ( .A(n326), .Y(n319) );
  INVX1 U926 ( .A(n325), .Y(n320) );
  INVX1 U927 ( .A(n325), .Y(n321) );
  INVX1 U928 ( .A(n325), .Y(n322) );
  INVX1 U929 ( .A(n326), .Y(n323) );
  INVX1 U930 ( .A(n270), .Y(n271) );
  INVX1 U931 ( .A(n287), .Y(n301) );
  INVX1 U932 ( .A(n283), .Y(n312) );
  INVX1 U933 ( .A(n281), .Y(n308) );
  INVX1 U934 ( .A(n281), .Y(n307) );
  INVX1 U935 ( .A(n281), .Y(n309) );
  INVX1 U936 ( .A(n280), .Y(n306) );
  INVX1 U937 ( .A(n280), .Y(n305) );
  INVX1 U938 ( .A(n280), .Y(n304) );
  INVX1 U939 ( .A(n282), .Y(n310) );
  INVX1 U940 ( .A(n282), .Y(n303) );
  INVX1 U941 ( .A(n282), .Y(n311) );
  INVX1 U942 ( .A(n138), .Y(n279) );
  INVX1 U943 ( .A(n201), .Y(n197) );
  INVX1 U944 ( .A(n266), .Y(n264) );
  INVX1 U945 ( .A(n266), .Y(n263) );
  INVX1 U946 ( .A(n266), .Y(n265) );
  INVX1 U947 ( .A(n267), .Y(n262) );
  INVX1 U948 ( .A(n208), .Y(n234) );
  INVX1 U949 ( .A(n203), .Y(n192) );
  INVX1 U950 ( .A(n202), .Y(n193) );
  INVX1 U951 ( .A(n203), .Y(n194) );
  INVX1 U952 ( .A(n202), .Y(n195) );
  INVX1 U953 ( .A(n209), .Y(n207) );
  INVX1 U954 ( .A(n209), .Y(n208) );
  INVX1 U955 ( .A(n209), .Y(n205) );
  INVX1 U956 ( .A(n209), .Y(n206) );
  INVX1 U957 ( .A(n679), .Y(n267) );
  INVX1 U958 ( .A(n282), .Y(n314) );
  INVX1 U959 ( .A(n184), .Y(n200) );
  INVX1 U960 ( .A(n301), .Y(n302) );
  INVX1 U961 ( .A(n196), .Y(n202) );
  INVX1 U962 ( .A(n184), .Y(n201) );
  INVX1 U963 ( .A(n674), .Y(n210) );
  INVX1 U964 ( .A(n678), .Y(n250) );
  INVX1 U965 ( .A(n678), .Y(n249) );
  INVX1 U966 ( .A(n284), .Y(n283) );
  INVX1 U967 ( .A(n285), .Y(n281) );
  INVX1 U968 ( .A(n286), .Y(n280) );
  INVX1 U969 ( .A(n284), .Y(n282) );
  INVX1 U970 ( .A(n198), .Y(n203) );
  INVX1 U971 ( .A(n674), .Y(n209) );
  INVX1 U972 ( .A(n2382), .Y(n710) );
  INVX1 U973 ( .A(n2448), .Y(n751) );
  INVX1 U974 ( .A(n2332), .Y(n746) );
  INVX1 U975 ( .A(n2400), .Y(n729) );
  NOR2X1 U976 ( .A(n730), .B(n749), .Y(n2313) );
  INVX1 U977 ( .A(n2372), .Y(n739) );
  NOR2X1 U978 ( .A(n756), .B(n752), .Y(n2285) );
  INVX1 U979 ( .A(n2257), .Y(n756) );
  INVX1 U980 ( .A(n2406), .Y(n716) );
  NAND4X1 U981 ( .A(n751), .B(n716), .C(n2322), .D(n727), .Y(n2365) );
  NAND2X1 U982 ( .A(n2389), .B(n140), .Y(n2323) );
  INVX1 U983 ( .A(n2399), .Y(n735) );
  AOI21X1 U984 ( .A0(n752), .A1(n719), .B0(n758), .Y(n2485) );
  INVX1 U985 ( .A(n2519), .Y(n708) );
  INVX1 U986 ( .A(n2347), .Y(n732) );
  NAND2X1 U987 ( .A(n725), .B(n717), .Y(n2374) );
  INVX1 U988 ( .A(n2429), .Y(n713) );
  INVX1 U989 ( .A(n2298), .Y(n707) );
  NAND2X1 U990 ( .A(n733), .B(n729), .Y(n2361) );
  NAND2X1 U991 ( .A(n726), .B(n756), .Y(n2398) );
  NOR2X1 U992 ( .A(n191), .B(n601), .Y(n602) );
  OAI2BB1X1 U993 ( .A0N(N877), .A1N(n246), .B0(n591), .Y(n2992) );
  NOR2X1 U994 ( .A(n191), .B(n589), .Y(n590) );
  AOI21XL U995 ( .A0(next_A[24]), .A1(n10), .B0(n598), .Y(n599) );
  INVX1 U996 ( .A(n138), .Y(n270) );
  INVX1 U997 ( .A(n2501), .Y(n758) );
  INVX1 U998 ( .A(n2271), .Y(n753) );
  NAND3X1 U999 ( .A(n330), .B(n333), .C(n1878), .Y(n1859) );
  AOI31X1 U1000 ( .A0(n2421), .A1(n2422), .A2(n2423), .B0(n268), .Y(N3017) );
  NOR3X1 U1001 ( .A(n2426), .B(n2342), .C(n2416), .Y(n2422) );
  AOI211X1 U1002 ( .A0(n2372), .A1(n1397), .B0(n2424), .C0(n2405), .Y(n2423)
         );
  AOI31X1 U1003 ( .A0(n724), .A1(n748), .A2(n2237), .B0(n268), .Y(N3033) );
  INVX1 U1004 ( .A(n2239), .Y(n748) );
  INVX1 U1005 ( .A(n2240), .Y(n724) );
  AND4X2 U1006 ( .A(n750), .B(n720), .C(n739), .D(n740), .Y(n2237) );
  NOR2X1 U1007 ( .A(n749), .B(n755), .Y(n2332) );
  NOR2X1 U1008 ( .A(n757), .B(n752), .Y(n2448) );
  NOR2X1 U1009 ( .A(n711), .B(n332), .Y(n2382) );
  NOR2X1 U1010 ( .A(n730), .B(n755), .Y(n2400) );
  OAI21XL U1011 ( .A0(n335), .A1(n710), .B0(n2495), .Y(n2509) );
  NAND4X1 U1012 ( .A(n2386), .B(n706), .C(n739), .D(n720), .Y(n2443) );
  INVX1 U1013 ( .A(n2445), .Y(n720) );
  NAND3BX1 U1014 ( .AN(n2297), .B(n710), .C(n706), .Y(n2293) );
  INVX1 U1015 ( .A(n2465), .Y(n711) );
  AOI21X1 U1016 ( .A0(n710), .A1(n2269), .B0(n330), .Y(n2359) );
  INVX1 U1017 ( .A(n2258), .Y(n717) );
  NOR2X1 U1018 ( .A(n744), .B(n717), .Y(n2406) );
  NOR2X1 U1019 ( .A(n747), .B(n730), .Y(n2300) );
  INVX1 U1020 ( .A(n2428), .Y(n749) );
  NOR2X1 U1021 ( .A(n757), .B(n742), .Y(n2297) );
  NOR2X1 U1022 ( .A(n742), .B(n755), .Y(n2372) );
  OAI222XL U1023 ( .A0(n742), .A1(n725), .B0(n757), .B1(n707), .C0(n335), .C1(
        n2288), .Y(n2424) );
  NOR3X1 U1024 ( .A(n330), .B(n752), .C(n754), .Y(n2274) );
  NAND2X1 U1025 ( .A(n2521), .B(n335), .Y(n2289) );
  INVX1 U1026 ( .A(n2343), .Y(n725) );
  NOR2X1 U1027 ( .A(n140), .B(n332), .Y(n2298) );
  NOR2X1 U1028 ( .A(n749), .B(n335), .Y(n2473) );
  NOR2X1 U1029 ( .A(n754), .B(n717), .Y(n2306) );
  OAI22X1 U1030 ( .A0(n335), .A1(n757), .B0(n730), .B1(n754), .Y(n2479) );
  NOR2X1 U1031 ( .A(n726), .B(n755), .Y(n2370) );
  NOR2X1 U1032 ( .A(n2456), .B(n335), .Y(n2347) );
  NOR2X1 U1033 ( .A(n730), .B(n757), .Y(n2342) );
  NOR2X1 U1034 ( .A(n754), .B(n738), .Y(n2389) );
  NAND2X1 U1035 ( .A(n2372), .B(n335), .Y(n2322) );
  INVX1 U1036 ( .A(n2435), .Y(n750) );
  NOR2X1 U1037 ( .A(n738), .B(n755), .Y(n2284) );
  INVX1 U1038 ( .A(n131), .Y(n752) );
  INVX1 U1039 ( .A(n2495), .Y(n743) );
  NOR2X1 U1040 ( .A(n717), .B(n755), .Y(n2429) );
  NOR4BBX1 U1041 ( .AN(n2282), .BN(n2386), .C(n2348), .D(n2406), .Y(n2536) );
  AOI31X1 U1042 ( .A0(n734), .A1(n753), .A2(n2255), .B0(n335), .Y(n2254) );
  INVX1 U1043 ( .A(n2437), .Y(n733) );
  OAI22X1 U1044 ( .A0(n332), .A1(n2272), .B0(n757), .B1(n712), .Y(n2469) );
  INVX1 U1045 ( .A(n1878), .Y(n731) );
  INVX1 U1046 ( .A(n2375), .Y(n719) );
  NOR2X1 U1047 ( .A(n738), .B(n758), .Y(n2399) );
  NAND3X1 U1048 ( .A(n731), .B(n732), .C(n714), .Y(n2483) );
  INVX1 U1049 ( .A(n2371), .Y(n718) );
  NOR2X1 U1050 ( .A(n757), .B(n330), .Y(n2257) );
  AOI21X1 U1051 ( .A0(n2282), .A1(n735), .B0(n335), .Y(n2415) );
  INVX1 U1052 ( .A(n2417), .Y(n727) );
  INVX1 U1053 ( .A(n2381), .Y(n712) );
  NAND2X1 U1054 ( .A(n2318), .B(n2261), .Y(n2333) );
  NAND3X1 U1055 ( .A(n2322), .B(n727), .C(n2386), .Y(n2414) );
  NAND3X1 U1056 ( .A(n2307), .B(n714), .C(n713), .Y(n2499) );
  NAND3X1 U1057 ( .A(n2307), .B(n740), .C(n2255), .Y(n2305) );
  AOI21X1 U1058 ( .A0(n739), .A1(n751), .B0(n335), .Y(n2471) );
  AOI21X1 U1059 ( .A0(n2279), .A1(n751), .B0(n1397), .Y(n2320) );
  NAND2X1 U1060 ( .A(n335), .B(n1878), .Y(n2356) );
  NAND3X1 U1061 ( .A(n732), .B(n740), .C(n2356), .Y(n2353) );
  AOI21X1 U1062 ( .A0(n706), .A1(n731), .B0(n332), .Y(n2419) );
  OAI21XL U1063 ( .A0(n129), .A1(n738), .B0(n718), .Y(n2358) );
  OAI2BB1X1 U1064 ( .A0N(n130), .A1N(n2260), .B0(n2456), .Y(n2503) );
  NAND3X1 U1065 ( .A(n2307), .B(n2282), .C(n2272), .Y(n2330) );
  INVX1 U1066 ( .A(n2312), .Y(n737) );
  NAND2X1 U1067 ( .A(n2465), .B(n2428), .Y(n2283) );
  OAI2BB1X1 U1068 ( .A0N(n330), .A1N(n2389), .B0(n714), .Y(n2444) );
  INVX1 U1069 ( .A(n129), .Y(n726) );
  INVX1 U1070 ( .A(n2344), .Y(n715) );
  NOR2X1 U1071 ( .A(n332), .B(n758), .Y(n2427) );
  NOR3X1 U1072 ( .A(n742), .B(n758), .C(n330), .Y(n2275) );
  NAND2X1 U1073 ( .A(n2258), .B(n131), .Y(n2304) );
  INVX1 U1074 ( .A(n2346), .Y(n722) );
  NAND2X1 U1075 ( .A(n738), .B(n752), .Y(n2245) );
  INVX1 U1076 ( .A(n2310), .Y(n721) );
  AOI31X1 U1077 ( .A0(n338), .A1(n341), .A2(n339), .B0(n1849), .Y(n679) );
  OAI221XL U1078 ( .A0(n27), .A1(n912), .B0(n1457), .B1(n945), .C0(n1461), .Y(
        n2574) );
  AOI21X1 U1079 ( .A0(N1103), .A1(n244), .B0(n273), .Y(n1461) );
  OAI221XL U1080 ( .A0(n17), .A1(n698), .B0(n223), .B1(n789), .C0(n1757), .Y(
        n2925) );
  AOI21X1 U1081 ( .A0(N912), .A1(n241), .B0(n278), .Y(n1757) );
  OAI221XL U1082 ( .A0(n14), .A1(n697), .B0(n223), .B1(n788), .C0(n1758), .Y(
        n2926) );
  AOI21X1 U1083 ( .A0(N911), .A1(n241), .B0(n278), .Y(n1758) );
  OAI221XL U1084 ( .A0(n27), .A1(n789), .B0(n228), .B1(n816), .C0(n1725), .Y(
        n2892) );
  AOI21X1 U1085 ( .A0(N944), .A1(n240), .B0(n276), .Y(n1725) );
  OAI221XL U1086 ( .A0(n16), .A1(n887), .B0(n233), .B1(n912), .C0(n1496), .Y(
        n2606) );
  AOI21X1 U1087 ( .A0(N1071), .A1(n243), .B0(n278), .Y(n1496) );
  OAI221XL U1088 ( .A0(n29), .A1(n788), .B0(n228), .B1(n815), .C0(n1726), .Y(
        n2893) );
  AOI21X1 U1089 ( .A0(N943), .A1(n239), .B0(n276), .Y(n1726) );
  OAI221XL U1090 ( .A0(n13), .A1(n816), .B0(n233), .B1(n849), .C0(n1693), .Y(
        n2860) );
  AOI21X1 U1091 ( .A0(N976), .A1(n240), .B0(n275), .Y(n1693) );
  OAI211X1 U1092 ( .A0(n34), .A1(n624), .B0(n623), .C0(n622), .Y(n3003) );
  OAI211X1 U1093 ( .A0(n32), .A1(n621), .B0(n620), .C0(n619), .Y(n3002) );
  INVXL U1094 ( .A(next_A[16]), .Y(n621) );
  AOI21X1 U1095 ( .A0(n213), .A1(n167), .B0(n272), .Y(n620) );
  NAND2X1 U1096 ( .A(N867), .B(n248), .Y(n619) );
  INVXL U1097 ( .A(next_A[19]), .Y(n614) );
  OAI211X1 U1098 ( .A0(n35), .A1(n627), .B0(n626), .C0(n625), .Y(n3004) );
  INVXL U1099 ( .A(next_A[14]), .Y(n627) );
  XOR3X2 U1100 ( .A(n179), .B(n168), .C(n160), .Y(f3_A_32[2]) );
  NAND3X1 U1101 ( .A(n595), .B(n594), .C(n593), .Y(n2993) );
  NAND2X1 U1102 ( .A(N876), .B(n248), .Y(n593) );
  NAND2XL U1103 ( .A(n10), .B(next_E[30]), .Y(n407) );
  NOR2X1 U1104 ( .A(n862), .B(n203), .Y(n432) );
  NOR2X1 U1105 ( .A(n191), .B(n410), .Y(n411) );
  OAI2BB1X1 U1106 ( .A0N(N1004), .A1N(n247), .B0(n428), .Y(n2832) );
  NOR2X1 U1107 ( .A(n697), .B(n191), .Y(n583) );
  INVXL U1108 ( .A(next_E[19]), .Y(n442) );
  OAI211X1 U1109 ( .A0(n28), .A1(n448), .B0(n447), .C0(n446), .Y(n2840) );
  INVXL U1110 ( .A(next_E[17]), .Y(n448) );
  AOI21XL U1111 ( .A0(next_E[27]), .A1(n11), .B0(n419), .Y(n420) );
  NOR2X1 U1112 ( .A(n191), .B(n418), .Y(n419) );
  OAI2BB1X1 U1113 ( .A0N(N869), .A1N(n236), .B0(n616), .Y(n3000) );
  AOI2BB2X1 U1114 ( .B0(n192), .B1(n165), .A0N(n21), .A1N(n615), .Y(n616) );
  INVXL U1115 ( .A(next_A[18]), .Y(n615) );
  OAI2BB1X1 U1116 ( .A0N(N1000), .A1N(n247), .B0(n437), .Y(n2836) );
  AOI2BB2X1 U1117 ( .B0(n193), .B1(n146), .A0N(n23), .A1N(n436), .Y(n437) );
  INVXL U1118 ( .A(next_E[21]), .Y(n436) );
  OAI2BB1X1 U1119 ( .A0N(N872), .A1N(n235), .B0(n609), .Y(n2997) );
  AOI2BB2X1 U1120 ( .B0(n192), .B1(n162), .A0N(n20), .A1N(n608), .Y(n609) );
  INVXL U1121 ( .A(next_A[21]), .Y(n608) );
  OAI2BB1X1 U1122 ( .A0N(N873), .A1N(n236), .B0(n607), .Y(n2996) );
  AOI21XL U1123 ( .A0(next_A[22]), .A1(n10), .B0(n606), .Y(n607) );
  NOR2X1 U1124 ( .A(n700), .B(n203), .Y(n575) );
  NOR2X1 U1125 ( .A(n191), .B(n511), .Y(n512) );
  OAI2BB1X1 U1126 ( .A0N(N871), .A1N(n238), .B0(n611), .Y(n2998) );
  AOI2BB2X1 U1127 ( .B0(n192), .B1(n163), .A0N(n19), .A1N(n610), .Y(n611) );
  INVXL U1128 ( .A(next_A[20]), .Y(n610) );
  OAI2BB1X1 U1129 ( .A0N(N999), .A1N(n245), .B0(n439), .Y(n2837) );
  AOI2BB2X1 U1130 ( .B0(n193), .B1(SHA256_result[116]), .A0N(n36), .A1N(n438), 
        .Y(n439) );
  INVXL U1131 ( .A(next_E[20]), .Y(n438) );
  OAI2BB1X1 U1132 ( .A0N(N868), .A1N(n247), .B0(n618), .Y(n3001) );
  AOI2BB2X1 U1133 ( .B0(n192), .B1(n166), .A0N(n15), .A1N(n617), .Y(n618) );
  INVXL U1134 ( .A(next_A[17]), .Y(n617) );
  OAI2BB1X1 U1135 ( .A0N(N1001), .A1N(n247), .B0(n435), .Y(n2835) );
  AOI21XL U1136 ( .A0(next_E[22]), .A1(n11), .B0(n434), .Y(n435) );
  NOR2X1 U1137 ( .A(n861), .B(n202), .Y(n434) );
  INVX1 U1138 ( .A(output_enable), .Y(n338) );
  OAI221XL U1139 ( .A0(n35), .A1(n644), .B0(n675), .B1(n643), .C0(n642), .Y(
        n3010) );
  NAND2X1 U1140 ( .A(n194), .B(n175), .Y(n642) );
  INVX1 U1141 ( .A(N859), .Y(n643) );
  INVX1 U1142 ( .A(N858), .Y(n646) );
  NAND2X1 U1143 ( .A(n194), .B(n176), .Y(n645) );
  OAI221XL U1144 ( .A0(n35), .A1(n911), .B0(n1457), .B1(n944), .C0(n1462), .Y(
        n2575) );
  AOI21X1 U1145 ( .A0(N1102), .A1(n244), .B0(n273), .Y(n1462) );
  OAI221XL U1146 ( .A0(n30), .A1(n909), .B0(n1457), .B1(n942), .C0(n1464), .Y(
        n2577) );
  AOI21X1 U1147 ( .A0(N1100), .A1(n244), .B0(n273), .Y(n1464) );
  OAI221XL U1148 ( .A0(n33), .A1(n908), .B0(n1457), .B1(n941), .C0(n1465), .Y(
        n2578) );
  AOI21X1 U1149 ( .A0(N1099), .A1(n244), .B0(n273), .Y(n1465) );
  OAI221XL U1150 ( .A0(n30), .A1(n907), .B0(n1457), .B1(n940), .C0(n1466), .Y(
        n2579) );
  OAI221XL U1151 ( .A0(n24), .A1(n906), .B0(n1457), .B1(n939), .C0(n1467), .Y(
        n2580) );
  OAI221XL U1152 ( .A0(n32), .A1(n905), .B0(n1457), .B1(n938), .C0(n1468), .Y(
        n2581) );
  OAI221XL U1153 ( .A0(n17), .A1(n899), .B0(n1457), .B1(n932), .C0(n1474), .Y(
        n2587) );
  AOI21X1 U1154 ( .A0(N1090), .A1(n244), .B0(n276), .Y(n1474) );
  OAI221XL U1155 ( .A0(n31), .A1(n898), .B0(n1457), .B1(n931), .C0(n1475), .Y(
        n2588) );
  OAI221XL U1156 ( .A0(n16), .A1(n895), .B0(n1457), .B1(n928), .C0(n1478), .Y(
        n2591) );
  AOI21X1 U1157 ( .A0(N1086), .A1(n244), .B0(n271), .Y(n1478) );
  OAI221XL U1158 ( .A0(n36), .A1(n894), .B0(n1457), .B1(n927), .C0(n1479), .Y(
        n2592) );
  OAI221XL U1159 ( .A0(n18), .A1(n892), .B0(n1457), .B1(n925), .C0(n1481), .Y(
        n2594) );
  OAI221XL U1160 ( .A0(n18), .A1(n696), .B0(n224), .B1(n787), .C0(n1759), .Y(
        n2927) );
  AOI21X1 U1161 ( .A0(N910), .A1(n241), .B0(n278), .Y(n1759) );
  OAI221XL U1162 ( .A0(n29), .A1(n692), .B0(n225), .B1(n778), .C0(n1768), .Y(
        n2936) );
  OAI221XL U1163 ( .A0(n15), .A1(n691), .B0(n227), .B1(n777), .C0(n1769), .Y(
        n2937) );
  OAI221XL U1164 ( .A0(n23), .A1(n683), .B0(n219), .B1(n769), .C0(n1777), .Y(
        n2945) );
  AOI21X1 U1165 ( .A0(N892), .A1(n242), .B0(n271), .Y(n1777) );
  OAI221XL U1166 ( .A0(n16), .A1(n695), .B0(n226), .B1(n781), .C0(n1765), .Y(
        n2933) );
  AOI21X1 U1167 ( .A0(N904), .A1(n241), .B0(n278), .Y(n1765) );
  OAI221XL U1168 ( .A0(n32), .A1(n689), .B0(n219), .B1(n775), .C0(n1771), .Y(
        n2939) );
  OAI221XL U1169 ( .A0(n21), .A1(n687), .B0(n218), .B1(n773), .C0(n1773), .Y(
        n2941) );
  AOI21X1 U1170 ( .A0(N896), .A1(n242), .B0(n278), .Y(n1773) );
  OAI221XL U1171 ( .A0(n23), .A1(n786), .B0(n228), .B1(n813), .C0(n1728), .Y(
        n2895) );
  AOI21X1 U1172 ( .A0(N941), .A1(n240), .B0(n276), .Y(n1728) );
  OAI221XL U1173 ( .A0(n20), .A1(n779), .B0(n220), .B1(n806), .C0(n1735), .Y(
        n2902) );
  OAI221XL U1174 ( .A0(n22), .A1(n778), .B0(n220), .B1(n805), .C0(n1736), .Y(
        n2903) );
  OAI221XL U1175 ( .A0(n29), .A1(n777), .B0(n220), .B1(n804), .C0(n1737), .Y(
        n2904) );
  OAI221XL U1176 ( .A0(n29), .A1(n768), .B0(n221), .B1(n795), .C0(n1746), .Y(
        n2913) );
  AOI21X1 U1177 ( .A0(N923), .A1(n241), .B0(n277), .Y(n1746) );
  OAI221XL U1178 ( .A0(n36), .A1(n782), .B0(n229), .B1(n809), .C0(n1732), .Y(
        n2899) );
  AOI21X1 U1179 ( .A0(N937), .A1(n235), .B0(n277), .Y(n1732) );
  OAI221XL U1180 ( .A0(n19), .A1(n775), .B0(n220), .B1(n802), .C0(n1739), .Y(
        n2906) );
  OAI221XL U1181 ( .A0(n17), .A1(n774), .B0(n232), .B1(n801), .C0(n1740), .Y(
        n2907) );
  OAI221XL U1182 ( .A0(n32), .A1(n773), .B0(n220), .B1(n800), .C0(n1741), .Y(
        n2908) );
  AOI21X1 U1183 ( .A0(N928), .A1(n241), .B0(n277), .Y(n1741) );
  OAI221XL U1184 ( .A0(n24), .A1(n772), .B0(n221), .B1(n799), .C0(n1742), .Y(
        n2909) );
  AOI21X1 U1185 ( .A0(N927), .A1(n242), .B0(n277), .Y(n1742) );
  OAI221XL U1186 ( .A0(n32), .A1(n765), .B0(n222), .B1(n792), .C0(n1749), .Y(
        n2916) );
  AOI21X1 U1187 ( .A0(N920), .A1(n241), .B0(n278), .Y(n1749) );
  OAI221XL U1188 ( .A0(n34), .A1(n764), .B0(n222), .B1(n791), .C0(n1750), .Y(
        n2917) );
  AOI21X1 U1189 ( .A0(N919), .A1(n242), .B0(n278), .Y(n1750) );
  OAI221XL U1190 ( .A0(n24), .A1(n886), .B0(n233), .B1(n911), .C0(n1497), .Y(
        n2607) );
  AOI21X1 U1191 ( .A0(N1070), .A1(n243), .B0(n275), .Y(n1497) );
  OAI221XL U1192 ( .A0(n33), .A1(n884), .B0(n234), .B1(n909), .C0(n1499), .Y(
        n2609) );
  AOI21X1 U1193 ( .A0(N1068), .A1(n243), .B0(n272), .Y(n1499) );
  OAI221XL U1194 ( .A0(n34), .A1(n883), .B0(n234), .B1(n908), .C0(n1500), .Y(
        n2610) );
  AOI21X1 U1195 ( .A0(N1067), .A1(n243), .B0(n274), .Y(n1500) );
  OAI221XL U1196 ( .A0(n12), .A1(n870), .B0(n230), .B1(n895), .C0(n1513), .Y(
        n2623) );
  OAI221XL U1197 ( .A0(n19), .A1(n867), .B0(n231), .B1(n892), .C0(n1516), .Y(
        n2626) );
  OAI221XL U1198 ( .A0(n15), .A1(n882), .B0(n234), .B1(n907), .C0(n1501), .Y(
        n2611) );
  OAI221XL U1199 ( .A0(n27), .A1(n874), .B0(n229), .B1(n899), .C0(n1509), .Y(
        n2619) );
  AOI21X1 U1200 ( .A0(N1058), .A1(n243), .B0(n274), .Y(n1509) );
  OAI221XL U1201 ( .A0(n26), .A1(n873), .B0(n230), .B1(n898), .C0(n1510), .Y(
        n2620) );
  AOI21X1 U1202 ( .A0(N1057), .A1(n243), .B0(n274), .Y(n1510) );
  OAI221XL U1203 ( .A0(n35), .A1(n863), .B0(n231), .B1(n883), .C0(n1617), .Y(
        n2801) );
  AOI21X1 U1204 ( .A0(N1035), .A1(n242), .B0(n274), .Y(n1617) );
  OAI221XL U1205 ( .A0(n22), .A1(n855), .B0(n231), .B1(n875), .C0(n1625), .Y(
        n2809) );
  AOI21X1 U1206 ( .A0(N1027), .A1(n240), .B0(n275), .Y(n1625) );
  OAI221XL U1207 ( .A0(n22), .A1(n853), .B0(n230), .B1(n873), .C0(n1627), .Y(
        n2811) );
  AOI21X1 U1208 ( .A0(N1025), .A1(n240), .B0(n275), .Y(n1627) );
  OAI221XL U1209 ( .A0(n25), .A1(n813), .B0(n232), .B1(n846), .C0(n1696), .Y(
        n2863) );
  AOI21X1 U1210 ( .A0(N973), .A1(n241), .B0(n275), .Y(n1696) );
  OAI221XL U1211 ( .A0(n25), .A1(n690), .B0(n218), .B1(n776), .C0(n1770), .Y(
        n2938) );
  OAI221XL U1212 ( .A0(n21), .A1(n685), .B0(n218), .B1(n771), .C0(n1775), .Y(
        n2943) );
  AOI21X1 U1213 ( .A0(N894), .A1(n242), .B0(n272), .Y(n1775) );
  OAI221XL U1214 ( .A0(n33), .A1(n684), .B0(n219), .B1(n770), .C0(n1776), .Y(
        n2944) );
  OAI221XL U1215 ( .A0(n17), .A1(n681), .B0(n219), .B1(n767), .C0(n1779), .Y(
        n2947) );
  OAI221XL U1216 ( .A0(n30), .A1(n787), .B0(n228), .B1(n814), .C0(n1727), .Y(
        n2894) );
  AOI21X1 U1217 ( .A0(N942), .A1(n235), .B0(n276), .Y(n1727) );
  OAI221XL U1218 ( .A0(n30), .A1(n769), .B0(n221), .B1(n796), .C0(n1745), .Y(
        n2912) );
  OAI221XL U1219 ( .A0(n18), .A1(n781), .B0(n219), .B1(n808), .C0(n1733), .Y(
        n2900) );
  AOI21X1 U1220 ( .A0(N936), .A1(n240), .B0(n277), .Y(n1733) );
  OAI221XL U1221 ( .A0(n31), .A1(n766), .B0(n222), .B1(n793), .C0(n1748), .Y(
        n2915) );
  OAI221XL U1222 ( .A0(n27), .A1(n802), .B0(n225), .B1(n835), .C0(n1707), .Y(
        n2874) );
  AOI21X1 U1223 ( .A0(N962), .A1(n239), .B0(n276), .Y(n1707) );
  OAI221XL U1224 ( .A0(n31), .A1(n885), .B0(n233), .B1(n910), .C0(n1498), .Y(
        n2608) );
  AOI21X1 U1225 ( .A0(N1069), .A1(n242), .B0(n274), .Y(n1498) );
  OAI221XL U1226 ( .A0(n18), .A1(n876), .B0(n218), .B1(n901), .C0(n1507), .Y(
        n2617) );
  AOI21X1 U1227 ( .A0(N1060), .A1(n243), .B0(n274), .Y(n1507) );
  OAI221XL U1228 ( .A0(n28), .A1(n875), .B0(n229), .B1(n900), .C0(n1508), .Y(
        n2618) );
  AOI21X1 U1229 ( .A0(N1059), .A1(n243), .B0(n274), .Y(n1508) );
  OAI221XL U1230 ( .A0(n25), .A1(n871), .B0(n230), .B1(n896), .C0(n1512), .Y(
        n2622) );
  OAI221XL U1231 ( .A0(n20), .A1(n866), .B0(n231), .B1(n891), .C0(n1517), .Y(
        n2627) );
  OAI221XL U1232 ( .A0(n31), .A1(n857), .B0(n221), .B1(n877), .C0(n1623), .Y(
        n2807) );
  AOI21X1 U1233 ( .A0(N1029), .A1(n241), .B0(n274), .Y(n1623) );
  OAI221XL U1234 ( .A0(n14), .A1(n811), .B0(n232), .B1(n844), .C0(n1698), .Y(
        n2865) );
  OAI221XL U1235 ( .A0(n23), .A1(n852), .B0(n232), .B1(n872), .C0(n1628), .Y(
        n2812) );
  OAI221XL U1236 ( .A0(n19), .A1(n804), .B0(n225), .B1(n837), .C0(n1705), .Y(
        n2872) );
  AOI21X1 U1237 ( .A0(N964), .A1(n240), .B0(n275), .Y(n1705) );
  OAI221XL U1238 ( .A0(n28), .A1(n803), .B0(n225), .B1(n836), .C0(n1706), .Y(
        n2873) );
  AOI21X1 U1239 ( .A0(N963), .A1(n237), .B0(n275), .Y(n1706) );
  OAI221XL U1240 ( .A0(n29), .A1(n797), .B0(n227), .B1(n830), .C0(n1712), .Y(
        n2879) );
  AOI21X1 U1241 ( .A0(N957), .A1(n239), .B0(n276), .Y(n1712) );
  OAI221XL U1242 ( .A0(n36), .A1(n795), .B0(n227), .B1(n828), .C0(n1714), .Y(
        n2881) );
  AOI21X1 U1243 ( .A0(N955), .A1(n235), .B0(n276), .Y(n1714) );
  OAI221XL U1244 ( .A0(n16), .A1(n809), .B0(n232), .B1(n842), .C0(n1700), .Y(
        n2867) );
  AOI21X1 U1245 ( .A0(N969), .A1(n242), .B0(n275), .Y(n1700) );
  OAI221XL U1246 ( .A0(n35), .A1(n801), .B0(n226), .B1(n834), .C0(n1708), .Y(
        n2875) );
  AOI21X1 U1247 ( .A0(N961), .A1(n240), .B0(n276), .Y(n1708) );
  OAI221XL U1248 ( .A0(n36), .A1(n799), .B0(n227), .B1(n832), .C0(n1710), .Y(
        n2877) );
  AOI21X1 U1249 ( .A0(N959), .A1(n239), .B0(n276), .Y(n1710) );
  OAI221XL U1250 ( .A0(n28), .A1(n792), .B0(n229), .B1(n825), .C0(n1717), .Y(
        n2884) );
  AOI21X1 U1251 ( .A0(N952), .A1(n237), .B0(n276), .Y(n1717) );
  OAI221XL U1252 ( .A0(n27), .A1(n791), .B0(n228), .B1(n824), .C0(n1718), .Y(
        n2885) );
  AOI21X1 U1253 ( .A0(N951), .A1(n239), .B0(n276), .Y(n1718) );
  OAI221XL U1254 ( .A0(n24), .A1(n806), .B0(n224), .B1(n839), .C0(n1703), .Y(
        n2870) );
  AOI21X1 U1255 ( .A0(N966), .A1(n240), .B0(n275), .Y(n1703) );
  OAI221XL U1256 ( .A0(n15), .A1(n805), .B0(n224), .B1(n838), .C0(n1704), .Y(
        n2871) );
  AOI21X1 U1257 ( .A0(N965), .A1(n242), .B0(n275), .Y(n1704) );
  OAI221XL U1258 ( .A0(n14), .A1(n800), .B0(n226), .B1(n833), .C0(n1709), .Y(
        n2876) );
  AOI21X1 U1259 ( .A0(N960), .A1(n237), .B0(n276), .Y(n1709) );
  NAND3BX1 U1260 ( .AN(n1849), .B(n1337), .C(n342), .Y(n343) );
  INVX1 U1261 ( .A(n1859), .Y(n342) );
  OAI211X1 U1262 ( .A0(n18), .A1(n630), .B0(n629), .C0(n628), .Y(n3005) );
  OAI211X1 U1263 ( .A0(n15), .A1(n472), .B0(n471), .C0(n470), .Y(n2848) );
  OAI211X1 U1264 ( .A0(n20), .A1(n477), .B0(n476), .C0(n475), .Y(n2849) );
  NAND2X1 U1265 ( .A(n153), .B(n195), .Y(n476) );
  OAI211X1 U1266 ( .A0(n12), .A1(n486), .B0(n485), .C0(n484), .Y(n2851) );
  OAI211X1 U1267 ( .A0(n19), .A1(n633), .B0(n632), .C0(n631), .Y(n3006) );
  INVX1 U1268 ( .A(next_A[12]), .Y(n633) );
  OAI211X1 U1269 ( .A0(n16), .A1(n641), .B0(n640), .C0(n639), .Y(n3009) );
  INVX1 U1270 ( .A(next_A[9]), .Y(n641) );
  OAI211X1 U1271 ( .A0(n28), .A1(n650), .B0(n649), .C0(n648), .Y(n3012) );
  NAND2X1 U1272 ( .A(N857), .B(n248), .Y(n649) );
  OAI211X1 U1273 ( .A0(n21), .A1(n654), .B0(n653), .C0(n652), .Y(n3013) );
  OAI211X1 U1274 ( .A0(n33), .A1(n659), .B0(n658), .C0(n657), .Y(n3014) );
  NAND2X1 U1275 ( .A(n179), .B(n197), .Y(n658) );
  OAI211X1 U1276 ( .A0(n24), .A1(n665), .B0(n664), .C0(n663), .Y(n3015) );
  NAND2X1 U1277 ( .A(n180), .B(n194), .Y(n664) );
  NAND2X1 U1278 ( .A(N854), .B(n245), .Y(n663) );
  OAI211X1 U1279 ( .A0(n26), .A1(n669), .B0(n668), .C0(n667), .Y(n3016) );
  INVX1 U1280 ( .A(next_A[2]), .Y(n669) );
  OAI211X1 U1281 ( .A0(n34), .A1(n673), .B0(n672), .C0(n671), .Y(n3017) );
  NAND2BX1 U1282 ( .AN(n540), .B(n539), .Y(n2952) );
  OAI21XL U1283 ( .A0(n762), .A1(n215), .B0(n636), .Y(n540) );
  XOR3X2 U1284 ( .A(n163), .B(n174), .C(n156), .Y(f3_A_32[7]) );
  XOR3X2 U1285 ( .A(n165), .B(n176), .C(n157), .Y(f3_A_32[5]) );
  XOR3X2 U1286 ( .A(n162), .B(n173), .C(n155), .Y(f3_A_32[8]) );
  XOR3X2 U1287 ( .A(n72), .B(n170), .C(n160), .Y(f3_A_32[11]) );
  XOR3X2 U1288 ( .A(n166), .B(n177), .C(n158), .Y(f3_A_32[4]) );
  XOR3X2 U1289 ( .A(n70), .B(n171), .C(n161), .Y(f3_A_32[10]) );
  XOR3X2 U1290 ( .A(n180), .B(n168), .C(n158), .Y(f3_A_32[13]) );
  OAI21XL U1291 ( .A0(n191), .A1(n786), .B0(n1760), .Y(n2928) );
  AOI22X1 U1292 ( .A0(N909), .A1(n237), .B0(n158), .B1(n11), .Y(n1760) );
  OAI21XL U1293 ( .A0(n190), .A1(n779), .B0(n1767), .Y(n2935) );
  OAI21XL U1294 ( .A0(n190), .A1(n768), .B0(n1778), .Y(n2946) );
  AOI22X1 U1295 ( .A0(N891), .A1(n237), .B0(n175), .B1(n11), .Y(n1778) );
  OAI21XL U1296 ( .A0(n190), .A1(n774), .B0(n1772), .Y(n2940) );
  AOI22X1 U1297 ( .A0(N897), .A1(n241), .B0(n169), .B1(n10), .Y(n1772) );
  OAI21XL U1298 ( .A0(n190), .A1(n772), .B0(n1774), .Y(n2942) );
  AOI22X1 U1299 ( .A0(N895), .A1(n237), .B0(n171), .B1(n11), .Y(n1774) );
  OAI21XL U1300 ( .A0(n190), .A1(n766), .B0(n1780), .Y(n2948) );
  AOI22X1 U1301 ( .A0(N889), .A1(n237), .B0(n177), .B1(n11), .Y(n1780) );
  OAI21XL U1302 ( .A0(n190), .A1(n765), .B0(n1781), .Y(n2949) );
  OAI21XL U1303 ( .A0(n190), .A1(n764), .B0(n1782), .Y(n2950) );
  OAI21XL U1304 ( .A0(n187), .A1(n876), .B0(n1624), .Y(n2808) );
  AOI22X1 U1305 ( .A0(N1028), .A1(n236), .B0(n148), .B1(n10), .Y(n1624) );
  OAI21XL U1306 ( .A0(n187), .A1(n867), .B0(n1633), .Y(n2817) );
  OAI21XL U1307 ( .A0(n187), .A1(n874), .B0(n1626), .Y(n2810) );
  OAI21XL U1308 ( .A0(n187), .A1(n871), .B0(n1629), .Y(n2813) );
  OAI21XL U1309 ( .A0(n191), .A1(n783), .B0(n1763), .Y(n2931) );
  OAI21XL U1310 ( .A0(n191), .A1(n780), .B0(n1766), .Y(n2934) );
  AOI22X1 U1311 ( .A0(N903), .A1(n237), .B0(n163), .B1(n10), .Y(n1766) );
  OAI21XL U1312 ( .A0(n190), .A1(n763), .B0(n1783), .Y(n2951) );
  OAI21XL U1313 ( .A0(n187), .A1(n878), .B0(n1622), .Y(n2806) );
  AOI22X1 U1314 ( .A0(N1030), .A1(n235), .B0(n147), .B1(n10), .Y(n1622) );
  OAI21XL U1315 ( .A0(n187), .A1(n869), .B0(n1631), .Y(n2815) );
  OAI21XL U1316 ( .A0(n187), .A1(n868), .B0(n1632), .Y(n2816) );
  OAI21XL U1317 ( .A0(n188), .A1(n880), .B0(n1620), .Y(n2804) );
  AOI22X1 U1318 ( .A0(N1032), .A1(n235), .B0(n146), .B1(n10), .Y(n1620) );
  OAI21XL U1319 ( .A0(n187), .A1(n879), .B0(n1621), .Y(n2805) );
  AOI22X1 U1320 ( .A0(N1031), .A1(n235), .B0(SHA256_result[116]), .B1(n11), 
        .Y(n1621) );
  OAI21XL U1321 ( .A0(n189), .A1(n865), .B0(n1635), .Y(n2819) );
  NAND3BX1 U1322 ( .AN(n533), .B(n532), .C(n531), .Y(n2929) );
  OAI21XL U1323 ( .A0(n785), .A1(n216), .B0(n636), .Y(n533) );
  NAND2BX1 U1324 ( .AN(n30), .B(n159), .Y(n532) );
  NAND2X1 U1325 ( .A(N908), .B(n247), .Y(n531) );
  NAND3BX1 U1326 ( .AN(n536), .B(n535), .C(n534), .Y(n2930) );
  OAI21XL U1327 ( .A0(n784), .A1(n215), .B0(n636), .Y(n536) );
  NAND2X1 U1328 ( .A(N907), .B(n247), .Y(n534) );
  NAND2BX1 U1329 ( .AN(n18), .B(n160), .Y(n535) );
  NAND3BX1 U1330 ( .AN(n346), .B(n345), .C(n344), .Y(n2598) );
  NAND2BX1 U1331 ( .AN(n921), .B(n350), .Y(n344) );
  NAND2BX1 U1334 ( .AN(n675), .B(N1079), .Y(n345) );
  OAI21XL U1337 ( .A0(n15), .A1(n400), .B0(n636), .Y(n346) );
  NAND3BX1 U1340 ( .AN(n349), .B(n348), .C(n347), .Y(n2599) );
  NAND2BX1 U1343 ( .AN(n920), .B(n350), .Y(n347) );
  NAND2BX1 U1344 ( .AN(n675), .B(N1078), .Y(n348) );
  OAI21XL U1347 ( .A0(n17), .A1(n402), .B0(n636), .Y(n349) );
  NAND3BX1 U1350 ( .AN(n353), .B(n352), .C(n351), .Y(n2602) );
  NAND2BX1 U1355 ( .AN(n917), .B(n350), .Y(n351) );
  NAND2BX1 U1360 ( .AN(n675), .B(N1075), .Y(n352) );
  OAI21XL U1361 ( .A0(n13), .A1(n94), .B0(n636), .Y(n353) );
  OAI211X1 U1364 ( .A0(n12), .A1(n468), .B0(n467), .C0(n466), .Y(n2847) );
  NAND2X1 U1367 ( .A(n151), .B(n195), .Y(n467) );
  NAND2X1 U1370 ( .A(n459), .B(n458), .Y(n2845) );
  NAND2BX1 U1373 ( .AN(n515), .B(n514), .Y(n2886) );
  OAI21XL U1374 ( .A0(n823), .A1(n215), .B0(n636), .Y(n515) );
  NAND2BX1 U1377 ( .AN(n517), .B(n516), .Y(n2888) );
  OAI21XL U1380 ( .A0(n821), .A1(n234), .B0(n636), .Y(n517) );
  NAND2BX1 U1385 ( .AN(n538), .B(n537), .Y(n2932) );
  OAI21XL U1391 ( .A0(n782), .A1(n215), .B0(n636), .Y(n538) );
  OAI2BB1X1 U1392 ( .A0N(N862), .A1N(n245), .B0(n635), .Y(n3007) );
  AOI2BB2X1 U1393 ( .B0(n192), .B1(n172), .A0N(n21), .A1N(n634), .Y(n635) );
  INVXL U1394 ( .A(next_A[11]), .Y(n634) );
  NAND2X1 U1397 ( .A(n677), .B(n676), .Y(n3018) );
  NAND2X1 U1400 ( .A(n638), .B(n637), .Y(n3008) );
  AOI21X1 U1403 ( .A0(n214), .A1(n173), .B0(n276), .Y(n637) );
  AOI22XL U1406 ( .A0(next_A[10]), .A1(n11), .B0(N861), .B1(n239), .Y(n638) );
  INVX1 U1407 ( .A(n662), .Y(n185) );
  OAI21XL U1410 ( .A0(first_block_core), .A1(n343), .B0(n1491), .Y(n662) );
  XOR3X2 U1413 ( .A(n179), .B(n167), .C(n157), .Y(f3_A_32[14]) );
  XOR3X2 U1419 ( .A(n164), .B(n176), .C(n155), .Y(f3_A_32[17]) );
  XOR3X2 U1425 ( .A(n70), .B(n174), .C(n162), .Y(f3_A_32[19]) );
  XOR3X2 U1426 ( .A(n181), .B(n169), .C(n159), .Y(f3_A_32[12]) );
  INVX1 U1429 ( .A(n1489), .Y(n705) );
  OAI21XL U1432 ( .A0(first_block_core), .A1(n1490), .B0(n1491), .Y(n1489) );
  NOR2X1 U1433 ( .A(n1975), .B(n1977), .Y(n1976) );
  NOR2X1 U1436 ( .A(round[2]), .B(round[3]), .Y(n2501) );
  AOI31X1 U1439 ( .A0(n2466), .A1(n2467), .A2(n2468), .B0(n268), .Y(N3012) );
  AOI2BB2X1 U1440 ( .B0(n2400), .B1(n332), .A0N(n758), .A1N(n2472), .Y(n2466)
         );
  AOI211X1 U1441 ( .A0(n2332), .A1(n1397), .B0(n2469), .C0(n2470), .Y(n2468)
         );
  AOI31X1 U1444 ( .A0(n2450), .A1(n2451), .A2(n2452), .B0(n268), .Y(N3014) );
  NOR3BX1 U1447 ( .AN(n2456), .B(n2348), .C(n2354), .Y(n2451) );
  AOI211X1 U1448 ( .A0(n2457), .A1(n2435), .B0(n2458), .C0(n2275), .Y(n2450)
         );
  AOI211X1 U1453 ( .A0(n2332), .A1(n336), .B0(n2453), .C0(n2454), .Y(n2452) );
  AOI31X1 U1454 ( .A0(n2393), .A1(n2394), .A2(n2395), .B0(n269), .Y(N3020) );
  AOI211X1 U1459 ( .A0(n2332), .A1(n336), .B0(n2396), .C0(n2281), .Y(n2395) );
  AOI211X1 U1461 ( .A0(n40), .A1(n2398), .B0(n2247), .C0(n2321), .Y(n2394) );
  AOI31X1 U1462 ( .A0(n2510), .A1(n2511), .A2(n2512), .B0(n268), .Y(N3006) );
  AOI221X1 U1463 ( .A0(n2406), .A1(n182), .B0(n2357), .B1(n1397), .C0(n2503), 
        .Y(n2510) );
  NOR4BX1 U1464 ( .AN(n2513), .B(n2285), .C(n2370), .D(n2437), .Y(n2512) );
  AOI31X1 U1465 ( .A0(n2362), .A1(n709), .A2(n2363), .B0(n269), .Y(N3023) );
  AOI222X1 U1466 ( .A0(n2372), .A1(n1397), .B0(n47), .B1(n2374), .C0(n2262), 
        .C1(n2375), .Y(n2362) );
  INVX1 U1467 ( .A(n2368), .Y(n709) );
  AOI211X1 U1468 ( .A0(n2244), .A1(n131), .B0(n2365), .C0(n2366), .Y(n2363) );
  AOI31X1 U1469 ( .A0(n2439), .A1(n2440), .A2(n2441), .B0(n268), .Y(N3015) );
  AOI222X1 U1470 ( .A0(n2448), .A1(n1397), .B0(n2299), .B1(n329), .C0(n2428), 
        .C1(n2449), .Y(n2439) );
  AOI211X1 U1471 ( .A0(n183), .A1(n2442), .B0(n2443), .C0(n2444), .Y(n2441) );
  AOI31X1 U1472 ( .A0(n2528), .A1(n2529), .A2(n2530), .B0(n268), .Y(N3003) );
  NOR3X1 U1473 ( .A(n2259), .B(n2300), .C(n743), .Y(n2529) );
  AOI211X1 U1474 ( .A0(n2344), .A1(n47), .B0(n2531), .C0(n2454), .Y(n2530) );
  AOI31X1 U1475 ( .A0(n2248), .A1(n2249), .A2(n2250), .B0(n269), .Y(N3032) );
  AOI22X1 U1476 ( .A0(n2261), .A1(n2262), .B0(n2263), .B1(n332), .Y(n2248) );
  AOI222X1 U1477 ( .A0(n2257), .A1(n182), .B0(n2258), .B1(n2259), .C0(n2260), 
        .C1(n335), .Y(n2249) );
  AOI211X1 U1478 ( .A0(n2251), .A1(n129), .B0(n2253), .C0(n2254), .Y(n2250) );
  AOI31X1 U1479 ( .A0(n2383), .A1(n2384), .A2(n2385), .B0(n269), .Y(N3021) );
  AOI222X1 U1480 ( .A0(n131), .A1(n2374), .B0(n2390), .B1(n336), .C0(n2391), 
        .C1(n2349), .Y(n2384) );
  NOR4BX1 U1481 ( .AN(n2386), .B(n2297), .C(n2387), .D(n2263), .Y(n2385) );
  AOI31X1 U1482 ( .A0(n2504), .A1(n2505), .A2(n2506), .B0(n268), .Y(N3007) );
  NOR4BX1 U1483 ( .AN(n739), .B(n2332), .C(n2507), .D(n2300), .Y(n2506) );
  AOI221X1 U1484 ( .A0(n2448), .A1(n336), .B0(n2417), .B1(n335), .C0(n2509), 
        .Y(n2504) );
  AOI31X1 U1485 ( .A0(n2326), .A1(n2327), .A2(n2328), .B0(n269), .Y(N3026) );
  AOI2BB2X1 U1486 ( .B0(n335), .B1(n2332), .A0N(n2333), .A1N(n333), .Y(n2326)
         );
  AOI211X1 U1487 ( .A0(n2329), .A1(n1397), .B0(n2330), .C0(n2331), .Y(n2328)
         );
  AOI31X1 U1488 ( .A0(n2474), .A1(n2475), .A2(n2476), .B0(n268), .Y(N3011) );
  NOR4BX1 U1489 ( .AN(n2289), .B(n2437), .C(n2477), .D(n2478), .Y(n2476) );
  AOI22X1 U1490 ( .A0(n2297), .A1(n329), .B0(n47), .B1(n2479), .Y(n2475) );
  NOR2X1 U1491 ( .A(n2420), .B(n2470), .Y(n2474) );
  AOI31X1 U1492 ( .A0(n2334), .A1(n2335), .A2(n2336), .B0(n269), .Y(N3025) );
  NOR3X1 U1493 ( .A(n2347), .B(n2285), .C(n2348), .Y(n2335) );
  AOI31X1 U1494 ( .A0(n2430), .A1(n2431), .A2(n2432), .B0(n268), .Y(N3016) );
  NOR4BX1 U1495 ( .AN(n2433), .B(n2434), .C(n2435), .D(n2348), .Y(n2432) );
  AOI31X1 U1496 ( .A0(n2411), .A1(n2412), .A2(n2413), .B0(n269), .Y(N3018) );
  NOR4BX1 U1497 ( .AN(n2288), .B(n2414), .C(n2415), .D(n2416), .Y(n2413) );
  AOI211X1 U1498 ( .A0(n2284), .A1(n2261), .B0(n2418), .C0(n2419), .Y(n2412)
         );
  AOI21X1 U1499 ( .A0(n2321), .A1(n328), .B0(n2420), .Y(n2411) );
  AOI31X1 U1500 ( .A0(n2276), .A1(n2277), .A2(n2278), .B0(n269), .Y(N3030) );
  NOR3BX1 U1501 ( .AN(n2283), .B(n2284), .C(n2285), .Y(n2277) );
  NOR3BX1 U1502 ( .AN(n2279), .B(n2280), .C(n2281), .Y(n2278) );
  AOI31X1 U1503 ( .A0(n2533), .A1(n2534), .A2(n2535), .B0(n268), .Y(N3002) );
  AOI222X1 U1504 ( .A0(n47), .A1(n2343), .B0(n2473), .B1(n2262), .C0(n2298), 
        .C1(round[3]), .Y(n2533) );
  AND4X2 U1505 ( .A(n2536), .B(n729), .C(n2288), .D(n2255), .Y(n2535) );
  AOI21X1 U1506 ( .A0(n2167), .A1(n2168), .B0(n1975), .Y(N3444) );
  NOR4X1 U1507 ( .A(n2169), .B(n2170), .C(n2171), .D(n2172), .Y(n2168) );
  NOR4X1 U1508 ( .A(n2207), .B(n2208), .C(n2209), .D(n2210), .Y(n2167) );
  NAND4X1 U1509 ( .A(n2201), .B(n2202), .C(n2203), .D(n2204), .Y(n2169) );
  AOI21X1 U1510 ( .A0(n2125), .A1(n2126), .B0(n1975), .Y(N3445) );
  NOR4X1 U1511 ( .A(n2127), .B(n2128), .C(n2129), .D(n2130), .Y(n2126) );
  NOR4X1 U1512 ( .A(n2147), .B(n2148), .C(n2149), .D(n2150), .Y(n2125) );
  NAND4X1 U1513 ( .A(n2143), .B(n2144), .C(n2145), .D(n2146), .Y(n2127) );
  AOI21X1 U1514 ( .A0(n2083), .A1(n2084), .B0(n1975), .Y(N3446) );
  NOR4X1 U1515 ( .A(n2085), .B(n2086), .C(n2087), .D(n2088), .Y(n2084) );
  NOR4X1 U1516 ( .A(n2105), .B(n2106), .C(n2107), .D(n2108), .Y(n2083) );
  NAND4X1 U1517 ( .A(n2101), .B(n2102), .C(n2103), .D(n2104), .Y(n2085) );
  AOI21X1 U1518 ( .A0(n1978), .A1(n1979), .B0(n1975), .Y(N3447) );
  NOR4X1 U1519 ( .A(n1980), .B(n1981), .C(n1982), .D(n1983), .Y(n1979) );
  NOR4X1 U1520 ( .A(n2031), .B(n2032), .C(n2033), .D(n2034), .Y(n1978) );
  NAND4X1 U1521 ( .A(n2020), .B(n2021), .C(n2022), .D(n2023), .Y(n1980) );
  XOR3X2 U1522 ( .A(n165), .B(n177), .C(n156), .Y(f3_A_32[16]) );
  XOR3X2 U1524 ( .A(n179), .B(n170), .C(n159), .Y(f3_A_32[23]) );
  XOR3X2 U1525 ( .A(n181), .B(n172), .C(n161), .Y(f3_A_32[21]) );
  XOR3X2 U1526 ( .A(n180), .B(n171), .C(n160), .Y(f3_A_32[22]) );
  AOI21X1 U1527 ( .A0(n2497), .A1(n2498), .B0(n268), .Y(N3008) );
  AOI211X1 U1528 ( .A0(n2446), .A1(round[3]), .B0(n2502), .C0(n2503), .Y(n2497) );
  AOI211X1 U1529 ( .A0(n2486), .A1(n335), .B0(n2499), .C0(n2500), .Y(n2498) );
  OAI222XL U1530 ( .A0(n1397), .A1(n741), .B0(n182), .B1(n2272), .C0(n2261), 
        .C1(n752), .Y(n2502) );
  INVX1 U1531 ( .A(n144), .Y(n269) );
  XOR3X2 U1532 ( .A(n178), .B(n169), .C(n158), .Y(f3_A_32[24]) );
  XOR3X2 U1533 ( .A(n166), .B(n175), .C(n156), .Y(f3_A_32[27]) );
  XOR3X2 U1534 ( .A(n168), .B(n177), .C(n157), .Y(f3_A_32[25]) );
  XOR3X2 U1535 ( .A(n165), .B(n174), .C(n155), .Y(f3_A_32[28]) );
  INVX1 U1536 ( .A(n334), .Y(n333) );
  INVX1 U1537 ( .A(n2263), .Y(n714) );
  OAI211X1 U1538 ( .A0(round[2]), .A1(n714), .B0(n2333), .C0(n2356), .Y(n2454)
         );
  NOR2X1 U1539 ( .A(n754), .B(n328), .Y(n2465) );
  INVX1 U1540 ( .A(n2438), .Y(n723) );
  NAND3X1 U1541 ( .A(n710), .B(n2256), .C(n2279), .Y(n2420) );
  NOR2X1 U1542 ( .A(n328), .B(n746), .Y(n2445) );
  XOR3X2 U1543 ( .A(n70), .B(n172), .C(n163), .Y(f3_A_32[30]) );
  OAI2BB1X1 U1544 ( .A0N(n183), .A1N(n2425), .B0(n720), .Y(n2405) );
  INVX1 U1545 ( .A(n2262), .Y(n757) );
  INVX1 U1546 ( .A(n2349), .Y(n755) );
  OAI2BB1X1 U1547 ( .A0N(n335), .A1N(n2427), .B0(n2526), .Y(n2525) );
  AOI31X1 U1548 ( .A0(n737), .A1(n751), .A2(n2397), .B0(round[0]), .Y(n2527)
         );
  NOR3X1 U1549 ( .A(n332), .B(round[0]), .C(n755), .Y(n2437) );
  NOR2X1 U1550 ( .A(n182), .B(n183), .Y(n2428) );
  OAI222XL U1551 ( .A0(n730), .A1(n744), .B0(n2436), .B1(n717), .C0(n40), .C1(
        n711), .Y(n2434) );
  NOR2X1 U1552 ( .A(n2259), .B(n2428), .Y(n2436) );
  OAI222XL U1553 ( .A0(n182), .A1(n716), .B0(n742), .B1(n721), .C0(n335), .C1(
        n2282), .Y(n2280) );
  NOR3X1 U1554 ( .A(n335), .B(round[2]), .C(n752), .Y(n2435) );
  OAI222XL U1555 ( .A0(round[0]), .A1(n2495), .B0(n726), .B1(n741), .C0(n335), 
        .C1(n733), .Y(n2491) );
  NOR2X1 U1556 ( .A(n2289), .B(round[2]), .Y(n2348) );
  OAI222XL U1557 ( .A0(n140), .A1(n2296), .B0(n2519), .B1(n745), .C0(n2532), 
        .C1(n726), .Y(n2531) );
  INVX1 U1558 ( .A(n2390), .Y(n745) );
  NOR3X1 U1559 ( .A(n2355), .B(n40), .C(n2447), .Y(n2532) );
  NOR2X1 U1560 ( .A(n2298), .B(n2300), .Y(n2367) );
  OAI31X1 U1561 ( .A0(n725), .A1(n183), .A2(round[3]), .B0(n2388), .Y(n2387)
         );
  AOI31X1 U1562 ( .A0(n726), .A1(n757), .A2(n47), .B0(n2389), .Y(n2388) );
  NOR2X1 U1563 ( .A(n742), .B(round[3]), .Y(n2299) );
  NOR3X1 U1564 ( .A(round[0]), .B(n182), .C(n754), .Y(n2416) );
  NAND2X1 U1565 ( .A(n2521), .B(round[0]), .Y(n2282) );
  NOR2X1 U1566 ( .A(n717), .B(round[2]), .Y(n2344) );
  NOR2X1 U1567 ( .A(n726), .B(round[2]), .Y(n2343) );
  NOR2X1 U1568 ( .A(n738), .B(round[2]), .Y(n2260) );
  OAI221XL U1569 ( .A0(n738), .A1(n2272), .B0(n726), .B1(n739), .C0(n2455), 
        .Y(n2453) );
  OAI21XL U1570 ( .A0(n2306), .A1(n2314), .B0(n333), .Y(n2455) );
  NOR2X1 U1571 ( .A(n738), .B(round[3]), .Y(n2312) );
  OAI211X1 U1572 ( .A0(n182), .A1(n725), .B0(n707), .C0(n719), .Y(n2324) );
  OAI22X1 U1573 ( .A0(n328), .A1(n750), .B0(n736), .B1(n140), .Y(n2470) );
  NOR3X1 U1574 ( .A(n328), .B(n182), .C(n757), .Y(n2496) );
  AOI221X1 U1575 ( .A0(n708), .A1(n182), .B0(n183), .B1(n335), .C0(n2473), .Y(
        n2472) );
  NAND2X1 U1576 ( .A(n129), .B(n2262), .Y(n2272) );
  INVX1 U1577 ( .A(n40), .Y(n742) );
  NOR2X1 U1578 ( .A(n749), .B(round[3]), .Y(n2521) );
  AOI211X1 U1579 ( .A0(n183), .A1(n2380), .B0(n2300), .C0(n2267), .Y(n2379) );
  OAI21XL U1580 ( .A0(n335), .A1(n755), .B0(n721), .Y(n2380) );
  NOR2X1 U1581 ( .A(n2397), .B(n730), .Y(n2354) );
  AOI31X1 U1582 ( .A0(n735), .A1(n741), .A2(n2296), .B0(n730), .Y(n2295) );
  INVX1 U1583 ( .A(n2259), .Y(n741) );
  NOR2X1 U1584 ( .A(n738), .B(n328), .Y(n2375) );
  NOR2X1 U1585 ( .A(n717), .B(n182), .Y(n2381) );
  OAI211X1 U1586 ( .A0(n182), .A1(round[2]), .B0(n737), .C0(n747), .Y(n2408)
         );
  INVX1 U1587 ( .A(n2251), .Y(n747) );
  NOR2X1 U1588 ( .A(n328), .B(n752), .Y(n2371) );
  NAND2X1 U1589 ( .A(n2371), .B(round[3]), .Y(n2288) );
  OAI211X1 U1590 ( .A0(n730), .A1(n736), .B0(n727), .C0(n2256), .Y(n2253) );
  NOR2X1 U1591 ( .A(n755), .B(n183), .Y(n2318) );
  OAI211X1 U1592 ( .A0(n2464), .A1(n1397), .B0(n2283), .C0(n731), .Y(n2462) );
  AOI21X1 U1593 ( .A0(n40), .A1(n754), .B0(n2390), .Y(n2464) );
  OAI2BB2X1 U1594 ( .B0(n335), .B1(n2397), .A0N(n328), .A1N(n2267), .Y(n2281)
         );
  NOR2X1 U1595 ( .A(n757), .B(round[0]), .Y(n2409) );
  NOR2X1 U1596 ( .A(n757), .B(n183), .Y(n2355) );
  OAI21XL U1597 ( .A0(round[0]), .A1(n758), .B0(n725), .Y(n2449) );
  NAND4X1 U1598 ( .A(n2151), .B(n2152), .C(n2153), .D(n2154), .Y(n2150) );
  AOI22X1 U1599 ( .A0(n2045), .A1(n159), .B0(n2046), .B1(n156), .Y(n2151) );
  AOI22X1 U1600 ( .A0(n2041), .A1(n174), .B0(n2042), .B1(n170), .Y(n2153) );
  AOI22X1 U1601 ( .A0(n2043), .A1(n166), .B0(n2044), .B1(n162), .Y(n2152) );
  OAI21XL U1602 ( .A0(n182), .A1(n756), .B0(n2289), .Y(n2239) );
  INVX1 U1603 ( .A(n2446), .Y(n706) );
  NAND2BX1 U1604 ( .AN(n2296), .B(n129), .Y(n2386) );
  NOR3X1 U1605 ( .A(n754), .B(round[0]), .C(n742), .Y(n2309) );
  INVX1 U1606 ( .A(n2357), .Y(n740) );
  NAND2X1 U1607 ( .A(n2267), .B(round[0]), .Y(n2456) );
  NAND2X1 U1608 ( .A(n2349), .B(n131), .Y(n2255) );
  NAND2X1 U1609 ( .A(n2244), .B(n40), .Y(n2495) );
  NOR2X1 U1610 ( .A(n750), .B(round[3]), .Y(n2273) );
  NOR2X1 U1611 ( .A(n2282), .B(round[2]), .Y(n2417) );
  AOI22X1 U1612 ( .A0(n2039), .A1(n72), .B0(n2040), .B1(n178), .Y(n2154) );
  AOI22X1 U1613 ( .A0(n2039), .A1(n181), .B0(n2040), .B1(n177), .Y(n2112) );
  AOI22X1 U1614 ( .A0(n2039), .A1(n180), .B0(n2040), .B1(n176), .Y(n2038) );
  AOI21X1 U1615 ( .A0(n2256), .A1(n747), .B0(n1397), .Y(n2484) );
  NAND3BX1 U1616 ( .AN(n2273), .B(n746), .C(n2392), .Y(n2338) );
  NAND3X1 U1617 ( .A(round[3]), .B(n328), .C(n40), .Y(n2392) );
  CLKINVX3 U1618 ( .A(n336), .Y(n335) );
  NAND3X1 U1619 ( .A(n713), .B(n2323), .C(n2508), .Y(n2507) );
  OAI21XL U1620 ( .A0(n2438), .A1(n2406), .B0(n182), .Y(n2508) );
  INVX1 U1621 ( .A(n2410), .Y(n736) );
  OAI221XL U1622 ( .A0(n335), .A1(n2269), .B0(round[2]), .B1(n718), .C0(n2270), 
        .Y(n2268) );
  OAI21XL U1623 ( .A0(n2271), .A1(n743), .B0(round[0]), .Y(n2270) );
  OAI21XL U1624 ( .A0(n2241), .A1(n182), .B0(n2242), .Y(n2240) );
  OAI21XL U1625 ( .A0(n136), .A1(n2244), .B0(n2245), .Y(n2242) );
  AOI2BB1X1 U1626 ( .A0N(n2267), .A1N(n2299), .B0(n730), .Y(n2478) );
  AOI21X1 U1627 ( .A0(n2289), .A1(n741), .B0(n329), .Y(n2286) );
  AOI21X1 U1628 ( .A0(n2322), .A1(n747), .B0(n328), .Y(n2458) );
  AOI21X1 U1629 ( .A0(n714), .A1(n712), .B0(round[2]), .Y(n2331) );
  INVX1 U1630 ( .A(n2325), .Y(n734) );
  INVX1 U1631 ( .A(n2329), .Y(n744) );
  NAND3BX1 U1632 ( .AN(n2321), .B(n2322), .C(n2323), .Y(n2319) );
  NAND3X1 U1633 ( .A(n2339), .B(n2340), .C(n2341), .Y(n2337) );
  OAI21XL U1634 ( .A0(n2344), .A1(n136), .B0(n40), .Y(n2339) );
  OAI21XL U1635 ( .A0(n2342), .A1(n2343), .B0(n183), .Y(n2341) );
  OAI21XL U1636 ( .A0(n2251), .A1(n2297), .B0(n2261), .Y(n2340) );
  AOI2BB1X1 U1637 ( .A0N(n2297), .A1N(n2284), .B0(round[0]), .Y(n2537) );
  AOI2BB1X1 U1638 ( .A0N(n2267), .A1N(n2447), .B0(n335), .Y(n2500) );
  XOR3X2 U1639 ( .A(n72), .B(n171), .C(n162), .Y(f3_A_32[31]) );
  OR2X2 U1640 ( .A(n328), .B(n335), .Y(n140) );
  INVX1 U1641 ( .A(n140), .Y(n2261) );
  INVX1 U1642 ( .A(n47), .Y(n738) );
  NOR3X1 U1643 ( .A(n726), .B(n182), .C(round[3]), .Y(n2477) );
  NAND2X1 U1644 ( .A(n131), .B(n328), .Y(n2346) );
  OAI21XL U1645 ( .A0(n182), .A1(n330), .B0(n2346), .Y(n2487) );
  NOR2X1 U1646 ( .A(n183), .B(n730), .Y(n2520) );
  INVX1 U1647 ( .A(n158), .Y(n589) );
  INVX1 U1648 ( .A(n161), .Y(n601) );
  INVX1 U1649 ( .A(n160), .Y(n597) );
  INVX1 U1650 ( .A(n172), .Y(n685) );
  INVX1 U1651 ( .A(n176), .Y(n681) );
  INVX1 U1652 ( .A(n166), .Y(n691) );
  INVX1 U1653 ( .A(n162), .Y(n695) );
  INVX1 U1654 ( .A(n165), .Y(n692) );
  INVX1 U1655 ( .A(n173), .Y(n684) );
  INVX1 U1656 ( .A(n174), .Y(n683) );
  INVX1 U1657 ( .A(n170), .Y(n687) );
  INVX1 U1658 ( .A(n167), .Y(n690) );
  INVX1 U1659 ( .A(n168), .Y(n689) );
  INVX1 U1660 ( .A(n157), .Y(n696) );
  INVX1 U1661 ( .A(n156), .Y(n698) );
  INVX1 U1662 ( .A(n181), .Y(n666) );
  INVX1 U1663 ( .A(inner_busy), .Y(n337) );
  XOR3X2 U1664 ( .A(SHA256_result[103]), .B(SHA256_result[116]), .C(
        SHA256_result[121]), .Y(f4_E_32[14]) );
  OAI211X1 U1665 ( .A0(n322), .A1(n782), .B0(n66), .C0(n1793), .Y(n2964) );
  NAND2X1 U1666 ( .A(H1[22]), .B(n254), .Y(n1793) );
  OAI211X1 U1667 ( .A0(n321), .A1(n787), .B0(n61), .C0(n1790), .Y(n2959) );
  NAND2X1 U1668 ( .A(H1[27]), .B(n254), .Y(n1790) );
  OAI211X1 U1669 ( .A0(n322), .A1(n778), .B0(n66), .C0(n1795), .Y(n2968) );
  NAND2X1 U1670 ( .A(H1[18]), .B(n253), .Y(n1795) );
  OAI211X1 U1671 ( .A0(n322), .A1(n777), .B0(n65), .C0(n1796), .Y(n2969) );
  NAND2X1 U1672 ( .A(H1[17]), .B(n253), .Y(n1796) );
  OAI211X1 U1673 ( .A0(n321), .A1(n789), .B0(n61), .C0(n1788), .Y(n2957) );
  NAND2X1 U1674 ( .A(H1[29]), .B(n254), .Y(n1788) );
  OAI211X1 U1675 ( .A0(n321), .A1(n788), .B0(n68), .C0(n1789), .Y(n2958) );
  NAND2X1 U1676 ( .A(H1[28]), .B(n254), .Y(n1789) );
  OAI211X1 U1677 ( .A0(n322), .A1(n781), .B0(n63), .C0(n1794), .Y(n2965) );
  NAND2X1 U1678 ( .A(H1[21]), .B(n254), .Y(n1794) );
  OAI211X1 U1679 ( .A0(n322), .A1(n775), .B0(n66), .C0(n1798), .Y(n2971) );
  NAND2X1 U1680 ( .A(H1[15]), .B(n253), .Y(n1798) );
  OAI211X1 U1681 ( .A0(n322), .A1(n773), .B0(n65), .C0(n1799), .Y(n2973) );
  NAND2X1 U1682 ( .A(H1[13]), .B(n253), .Y(n1799) );
  OAI211X1 U1683 ( .A0(n319), .A1(n813), .B0(n61), .C0(n1546), .Y(n2672) );
  NAND2X1 U1684 ( .A(H2[26]), .B(n258), .Y(n1546) );
  OAI211X1 U1685 ( .A0(n319), .A1(n806), .B0(n68), .C0(n1549), .Y(n2679) );
  NAND2X1 U1686 ( .A(H2[19]), .B(n258), .Y(n1549) );
  OAI211X1 U1687 ( .A0(n319), .A1(n805), .B0(n61), .C0(n1550), .Y(n2680) );
  NAND2X1 U1688 ( .A(H2[18]), .B(n258), .Y(n1550) );
  OAI211X1 U1689 ( .A0(n319), .A1(n804), .B0(n68), .C0(n1551), .Y(n2681) );
  NAND2X1 U1690 ( .A(H2[17]), .B(n258), .Y(n1551) );
  OAI211X1 U1691 ( .A0(n319), .A1(n816), .B0(n64), .C0(n1543), .Y(n2669) );
  NAND2X1 U1692 ( .A(H2[29]), .B(n260), .Y(n1543) );
  OAI211X1 U1693 ( .A0(n319), .A1(n809), .B0(n65), .C0(n1547), .Y(n2676) );
  NAND2X1 U1694 ( .A(H2[22]), .B(n258), .Y(n1547) );
  OAI211X1 U1695 ( .A0(n319), .A1(n802), .B0(n66), .C0(n1552), .Y(n2683) );
  NAND2X1 U1696 ( .A(H2[15]), .B(n258), .Y(n1552) );
  OAI211X1 U1697 ( .A0(n319), .A1(n801), .B0(n68), .C0(n1553), .Y(n2684) );
  NAND2X1 U1698 ( .A(H2[14]), .B(n257), .Y(n1553) );
  OAI211X1 U1699 ( .A0(n319), .A1(n800), .B0(n67), .C0(n1554), .Y(n2685) );
  NAND2X1 U1700 ( .A(H2[13]), .B(n257), .Y(n1554) );
  OAI211X1 U1701 ( .A0(n320), .A1(n799), .B0(n62), .C0(n1555), .Y(n2686) );
  NAND2X1 U1702 ( .A(H2[12]), .B(n257), .Y(n1555) );
  NAND2X1 U1703 ( .A(H2[5]), .B(n257), .Y(n1559) );
  OAI211X1 U1704 ( .A0(n318), .A1(n911), .B0(n63), .C0(n1525), .Y(n2638) );
  NAND2X1 U1705 ( .A(H6[27]), .B(n257), .Y(n1525) );
  OAI211X1 U1706 ( .A0(n318), .A1(n909), .B0(n61), .C0(n1527), .Y(n2640) );
  NAND2X1 U1707 ( .A(H6[25]), .B(n255), .Y(n1527) );
  OAI211X1 U1708 ( .A0(n318), .A1(n908), .B0(n62), .C0(n1528), .Y(n2641) );
  NAND2X1 U1709 ( .A(H6[24]), .B(n258), .Y(n1528) );
  OAI211X1 U1710 ( .A0(n318), .A1(n912), .B0(n68), .C0(n1524), .Y(n2637) );
  NAND2X1 U1711 ( .A(H6[28]), .B(n260), .Y(n1524) );
  OAI211X1 U1712 ( .A0(n318), .A1(n907), .B0(n67), .C0(n1529), .Y(n2642) );
  NAND2X1 U1713 ( .A(H6[23]), .B(n260), .Y(n1529) );
  OAI211X1 U1714 ( .A0(n318), .A1(n899), .B0(n65), .C0(n1532), .Y(n2650) );
  NAND2X1 U1715 ( .A(H6[15]), .B(n259), .Y(n1532) );
  OAI211X1 U1716 ( .A0(n318), .A1(n898), .B0(n63), .C0(n1533), .Y(n2651) );
  NAND2X1 U1717 ( .A(H6[14]), .B(n259), .Y(n1533) );
  OAI211X1 U1718 ( .A0(n321), .A1(n883), .B0(n66), .C0(n1601), .Y(n2769) );
  NAND2X1 U1719 ( .A(H5[24]), .B(n255), .Y(n1601) );
  OAI211X1 U1720 ( .A0(n321), .A1(n875), .B0(n65), .C0(n1603), .Y(n2777) );
  NAND2X1 U1721 ( .A(H5[16]), .B(n255), .Y(n1603) );
  OAI211X1 U1722 ( .A0(n321), .A1(n873), .B0(n67), .C0(n1604), .Y(n2779) );
  NAND2X1 U1723 ( .A(H5[14]), .B(n255), .Y(n1604) );
  OAI211X1 U1724 ( .A0(n322), .A1(n760), .B0(n58), .C0(n1805), .Y(n2986) );
  NAND2X1 U1725 ( .A(n91), .B(n253), .Y(n1805) );
  OAI211X1 U1726 ( .A0(n323), .A1(n506), .B0(n66), .C0(n1596), .Y(n2761) );
  NAND2X1 U1727 ( .A(H4[0]), .B(n255), .Y(n1596) );
  OAI211X1 U1728 ( .A0(n317), .A1(n853), .B0(n68), .C0(n1587), .Y(n2747) );
  NAND2X1 U1729 ( .A(H4[14]), .B(n256), .Y(n1587) );
  NAND2X1 U1730 ( .A(H4[5]), .B(n256), .Y(n1591) );
  NAND2X1 U1731 ( .A(H4[4]), .B(n255), .Y(n1592) );
  OAI211X1 U1732 ( .A0(n321), .A1(n785), .B0(n68), .C0(n1791), .Y(n2961) );
  NAND2X1 U1733 ( .A(H1[25]), .B(n254), .Y(n1791) );
  OAI211X1 U1734 ( .A0(n322), .A1(n784), .B0(n58), .C0(n1792), .Y(n2962) );
  NAND2X1 U1735 ( .A(H1[24]), .B(n254), .Y(n1792) );
  OAI211X1 U1736 ( .A0(n323), .A1(n495), .B0(n65), .C0(n1593), .Y(n2758) );
  NAND2X1 U1737 ( .A(H4[3]), .B(n255), .Y(n1593) );
  OAI211X1 U1738 ( .A0(n323), .A1(n502), .B0(n65), .C0(n1595), .Y(n2760) );
  NAND2X1 U1739 ( .A(H4[1]), .B(n255), .Y(n1595) );
  OAI211X1 U1740 ( .A0(n317), .A1(n863), .B0(n66), .C0(n1583), .Y(n2737) );
  NAND2X1 U1741 ( .A(H4[24]), .B(n256), .Y(n1583) );
  OAI211X1 U1742 ( .A0(n317), .A1(n857), .B0(n64), .C0(n1585), .Y(n2743) );
  NAND2X1 U1743 ( .A(H4[18]), .B(n256), .Y(n1585) );
  NAND2X1 U1744 ( .A(H1[2]), .B(n253), .Y(n1804) );
  OAI211X1 U1745 ( .A0(n324), .A1(n78), .B0(n68), .C0(n1594), .Y(n2759) );
  NAND2X1 U1746 ( .A(H4[2]), .B(n255), .Y(n1594) );
  OAI211X1 U1747 ( .A0(n35), .A1(n413), .B0(n369), .C0(n368), .Y(n2797) );
  AOI21X1 U1748 ( .A0(n214), .A1(SHA256_result[92]), .B0(n271), .Y(n369) );
  NAND2X1 U1749 ( .A(N1039), .B(n245), .Y(n368) );
  NAND2X1 U1750 ( .A(H4[28]), .B(n256), .Y(n1582) );
  NAND2X1 U1751 ( .A(H3[3]), .B(n256), .Y(n1579) );
  OAI211X1 U1752 ( .A0(n320), .A1(n846), .B0(n63), .C0(n1564), .Y(n2703) );
  NAND2X1 U1753 ( .A(H3[26]), .B(n257), .Y(n1564) );
  OAI211X1 U1754 ( .A0(n322), .A1(n776), .B0(n58), .C0(n1797), .Y(n2970) );
  NAND2X1 U1755 ( .A(H1[16]), .B(n253), .Y(n1797) );
  NAND2X1 U1756 ( .A(H1[10]), .B(n253), .Y(n1801) );
  OAI211X1 U1757 ( .A0(n321), .A1(n759), .B0(n61), .C0(n1787), .Y(n2955) );
  NAND2X1 U1758 ( .A(H1[31]), .B(n254), .Y(n1787) );
  OAI211X1 U1759 ( .A0(n319), .A1(n814), .B0(n61), .C0(n1545), .Y(n2671) );
  NAND2X1 U1760 ( .A(H2[27]), .B(n258), .Y(n1545) );
  OAI211X1 U1761 ( .A0(n319), .A1(n815), .B0(n66), .C0(n1544), .Y(n2670) );
  NAND2X1 U1762 ( .A(H2[28]), .B(n255), .Y(n1544) );
  OAI211X1 U1763 ( .A0(n319), .A1(n808), .B0(n58), .C0(n1548), .Y(n2677) );
  NAND2X1 U1764 ( .A(H2[21]), .B(n258), .Y(n1548) );
  OAI211X1 U1765 ( .A0(n320), .A1(n835), .B0(n62), .C0(n1571), .Y(n2714) );
  NAND2X1 U1766 ( .A(H3[15]), .B(n256), .Y(n1571) );
  OAI211X1 U1767 ( .A0(n318), .A1(n910), .B0(n65), .C0(n1526), .Y(n2639) );
  NAND2X1 U1768 ( .A(H6[26]), .B(n254), .Y(n1526) );
  OAI211X1 U1769 ( .A0(n318), .A1(n901), .B0(n62), .C0(n1530), .Y(n2648) );
  NAND2X1 U1770 ( .A(H6[17]), .B(n253), .Y(n1530) );
  OAI211X1 U1771 ( .A0(n318), .A1(n900), .B0(n65), .C0(n1531), .Y(n2649) );
  NAND2X1 U1772 ( .A(H6[16]), .B(n259), .Y(n1531) );
  OAI211X1 U1773 ( .A0(n321), .A1(n886), .B0(n62), .C0(n1599), .Y(n2766) );
  NAND2X1 U1774 ( .A(H5[27]), .B(n255), .Y(n1599) );
  OAI211X1 U1775 ( .A0(n321), .A1(n884), .B0(n57), .C0(n1600), .Y(n2768) );
  NAND2X1 U1776 ( .A(H5[25]), .B(n255), .Y(n1600) );
  OAI211X1 U1777 ( .A0(n319), .A1(n896), .B0(n57), .C0(n1534), .Y(n2653) );
  NAND2X1 U1778 ( .A(H6[12]), .B(n258), .Y(n1534) );
  OAI211X1 U1779 ( .A0(n321), .A1(n887), .B0(n66), .C0(n1598), .Y(n2765) );
  NAND2X1 U1780 ( .A(H5[28]), .B(n255), .Y(n1598) );
  OAI211X1 U1781 ( .A0(n321), .A1(n877), .B0(n61), .C0(n1602), .Y(n2775) );
  NAND2X1 U1782 ( .A(H5[18]), .B(n255), .Y(n1602) );
  OAI211X1 U1783 ( .A0(n320), .A1(n844), .B0(n57), .C0(n1565), .Y(n2705) );
  NAND2X1 U1784 ( .A(H3[24]), .B(n257), .Y(n1565) );
  OAI211X1 U1785 ( .A0(n321), .A1(n872), .B0(n67), .C0(n1605), .Y(n2780) );
  NAND2X1 U1786 ( .A(H5[13]), .B(n254), .Y(n1605) );
  OAI211X1 U1787 ( .A0(n323), .A1(n85), .B0(n64), .C0(n1561), .Y(n2697) );
  OAI211X1 U1788 ( .A0(n317), .A1(n944), .B0(n67), .C0(n1440), .Y(n2543) );
  NAND2X1 U1789 ( .A(H7[27]), .B(n260), .Y(n1440) );
  OAI211X1 U1790 ( .A0(n317), .A1(n942), .B0(n68), .C0(n1441), .Y(n2545) );
  NAND2X1 U1791 ( .A(H7[25]), .B(n260), .Y(n1441) );
  OAI211X1 U1792 ( .A0(n320), .A1(n837), .B0(n61), .C0(n1569), .Y(n2712) );
  NAND2X1 U1793 ( .A(H3[17]), .B(n256), .Y(n1569) );
  OAI211X1 U1794 ( .A0(n320), .A1(n836), .B0(n65), .C0(n1570), .Y(n2713) );
  NAND2X1 U1795 ( .A(H3[16]), .B(n252), .Y(n1570) );
  NAND2X1 U1796 ( .A(H3[10]), .B(n254), .Y(n1575) );
  OAI211X1 U1797 ( .A0(n317), .A1(n947), .B0(n58), .C0(n1438), .Y(n2540) );
  NAND2X1 U1798 ( .A(H7[30]), .B(n260), .Y(n1438) );
  OAI211X1 U1799 ( .A0(n317), .A1(n945), .B0(n66), .C0(n1439), .Y(n2542) );
  NAND2X1 U1800 ( .A(H7[28]), .B(n259), .Y(n1439) );
  OAI211X1 U1801 ( .A0(n317), .A1(n932), .B0(n57), .C0(n1446), .Y(n2555) );
  NAND2X1 U1802 ( .A(H7[15]), .B(n260), .Y(n1446) );
  OAI211X1 U1803 ( .A0(n318), .A1(n931), .B0(n57), .C0(n1447), .Y(n2556) );
  NAND2X1 U1804 ( .A(H7[14]), .B(n260), .Y(n1447) );
  OAI211X1 U1805 ( .A0(n320), .A1(n849), .B0(n57), .C0(n1563), .Y(n2700) );
  NAND2X1 U1806 ( .A(H3[29]), .B(n257), .Y(n1563) );
  OAI211X1 U1807 ( .A0(n320), .A1(n842), .B0(n68), .C0(n1566), .Y(n2707) );
  NAND2X1 U1808 ( .A(H3[22]), .B(n255), .Y(n1566) );
  OAI211X1 U1809 ( .A0(n317), .A1(n834), .B0(n68), .C0(n1572), .Y(n2715) );
  NAND2X1 U1810 ( .A(H3[14]), .B(n257), .Y(n1572) );
  OAI211X1 U1811 ( .A0(n317), .A1(n832), .B0(n63), .C0(n1574), .Y(n2717) );
  NAND2X1 U1812 ( .A(H3[12]), .B(n254), .Y(n1574) );
  NAND2X1 U1813 ( .A(H3[5]), .B(n253), .Y(n1577) );
  OAI211X1 U1814 ( .A0(n320), .A1(n819), .B0(n58), .C0(n1562), .Y(n2698) );
  NAND2X1 U1815 ( .A(H3[31]), .B(n257), .Y(n1562) );
  OAI211X1 U1816 ( .A0(n320), .A1(n839), .B0(n61), .C0(n1567), .Y(n2710) );
  NAND2X1 U1817 ( .A(H3[19]), .B(n256), .Y(n1567) );
  OAI211X1 U1818 ( .A0(n320), .A1(n838), .B0(n58), .C0(n1568), .Y(n2711) );
  NAND2X1 U1819 ( .A(H3[18]), .B(n252), .Y(n1568) );
  OAI211X1 U1820 ( .A0(n317), .A1(n833), .B0(n64), .C0(n1573), .Y(n2716) );
  NAND2X1 U1821 ( .A(H3[13]), .B(n259), .Y(n1573) );
  NAND2X1 U1822 ( .A(H7[3]), .B(n258), .Y(n1452) );
  NAND2X1 U1823 ( .A(H7[4]), .B(n260), .Y(n1451) );
  OAI211X1 U1824 ( .A0(n321), .A1(n864), .B0(n64), .C0(n1597), .Y(n2762) );
  INVX1 U1825 ( .A(SHA256_result[95]), .Y(n864) );
  NAND2X1 U1826 ( .A(H5[31]), .B(n255), .Y(n1597) );
  OAI211X1 U1827 ( .A0(n322), .A1(n858), .B0(n68), .C0(n1584), .Y(n2742) );
  INVX1 U1828 ( .A(n147), .Y(n858) );
  NAND2X1 U1829 ( .A(H4[19]), .B(n256), .Y(n1584) );
  OAI211X1 U1830 ( .A0(n320), .A1(n856), .B0(n57), .C0(n1586), .Y(n2744) );
  INVX1 U1831 ( .A(n148), .Y(n856) );
  NAND2X1 U1832 ( .A(H4[17]), .B(n256), .Y(n1586) );
  OAI211X1 U1833 ( .A0(n317), .A1(n851), .B0(n65), .C0(n1588), .Y(n2749) );
  NAND2X1 U1834 ( .A(H4[12]), .B(n256), .Y(n1588) );
  OAI211X1 U1835 ( .A0(n322), .A1(n699), .B0(n58), .C0(n1861), .Y(n3020) );
  INVX1 U1836 ( .A(n155), .Y(n699) );
  NAND2X1 U1837 ( .A(H0[30]), .B(n253), .Y(n1861) );
  OAI211X1 U1838 ( .A0(n322), .A1(n698), .B0(n65), .C0(n1862), .Y(n3021) );
  NAND2X1 U1839 ( .A(H0[29]), .B(n253), .Y(n1862) );
  OAI211X1 U1840 ( .A0(n323), .A1(n696), .B0(n66), .C0(n1863), .Y(n3023) );
  NAND2X1 U1841 ( .A(H0[27]), .B(n252), .Y(n1863) );
  OAI211X1 U1842 ( .A0(n323), .A1(n592), .B0(n67), .C0(n1864), .Y(n3025) );
  INVX1 U1843 ( .A(n159), .Y(n592) );
  NAND2X1 U1844 ( .A(H0[25]), .B(n252), .Y(n1864) );
  OAI211X1 U1845 ( .A0(n323), .A1(n693), .B0(n61), .C0(n1865), .Y(n3031) );
  INVX1 U1846 ( .A(n164), .Y(n693) );
  NAND2X1 U1847 ( .A(H0[19]), .B(n252), .Y(n1865) );
  OAI211X1 U1848 ( .A0(n323), .A1(n690), .B0(n65), .C0(n1866), .Y(n3034) );
  NAND2X1 U1849 ( .A(H0[16]), .B(n252), .Y(n1866) );
  OAI211X1 U1850 ( .A0(n323), .A1(n689), .B0(n58), .C0(n1867), .Y(n3035) );
  NAND2X1 U1851 ( .A(H0[15]), .B(n252), .Y(n1867) );
  OAI211X1 U1852 ( .A0(n323), .A1(n688), .B0(n68), .C0(n1868), .Y(n3036) );
  INVX1 U1853 ( .A(n169), .Y(n688) );
  NAND2X1 U1854 ( .A(H0[14]), .B(n252), .Y(n1868) );
  OAI211X1 U1855 ( .A0(n323), .A1(n687), .B0(n65), .C0(n1869), .Y(n3037) );
  NAND2X1 U1856 ( .A(H0[13]), .B(n252), .Y(n1869) );
  OAI211X1 U1857 ( .A0(n323), .A1(n684), .B0(n68), .C0(n1870), .Y(n3040) );
  NAND2X1 U1858 ( .A(H0[10]), .B(n252), .Y(n1870) );
  OAI211X1 U1859 ( .A0(n323), .A1(n683), .B0(n66), .C0(n1871), .Y(n3041) );
  NAND2X1 U1860 ( .A(H0[9]), .B(n252), .Y(n1871) );
  OAI211X1 U1861 ( .A0(n323), .A1(n680), .B0(n63), .C0(n1872), .Y(n3044) );
  INVX1 U1862 ( .A(n177), .Y(n680) );
  NAND2X1 U1863 ( .A(H0[6]), .B(n252), .Y(n1872) );
  OAI211X1 U1864 ( .A0(n323), .A1(n666), .B0(n62), .C0(n1874), .Y(n3048) );
  NAND2X1 U1865 ( .A(H0[2]), .B(n252), .Y(n1874) );
  OAI211X1 U1866 ( .A0(n323), .A1(n93), .B0(n61), .C0(n1876), .Y(n3050) );
  NAND2X1 U1867 ( .A(H0[0]), .B(n252), .Y(n1876) );
  XOR3X2 U1868 ( .A(SHA256_result[101]), .B(SHA256_result[114]), .C(
        SHA256_result[119]), .Y(f4_E_32[12]) );
  OAI21XL U1869 ( .A0(n705), .A1(n946), .B0(n1460), .Y(n2573) );
  AOI22X1 U1870 ( .A0(N1104), .A1(n237), .B0(SHA256_result[61]), .B1(n10), .Y(
        n1460) );
  XOR3X2 U1871 ( .A(SHA256_result[99]), .B(SHA256_result[112]), .C(n146), .Y(
        f4_E_32[10]) );
  XOR3X2 U1872 ( .A(n74), .B(SHA256_result[110]), .C(n147), .Y(f4_E_32[8]) );
  XOR3X2 U1873 ( .A(SHA256_result[98]), .B(n149), .C(SHA256_result[116]), .Y(
        f4_E_32[9]) );
  OAI2BB2X1 U1874 ( .B0(n327), .B1(n700), .A0N(H0[31]), .A1N(n261), .Y(n3019)
         );
  OAI2BB2X1 U1875 ( .B0(n327), .B1(n697), .A0N(H0[28]), .A1N(n261), .Y(n3022)
         );
  OAI2BB2X1 U1876 ( .B0(n327), .B1(n786), .A0N(H1[26]), .A1N(n262), .Y(n2960)
         );
  OAI2BB2X1 U1877 ( .B0(n327), .B1(n779), .A0N(H1[19]), .A1N(n262), .Y(n2967)
         );
  OAI2BB2X1 U1878 ( .B0(n327), .B1(n774), .A0N(H1[14]), .A1N(n261), .Y(n2972)
         );
  OAI2BB2X1 U1879 ( .B0(n327), .B1(n772), .A0N(H1[12]), .A1N(n262), .Y(n2974)
         );
  OAI2BB2X1 U1880 ( .B0(n327), .B1(n765), .A0N(H1[5]), .A1N(n261), .Y(n2981)
         );
  OAI2BB2X1 U1881 ( .B0(n327), .B1(n811), .A0N(H2[24]), .A1N(n263), .Y(n2674)
         );
  OAI2BB2X1 U1882 ( .B0(n327), .B1(n803), .A0N(H2[16]), .A1N(n264), .Y(n2682)
         );
  OAI2BB2X1 U1883 ( .B0(n327), .B1(n818), .A0N(H2[31]), .A1N(n265), .Y(n2667)
         );
  OAI2BB2X1 U1884 ( .B0(n327), .B1(n914), .A0N(H6[30]), .A1N(n264), .Y(n2635)
         );
  OAI2BB2X1 U1885 ( .B0(n327), .B1(n906), .A0N(H6[22]), .A1N(n265), .Y(n2643)
         );
  OAI2BB2X1 U1886 ( .B0(n327), .B1(n905), .A0N(H6[21]), .A1N(n265), .Y(n2644)
         );
  OAI2BB2X1 U1887 ( .B0(n327), .B1(n885), .A0N(H5[26]), .A1N(n264), .Y(n2767)
         );
  OAI2BB2X1 U1888 ( .B0(n327), .B1(n876), .A0N(H5[17]), .A1N(n263), .Y(n2776)
         );
  OAI2BB2X1 U1889 ( .B0(n327), .B1(n882), .A0N(H5[23]), .A1N(n263), .Y(n2770)
         );
  OAI2BB2X1 U1890 ( .B0(n327), .B1(n874), .A0N(H5[15]), .A1N(n263), .Y(n2778)
         );
  OAI2BB2X1 U1891 ( .B0(n327), .B1(n871), .A0N(H5[12]), .A1N(n263), .Y(n2781)
         );
  OAI2BB2X1 U1892 ( .B0(n327), .B1(n862), .A0N(H4[23]), .A1N(n265), .Y(n2738)
         );
  OAI2BB2X1 U1893 ( .B0(n327), .B1(n861), .A0N(H4[22]), .A1N(n264), .Y(n2739)
         );
  OAI2BB2X1 U1894 ( .B0(n327), .B1(n855), .A0N(H4[16]), .A1N(n264), .Y(n2745)
         );
  OAI2BB2X1 U1895 ( .B0(n327), .B1(n852), .A0N(H4[13]), .A1N(n264), .Y(n2748)
         );
  OAI2BB2X1 U1896 ( .B0(n327), .B1(n790), .A0N(H1[30]), .A1N(n262), .Y(n2956)
         );
  OAI2BB2X1 U1897 ( .B0(n327), .B1(n783), .A0N(H1[23]), .A1N(n262), .Y(n2963)
         );
  OAI2BB2X1 U1898 ( .B0(n327), .B1(n780), .A0N(H1[20]), .A1N(n262), .Y(n2966)
         );
  OAI2BB2X1 U1899 ( .B0(n327), .B1(n763), .A0N(H1[3]), .A1N(n261), .Y(n2983)
         );
  OAI2BB2X1 U1900 ( .B0(n327), .B1(n847), .A0N(H3[27]), .A1N(n252), .Y(n2702)
         );
  OAI2BB2X1 U1901 ( .B0(n327), .B1(n848), .A0N(H3[28]), .A1N(n255), .Y(n2701)
         );
  OAI2BB2X1 U1902 ( .B0(n327), .B1(n812), .A0N(H2[25]), .A1N(n258), .Y(n2673)
         );
  OAI2BB2X1 U1903 ( .B0(n327), .B1(n817), .A0N(H2[30]), .A1N(n252), .Y(n2668)
         );
  OAI2BB2X1 U1904 ( .B0(n327), .B1(n810), .A0N(H2[23]), .A1N(n263), .Y(n2675)
         );
  OAI2BB2X1 U1905 ( .B0(n327), .B1(n807), .A0N(H2[20]), .A1N(n261), .Y(n2678)
         );
  OAI2BB2X1 U1906 ( .B0(n327), .B1(n903), .A0N(H6[19]), .A1N(n265), .Y(n2646)
         );
  OAI2BB2X1 U1907 ( .B0(n327), .B1(n902), .A0N(H6[18]), .A1N(n265), .Y(n2647)
         );
  OAI2BB2X1 U1908 ( .B0(n327), .B1(n840), .A0N(H3[20]), .A1N(n265), .Y(n2709)
         );
  OAI2BB2X1 U1909 ( .B0(n327), .B1(n915), .A0N(H6[31]), .A1N(n264), .Y(n2634)
         );
  OAI2BB2X1 U1910 ( .B0(n327), .B1(n913), .A0N(H6[29]), .A1N(n264), .Y(n2636)
         );
  OAI2BB2X1 U1911 ( .B0(n327), .B1(n904), .A0N(H6[20]), .A1N(n265), .Y(n2645)
         );
  OAI2BB2X1 U1912 ( .B0(n327), .B1(n897), .A0N(H6[13]), .A1N(n265), .Y(n2652)
         );
  OAI2BB2X1 U1913 ( .B0(n327), .B1(n878), .A0N(H5[19]), .A1N(n263), .Y(n2774)
         );
  OAI2BB2X1 U1914 ( .B0(n327), .B1(n889), .A0N(H5[30]), .A1N(n264), .Y(n2763)
         );
  OAI2BB2X1 U1915 ( .B0(n327), .B1(n888), .A0N(H5[29]), .A1N(n264), .Y(n2764)
         );
  OAI2BB2X1 U1916 ( .B0(n327), .B1(n881), .A0N(H5[22]), .A1N(n263), .Y(n2771)
         );
  OAI2BB2X1 U1917 ( .B0(n327), .B1(n880), .A0N(H5[21]), .A1N(n263), .Y(n2772)
         );
  OAI2BB2X1 U1918 ( .B0(n327), .B1(n879), .A0N(H5[20]), .A1N(n263), .Y(n2773)
         );
  OAI2BB2X1 U1919 ( .B0(n327), .B1(n841), .A0N(H3[21]), .A1N(n265), .Y(n2708)
         );
  OAI2BB2X1 U1920 ( .B0(n327), .B1(n943), .A0N(H7[26]), .A1N(n262), .Y(n2544)
         );
  OAI2BB2X1 U1921 ( .B0(n327), .B1(n936), .A0N(H7[19]), .A1N(n263), .Y(n2551)
         );
  OAI2BB2X1 U1922 ( .B0(n327), .B1(n935), .A0N(H7[18]), .A1N(n263), .Y(n2552)
         );
  OAI2BB2X1 U1923 ( .B0(n327), .B1(n934), .A0N(H7[17]), .A1N(n263), .Y(n2553)
         );
  OAI2BB2X1 U1924 ( .B0(n327), .B1(n933), .A0N(H7[16]), .A1N(n263), .Y(n2554)
         );
  OAI2BB2X1 U1925 ( .B0(n327), .B1(n919), .A0N(H7[2]), .A1N(n264), .Y(n2568)
         );
  OAI2BB2X1 U1926 ( .B0(n327), .B1(n822), .A0N(H3[2]), .A1N(n265), .Y(n2727)
         );
  OAI2BB2X1 U1927 ( .B0(n327), .B1(n946), .A0N(H7[29]), .A1N(n262), .Y(n2541)
         );
  OAI2BB2X1 U1928 ( .B0(n327), .B1(n937), .A0N(H7[20]), .A1N(n262), .Y(n2550)
         );
  OAI2BB2X1 U1929 ( .B0(n327), .B1(n930), .A0N(H7[13]), .A1N(n263), .Y(n2557)
         );
  OAI2BB2X1 U1930 ( .B0(n327), .B1(n929), .A0N(H7[12]), .A1N(n263), .Y(n2558)
         );
  OAI2BB2X1 U1931 ( .B0(n327), .B1(n850), .A0N(H3[30]), .A1N(n255), .Y(n2699)
         );
  OAI2BB2X1 U1932 ( .B0(n327), .B1(n843), .A0N(H3[23]), .A1N(n265), .Y(n2706)
         );
  OAI2BB2X1 U1933 ( .B0(n327), .B1(n916), .A0N(H7[31]), .A1N(n262), .Y(n2539)
         );
  OAI2BB2X1 U1934 ( .B0(n327), .B1(n845), .A0N(H3[25]), .A1N(n265), .Y(n2704)
         );
  XOR3X2 U1935 ( .A(SHA256_result[127]), .B(n150), .C(n148), .Y(f4_E_32[6]) );
  OAI21XL U1936 ( .A0(n327), .A1(n605), .B0(n604), .Y(n3028) );
  NAND2X1 U1937 ( .A(H0[22]), .B(n259), .Y(n604) );
  OAI2BB2X1 U1938 ( .B0(n327), .B1(n681), .A0N(H0[7]), .A1N(n261), .Y(n3043)
         );
  OAI2BB2X1 U1939 ( .B0(n327), .B1(n695), .A0N(H0[21]), .A1N(n261), .Y(n3029)
         );
  OAI2BB2X1 U1940 ( .B0(n327), .B1(n692), .A0N(H0[18]), .A1N(n261), .Y(n3032)
         );
  OAI21XL U1941 ( .A0(n327), .A1(n418), .B0(n417), .Y(n2734) );
  NAND2X1 U1942 ( .A(H4[27]), .B(n259), .Y(n417) );
  OAI21XL U1943 ( .A0(n327), .A1(n426), .B0(n425), .Y(n2736) );
  NAND2X1 U1944 ( .A(H4[25]), .B(n259), .Y(n425) );
  OAI2BB2X1 U1945 ( .B0(n327), .B1(n860), .A0N(H4[21]), .A1N(n264), .Y(n2740)
         );
  INVX1 U1946 ( .A(n146), .Y(n860) );
  OAI2BB2X1 U1947 ( .B0(n327), .B1(n859), .A0N(H4[20]), .A1N(n264), .Y(n2741)
         );
  INVX1 U1948 ( .A(SHA256_result[116]), .Y(n859) );
  OAI2BB2X1 U1949 ( .B0(n327), .B1(n854), .A0N(H4[15]), .A1N(n264), .Y(n2746)
         );
  OAI2BB2X1 U1950 ( .B0(n327), .B1(n694), .A0N(H0[20]), .A1N(n262), .Y(n3030)
         );
  INVX1 U1951 ( .A(n163), .Y(n694) );
  OAI21XL U1952 ( .A0(n327), .A1(n511), .B0(n510), .Y(n2730) );
  NAND2X1 U1953 ( .A(H4[31]), .B(n253), .Y(n510) );
  OAI2BB2X1 U1954 ( .B0(n327), .B1(n686), .A0N(H0[12]), .A1N(n261), .Y(n3038)
         );
  INVX1 U1955 ( .A(n171), .Y(n686) );
  INVX1 U1956 ( .A(n175), .Y(n682) );
  OAI21XL U1957 ( .A0(n327), .A1(n400), .B0(n356), .Y(n2661) );
  OAI21XL U1958 ( .A0(n327), .A1(n106), .B0(n391), .Y(n2793) );
  OAI21XL U1959 ( .A0(n327), .A1(n116), .B0(n388), .Y(n2792) );
  OAI21XL U1960 ( .A0(n327), .A1(n397), .B0(n378), .Y(n2788) );
  OAI21XL U1961 ( .A0(n327), .A1(n399), .B0(n381), .Y(n2789) );
  AOI21X1 U1962 ( .A0(SHA256_result[124]), .A1(n212), .B0(n275), .Y(n416) );
  OAI21XL U1963 ( .A0(n327), .A1(n422), .B0(n421), .Y(n2735) );
  NAND2X1 U1964 ( .A(H4[26]), .B(n257), .Y(n421) );
  OAI21XL U1965 ( .A0(n327), .A1(n410), .B0(n409), .Y(n2732) );
  NAND2X1 U1966 ( .A(H4[29]), .B(n254), .Y(n409) );
  XOR3X2 U1967 ( .A(SHA256_result[100]), .B(n148), .C(SHA256_result[118]), .Y(
        f4_E_32[11]) );
  OAI21XL U1968 ( .A0(n189), .A1(n848), .B0(n1694), .Y(n2861) );
  AOI22X1 U1969 ( .A0(N975), .A1(n237), .B0(SHA256_result[188]), .B1(n10), .Y(
        n1694) );
  OAI21XL U1970 ( .A0(n327), .A1(n461), .B0(n460), .Y(n2750) );
  NAND2X1 U1971 ( .A(H4[11]), .B(n259), .Y(n460) );
  OAI21XL U1972 ( .A0(n327), .A1(n479), .B0(n478), .Y(n2754) );
  NAND2X1 U1973 ( .A(H4[7]), .B(n259), .Y(n478) );
  OAI21XL U1974 ( .A0(n186), .A1(n913), .B0(n1495), .Y(n2605) );
  AOI22X1 U1975 ( .A0(N1072), .A1(n235), .B0(SHA256_result[93]), .B1(n10), .Y(
        n1495) );
  OAI21XL U1976 ( .A0(n186), .A1(n888), .B0(n1612), .Y(n2796) );
  OAI21XL U1977 ( .A0(n327), .A1(n404), .B0(n361), .Y(n2663) );
  OAI21XL U1978 ( .A0(n327), .A1(n519), .B0(n518), .Y(n2695) );
  OAI21XL U1979 ( .A0(n327), .A1(n589), .B0(n588), .Y(n3024) );
  NAND2X1 U1980 ( .A(H0[26]), .B(n254), .Y(n588) );
  OAI21XL U1981 ( .A0(n327), .A1(n597), .B0(n596), .Y(n3026) );
  NAND2X1 U1982 ( .A(H0[24]), .B(n260), .Y(n596) );
  OAI21XL U1983 ( .A0(n327), .A1(n601), .B0(n600), .Y(n3027) );
  NAND2X1 U1984 ( .A(H0[23]), .B(n260), .Y(n600) );
  OAI21XL U1985 ( .A0(n327), .A1(n523), .B0(n522), .Y(n2696) );
  OAI21XL U1986 ( .A0(n327), .A1(n88), .B0(n530), .Y(n2922) );
  OAI21XL U1987 ( .A0(n327), .A1(n656), .B0(n655), .Y(n3046) );
  NAND2X1 U1988 ( .A(H0[4]), .B(n260), .Y(n655) );
  OAI21XL U1989 ( .A0(n327), .A1(n661), .B0(n660), .Y(n3047) );
  NAND2X1 U1990 ( .A(H0[3]), .B(n260), .Y(n660) );
  OAI21XL U1991 ( .A0(n327), .A1(n465), .B0(n464), .Y(n2751) );
  NAND2X1 U1992 ( .A(H4[10]), .B(n259), .Y(n464) );
  OAI21XL U1993 ( .A0(n327), .A1(n474), .B0(n473), .Y(n2753) );
  NAND2X1 U1994 ( .A(H4[8]), .B(n253), .Y(n473) );
  NAND2X1 U1995 ( .A(H4[9]), .B(n256), .Y(n1589) );
  INVX1 U1996 ( .A(n152), .Y(n469) );
  NAND2X1 U1997 ( .A(H4[6]), .B(n256), .Y(n1590) );
  INVX1 U1998 ( .A(n154), .Y(n483) );
  NAND2X1 U1999 ( .A(H0[5]), .B(n252), .Y(n1873) );
  INVX1 U2000 ( .A(n178), .Y(n651) );
  NAND2X1 U2001 ( .A(H0[1]), .B(n252), .Y(n1875) );
  NOR2X1 U2002 ( .A(n317), .B(n102), .Y(n670) );
  NAND2X1 U2003 ( .A(H4[30]), .B(n256), .Y(n1581) );
  INVX1 U2004 ( .A(n145), .Y(n396) );
  NAND3X1 U2005 ( .A(n431), .B(n430), .C(n429), .Y(n2833) );
  NAND2XL U2006 ( .A(next_E[24]), .B(n11), .Y(n430) );
  OAI211X1 U2007 ( .A0(n12), .A1(n445), .B0(n444), .C0(n443), .Y(n2839) );
  INVXL U2008 ( .A(next_E[18]), .Y(n445) );
  OAI211X1 U2009 ( .A0(n31), .A1(n455), .B0(n454), .C0(n453), .Y(n2843) );
  INVXL U2010 ( .A(next_E[14]), .Y(n455) );
  AOI21X1 U2011 ( .A0(n213), .A1(SHA256_result[110]), .B0(n276), .Y(n454) );
  AOI2BB2X1 U2012 ( .B0(n193), .B1(SHA256_result[112]), .A0N(n12), .A1N(n449), 
        .Y(n450) );
  OAI2BB1X1 U2013 ( .A0N(SHA256_result[192]), .A1N(n70), .B0(n574), .Y(
        f2_ABC_32[0]) );
  OAI21XL U2014 ( .A0(n70), .A1(SHA256_result[192]), .B0(n90), .Y(n574) );
  OAI211X1 U2015 ( .A0(n761), .A1(n20), .B0(n527), .C0(n526), .Y(n2920) );
  OAI211X1 U2016 ( .A0(n15), .A1(n418), .B0(n371), .C0(n370), .Y(n2798) );
  NAND2X1 U2017 ( .A(N1038), .B(n245), .Y(n370) );
  OAI211X1 U2018 ( .A0(n33), .A1(n426), .B0(n373), .C0(n372), .Y(n2800) );
  NAND2X1 U2019 ( .A(N1036), .B(n245), .Y(n372) );
  AOI21X1 U2020 ( .A0(n213), .A1(SHA256_result[89]), .B0(n271), .Y(n373) );
  NAND2X1 U2021 ( .A(N1043), .B(n245), .Y(n367) );
  OAI211XL U2022 ( .A0(n27), .A1(n116), .B0(n365), .C0(n364), .Y(n2633) );
  NAND2X1 U2023 ( .A(N1048), .B(n245), .Y(n355) );
  NAND2X1 U2024 ( .A(N1046), .B(n245), .Y(n360) );
  OAI211X1 U2025 ( .A0(n25), .A1(n403), .B0(n363), .C0(n362), .Y(n2632) );
  NAND2XL U2026 ( .A(SHA256_result[34]), .B(n197), .Y(n363) );
  NAND2X1 U2027 ( .A(N1045), .B(n245), .Y(n362) );
  OAI211X1 U2028 ( .A0(n19), .A1(n461), .B0(n375), .C0(n374), .Y(n2814) );
  OAI211X1 U2029 ( .A0(n13), .A1(n479), .B0(n377), .C0(n376), .Y(n2818) );
  OAI211X1 U2030 ( .A0(n21), .A1(n506), .B0(n393), .C0(n392), .Y(n2825) );
  OAI211X1 U2031 ( .A0(n24), .A1(n487), .B0(n380), .C0(n379), .Y(n2820) );
  OAI211X1 U2032 ( .A0(n20), .A1(n491), .B0(n383), .C0(n382), .Y(n2821) );
  OAI211X1 U2033 ( .A0(n30), .A1(n495), .B0(n385), .C0(n384), .Y(n2822) );
  OAI211X1 U2034 ( .A0(n22), .A1(n502), .B0(n390), .C0(n389), .Y(n2824) );
  OAI211X1 U2035 ( .A0(n13), .A1(n78), .B0(n387), .C0(n386), .Y(n2823) );
  OAI211X1 U2036 ( .A0(n33), .A1(n482), .B0(n481), .C0(n480), .Y(n2850) );
  NAND2XL U2037 ( .A(SHA256_result[103]), .B(n196), .Y(n481) );
  OAI211X1 U2038 ( .A0(n32), .A1(n490), .B0(n489), .C0(n488), .Y(n2852) );
  NAND2X1 U2039 ( .A(N984), .B(n247), .Y(n489) );
  OAI211X1 U2040 ( .A0(n14), .A1(n494), .B0(n493), .C0(n492), .Y(n2853) );
  NAND2X1 U2041 ( .A(N983), .B(n247), .Y(n493) );
  OAI211X1 U2042 ( .A0(n36), .A1(n498), .B0(n497), .C0(n496), .Y(n2854) );
  NAND2X1 U2043 ( .A(N982), .B(n247), .Y(n497) );
  AOI21XL U2044 ( .A0(SHA256_result[99]), .A1(n211), .B0(n278), .Y(n496) );
  OAI211X1 U2045 ( .A0(n13), .A1(n501), .B0(n500), .C0(n499), .Y(n2855) );
  NAND2X1 U2046 ( .A(N981), .B(n247), .Y(n500) );
  AOI21XL U2047 ( .A0(SHA256_result[98]), .A1(n211), .B0(n272), .Y(n499) );
  OAI211X1 U2048 ( .A0(n12), .A1(n505), .B0(n504), .C0(n503), .Y(n2856) );
  NAND2X1 U2049 ( .A(N980), .B(n247), .Y(n504) );
  AOI21XL U2050 ( .A0(n74), .A1(n211), .B0(n272), .Y(n503) );
  OAI211X1 U2051 ( .A0(n22), .A1(n509), .B0(n508), .C0(n507), .Y(n2857) );
  INVX1 U2052 ( .A(next_E[0]), .Y(n509) );
  OAI211X1 U2053 ( .A0(n31), .A1(n763), .B0(n521), .C0(n520), .Y(n2918) );
  OAI211X1 U2054 ( .A0(n17), .A1(n762), .B0(n525), .C0(n524), .Y(n2919) );
  OAI211X1 U2055 ( .A0(n23), .A1(n760), .B0(n529), .C0(n528), .Y(n2921) );
  NAND2X1 U2056 ( .A(N915), .B(n247), .Y(n528) );
  OAI21XL U2057 ( .A0(n705), .A1(n943), .B0(n1463), .Y(n2576) );
  AOI22X1 U2058 ( .A0(N1101), .A1(n237), .B0(SHA256_result[58]), .B1(n11), .Y(
        n1463) );
  OAI21XL U2059 ( .A0(n705), .A1(n937), .B0(n1469), .Y(n2582) );
  OAI2BB1X1 U2060 ( .A0N(SHA256_result[201]), .A1N(n174), .B0(n565), .Y(
        f2_ABC_32[9]) );
  OAI21XL U2061 ( .A0(SHA256_result[201]), .A1(n174), .B0(SHA256_result[169]), 
        .Y(n565) );
  OAI2BB1X1 U2062 ( .A0N(SHA256_result[203]), .A1N(n172), .B0(n563), .Y(
        f2_ABC_32[11]) );
  OAI21XL U2063 ( .A0(SHA256_result[203]), .A1(n172), .B0(SHA256_result[171]), 
        .Y(n563) );
  OAI2BB1X1 U2064 ( .A0N(SHA256_result[199]), .A1N(n176), .B0(n567), .Y(
        f2_ABC_32[7]) );
  OAI21XL U2065 ( .A0(SHA256_result[199]), .A1(n176), .B0(SHA256_result[167]), 
        .Y(n567) );
  OAI2BB1X1 U2066 ( .A0N(SHA256_result[198]), .A1N(n177), .B0(n568), .Y(
        f2_ABC_32[6]) );
  OAI21XL U2067 ( .A0(SHA256_result[198]), .A1(n177), .B0(SHA256_result[166]), 
        .Y(n568) );
  OAI2BB1X1 U2068 ( .A0N(SHA256_result[200]), .A1N(n175), .B0(n566), .Y(
        f2_ABC_32[8]) );
  OAI21XL U2069 ( .A0(SHA256_result[200]), .A1(n175), .B0(SHA256_result[168]), 
        .Y(n566) );
  OAI2BB1X1 U2070 ( .A0N(SHA256_result[202]), .A1N(n173), .B0(n564), .Y(
        f2_ABC_32[10]) );
  OAI21XL U2071 ( .A0(SHA256_result[202]), .A1(n173), .B0(SHA256_result[170]), 
        .Y(n564) );
  OAI2BB1X1 U2072 ( .A0N(SHA256_result[196]), .A1N(n179), .B0(n570), .Y(
        f2_ABC_32[4]) );
  OAI21XL U2073 ( .A0(SHA256_result[196]), .A1(n179), .B0(SHA256_result[164]), 
        .Y(n570) );
  XOR3X2 U2074 ( .A(n77), .B(SHA256_result[110]), .C(n73), .Y(f4_E_32[21]) );
  XOR3X2 U2075 ( .A(SHA256_result[107]), .B(SHA256_result[120]), .C(
        SHA256_result[125]), .Y(f4_E_32[18]) );
  XOR3X2 U2076 ( .A(n152), .B(SHA256_result[118]), .C(n73), .Y(f4_E_32[16]) );
  XOR3X2 U2077 ( .A(n151), .B(SHA256_result[119]), .C(SHA256_result[124]), .Y(
        f4_E_32[17]) );
  MX2X1 U2078 ( .A(SHA256_result[48]), .B(SHA256_result[80]), .S0(
        SHA256_result[112]), .Y(f1_EFG_32[16]) );
  MX2X1 U2079 ( .A(SHA256_result[50]), .B(SHA256_result[82]), .S0(
        SHA256_result[114]), .Y(f1_EFG_32[18]) );
  XOR3X2 U2080 ( .A(n164), .B(n175), .C(SHA256_result[252]), .Y(f3_A_32[6]) );
  XOR3X2 U2081 ( .A(n37), .B(n172), .C(SHA256_result[255]), .Y(f3_A_32[9]) );
  XOR3X2 U2082 ( .A(SHA256_result[121]), .B(n150), .C(n145), .Y(f4_E_32[19])
         );
  XOR3X2 U2083 ( .A(n154), .B(n147), .C(SHA256_result[120]), .Y(f4_E_32[13])
         );
  XOR3X2 U2084 ( .A(n74), .B(n149), .C(SHA256_result[124]), .Y(f4_E_32[22]) );
  XOR3X2 U2085 ( .A(n153), .B(n146), .C(SHA256_result[122]), .Y(f4_E_32[15])
         );
  MX2X1 U2086 ( .A(SHA256_result[44]), .B(SHA256_result[76]), .S0(n150), .Y(
        f1_EFG_32[12]) );
  MX2X1 U2087 ( .A(SHA256_result[47]), .B(SHA256_result[79]), .S0(n149), .Y(
        f1_EFG_32[15]) );
  XOR3X2 U2088 ( .A(n151), .B(SHA256_result[101]), .C(SHA256_result[120]), .Y(
        f4_E_32[31]) );
  OAI21XL U2089 ( .A0(n189), .A1(n811), .B0(n1730), .Y(n2897) );
  AOI22X1 U2090 ( .A0(N939), .A1(n237), .B0(SHA256_result[216]), .B1(n10), .Y(
        n1730) );
  OAI21XL U2091 ( .A0(n189), .A1(n803), .B0(n1738), .Y(n2905) );
  OAI21XL U2092 ( .A0(n189), .A1(n797), .B0(n1744), .Y(n2911) );
  OAI21XL U2093 ( .A0(n186), .A1(n894), .B0(n1514), .Y(n2624) );
  OAI21XL U2094 ( .A0(n187), .A1(n906), .B0(n1502), .Y(n2612) );
  OAI21XL U2095 ( .A0(n187), .A1(n905), .B0(n1503), .Y(n2613) );
  AOI22X1 U2096 ( .A0(N1064), .A1(n240), .B0(SHA256_result[85]), .B1(n11), .Y(
        n1503) );
  OAI21XL U2097 ( .A0(n186), .A1(n885), .B0(n1615), .Y(n2799) );
  AOI22X1 U2098 ( .A0(N1037), .A1(n247), .B0(SHA256_result[122]), .B1(n10), 
        .Y(n1615) );
  OAI21XL U2099 ( .A0(n188), .A1(n882), .B0(n1618), .Y(n2802) );
  OAI21XL U2100 ( .A0(n189), .A1(n847), .B0(n1695), .Y(n2862) );
  AOI22X1 U2101 ( .A0(N974), .A1(n237), .B0(SHA256_result[187]), .B1(n11), .Y(
        n1695) );
  OAI21XL U2102 ( .A0(n189), .A1(n812), .B0(n1729), .Y(n2896) );
  AOI22X1 U2103 ( .A0(N940), .A1(n238), .B0(SHA256_result[217]), .B1(n11), .Y(
        n1729) );
  OAI21XL U2104 ( .A0(n189), .A1(n798), .B0(n1743), .Y(n2910) );
  OAI21XL U2105 ( .A0(n189), .A1(n810), .B0(n1731), .Y(n2898) );
  OAI21XL U2106 ( .A0(n189), .A1(n807), .B0(n1734), .Y(n2901) );
  AOI22X1 U2107 ( .A0(N935), .A1(n237), .B0(SHA256_result[212]), .B1(n11), .Y(
        n1734) );
  OAI21XL U2108 ( .A0(n189), .A1(n794), .B0(n1747), .Y(n2914) );
  OAI21XL U2109 ( .A0(n186), .A1(n903), .B0(n1505), .Y(n2615) );
  AOI22X1 U2110 ( .A0(N1062), .A1(n245), .B0(SHA256_result[83]), .B1(n11), .Y(
        n1505) );
  OAI21XL U2111 ( .A0(n186), .A1(n902), .B0(n1506), .Y(n2616) );
  OAI21XL U2112 ( .A0(n186), .A1(n893), .B0(n1515), .Y(n2625) );
  OAI21XL U2113 ( .A0(n188), .A1(n840), .B0(n1702), .Y(n2869) );
  AOI22X1 U2114 ( .A0(N967), .A1(n237), .B0(SHA256_result[180]), .B1(n11), .Y(
        n1702) );
  OAI21XL U2115 ( .A0(n187), .A1(n904), .B0(n1504), .Y(n2614) );
  AOI22X1 U2116 ( .A0(N1063), .A1(n239), .B0(SHA256_result[84]), .B1(n10), .Y(
        n1504) );
  OAI21XL U2117 ( .A0(n186), .A1(n897), .B0(n1511), .Y(n2621) );
  OAI21XL U2118 ( .A0(n186), .A1(n890), .B0(n1518), .Y(n2628) );
  OAI21XL U2119 ( .A0(n188), .A1(n881), .B0(n1619), .Y(n2803) );
  OAI21XL U2121 ( .A0(n188), .A1(n841), .B0(n1701), .Y(n2868) );
  AOI22X1 U2122 ( .A0(N968), .A1(n237), .B0(SHA256_result[181]), .B1(n10), .Y(
        n1701) );
  OAI21XL U2123 ( .A0(n705), .A1(n936), .B0(n1470), .Y(n2583) );
  OAI21XL U2124 ( .A0(n705), .A1(n935), .B0(n1471), .Y(n2584) );
  OAI21XL U2125 ( .A0(n705), .A1(n934), .B0(n1472), .Y(n2585) );
  OAI21XL U2126 ( .A0(n705), .A1(n933), .B0(n1473), .Y(n2586) );
  OAI21XL U2127 ( .A0(n705), .A1(n926), .B0(n1480), .Y(n2593) );
  OAI21XL U2128 ( .A0(n705), .A1(n919), .B0(n1487), .Y(n2600) );
  OAI21XL U2129 ( .A0(n705), .A1(n918), .B0(n1488), .Y(n2601) );
  OAI21XL U2130 ( .A0(n190), .A1(n822), .B0(n1720), .Y(n2887) );
  AOI22XL U2131 ( .A0(N949), .A1(n238), .B0(SHA256_result[162]), .B1(n10), .Y(
        n1720) );
  OAI21XL U2132 ( .A0(n190), .A1(n820), .B0(n1722), .Y(n2889) );
  OAI21XL U2133 ( .A0(n705), .A1(n930), .B0(n1476), .Y(n2589) );
  OAI21XL U2134 ( .A0(n705), .A1(n929), .B0(n1477), .Y(n2590) );
  OAI21XL U2135 ( .A0(n705), .A1(n924), .B0(n1482), .Y(n2595) );
  OAI21XL U2136 ( .A0(n705), .A1(n923), .B0(n1483), .Y(n2596) );
  OAI21XL U2137 ( .A0(n705), .A1(n922), .B0(n1484), .Y(n2597) );
  OAI21XL U2138 ( .A0(n188), .A1(n843), .B0(n1699), .Y(n2866) );
  AOI22X1 U2139 ( .A0(N970), .A1(n237), .B0(SHA256_result[183]), .B1(n10), .Y(
        n1699) );
  OAI21XL U2140 ( .A0(n188), .A1(n827), .B0(n1715), .Y(n2882) );
  OAI21XL U2141 ( .A0(n188), .A1(n826), .B0(n1716), .Y(n2883) );
  OAI21XL U2142 ( .A0(n188), .A1(n845), .B0(n1697), .Y(n2864) );
  AOI22X1 U2143 ( .A0(N972), .A1(n237), .B0(SHA256_result[185]), .B1(n11), .Y(
        n1697) );
  OAI21XL U2144 ( .A0(n188), .A1(n831), .B0(n1711), .Y(n2878) );
  OAI21XL U2145 ( .A0(n188), .A1(n829), .B0(n1713), .Y(n2880) );
  OAI2BB1X1 U2146 ( .A0N(N990), .A1N(n235), .B0(n463), .Y(n2846) );
  AOI2BB2X1 U2147 ( .B0(SHA256_result[107]), .B1(n195), .A0N(n12), .A1N(n462), 
        .Y(n463) );
  INVXL U2148 ( .A(next_E[11]), .Y(n462) );
  OAI2BB1X1 U2149 ( .A0N(N992), .A1N(n248), .B0(n457), .Y(n2844) );
  INVXL U2150 ( .A(next_E[13]), .Y(n456) );
  NAND2BX1 U2151 ( .AN(n542), .B(n541), .Y(n2954) );
  OAI21XL U2152 ( .A0(n760), .A1(n234), .B0(n636), .Y(n542) );
  OAI2BB1X1 U2153 ( .A0N(SHA256_result[209]), .A1N(n166), .B0(n557), .Y(
        f2_ABC_32[17]) );
  OAI21XL U2154 ( .A0(SHA256_result[209]), .A1(n166), .B0(SHA256_result[177]), 
        .Y(n557) );
  OAI2BB1X1 U2155 ( .A0N(SHA256_result[206]), .A1N(n169), .B0(n560), .Y(
        f2_ABC_32[14]) );
  OAI21XL U2156 ( .A0(SHA256_result[206]), .A1(n169), .B0(SHA256_result[174]), 
        .Y(n560) );
  OAI2BB1X1 U2157 ( .A0N(SHA256_result[207]), .A1N(n168), .B0(n559), .Y(
        f2_ABC_32[15]) );
  OAI21XL U2158 ( .A0(SHA256_result[207]), .A1(n168), .B0(SHA256_result[175]), 
        .Y(n559) );
  OAI2BB1X1 U2159 ( .A0N(SHA256_result[204]), .A1N(n171), .B0(n562), .Y(
        f2_ABC_32[12]) );
  OAI21XL U2160 ( .A0(SHA256_result[204]), .A1(n171), .B0(SHA256_result[172]), 
        .Y(n562) );
  OAI2BB1X1 U2161 ( .A0N(SHA256_result[205]), .A1N(n170), .B0(n561), .Y(
        f2_ABC_32[13]) );
  OAI21XL U2162 ( .A0(SHA256_result[205]), .A1(n170), .B0(SHA256_result[173]), 
        .Y(n561) );
  XOR3X2 U2163 ( .A(SHA256_result[98]), .B(SHA256_result[112]), .C(
        SHA256_result[125]), .Y(f4_E_32[23]) );
  XOR3X2 U2164 ( .A(SHA256_result[127]), .B(SHA256_result[109]), .C(
        SHA256_result[122]), .Y(f4_E_32[20]) );
  MX2X1 U2165 ( .A(SHA256_result[56]), .B(SHA256_result[88]), .S0(
        SHA256_result[120]), .Y(f1_EFG_32[24]) );
  MX2X1 U2166 ( .A(SHA256_result[55]), .B(SHA256_result[87]), .S0(
        SHA256_result[119]), .Y(f1_EFG_32[23]) );
  MX2X1 U2167 ( .A(SHA256_result[54]), .B(SHA256_result[86]), .S0(
        SHA256_result[118]), .Y(f1_EFG_32[22]) );
  XOR3X2 U2168 ( .A(n178), .B(n166), .C(SHA256_result[252]), .Y(f3_A_32[15])
         );
  XOR3X2 U2169 ( .A(n163), .B(n175), .C(SHA256_result[255]), .Y(f3_A_32[18])
         );
  XOR3X2 U2170 ( .A(SHA256_result[99]), .B(n148), .C(n145), .Y(f4_E_32[24]) );
  MX2X1 U2171 ( .A(SHA256_result[52]), .B(SHA256_result[84]), .S0(
        SHA256_result[116]), .Y(f1_EFG_32[20]) );
  AOI31X1 U2172 ( .A0(n2522), .A1(n2523), .A2(n2524), .B0(n268), .Y(N3004) );
  AND3X2 U2173 ( .A(n2288), .B(n2256), .C(n746), .Y(n2523) );
  AOI211X1 U2174 ( .A0(n2371), .A1(n1389), .B0(n2525), .C0(n2239), .Y(n2524)
         );
  AOI31X1 U2175 ( .A0(n2488), .A1(n2489), .A2(n2490), .B0(n268), .Y(N3009) );
  NOR3X1 U2176 ( .A(n2347), .B(n2372), .C(n2314), .Y(n2489) );
  AOI211X1 U2177 ( .A0(n2391), .A1(n1389), .B0(n2491), .C0(n2492), .Y(n2490)
         );
  AOI31X1 U2178 ( .A0(n2401), .A1(n2402), .A2(n2403), .B0(n269), .Y(N3019) );
  AOI211X1 U2179 ( .A0(n2343), .A1(n1371), .B0(n2404), .C0(n2405), .Y(n2403)
         );
  AOI31X1 U2180 ( .A0(n2264), .A1(n2265), .A2(n2266), .B0(n269), .Y(N3031) );
  AOI31X1 U2181 ( .A0(n738), .A1(n1384), .A2(n2258), .B0(n2275), .Y(n2264) );
  NOR3BX1 U2182 ( .AN(n2272), .B(n2273), .C(n2274), .Y(n2265) );
  AOI211X1 U2183 ( .A0(n2267), .A1(n129), .B0(n2268), .C0(n728), .Y(n2266) );
  AOI31X1 U2184 ( .A0(n2459), .A1(n2460), .A2(n2461), .B0(n268), .Y(N3013) );
  AOI2BB2X1 U2185 ( .B0(n2260), .B1(n328), .A0N(n2269), .A1N(n730), .Y(n2459)
         );
  AOI22X1 U2186 ( .A0(n2381), .A1(n1384), .B0(n2312), .B1(n335), .Y(n2460) );
  AOI31X1 U2187 ( .A0(n2315), .A1(n2316), .A2(n2317), .B0(n269), .Y(N3027) );
  AOI2BB2X1 U2188 ( .B0(n2299), .B1(n130), .A0N(n2307), .A1N(n333), .Y(n2315)
         );
  AOI22X1 U2189 ( .A0(n2324), .A1(n1384), .B0(n2325), .B1(n2261), .Y(n2316) );
  AOI211X1 U2190 ( .A0(n2318), .A1(n1397), .B0(n2319), .C0(n2320), .Y(n2317)
         );
  AOI31X1 U2191 ( .A0(n2514), .A1(n2515), .A2(n2516), .B0(n268), .Y(N3005) );
  AOI32X1 U2192 ( .A0(n328), .A1(n1389), .A2(n2428), .B0(n129), .B1(n2521), 
        .Y(n2514) );
  AOI211X1 U2193 ( .A0(n2445), .A1(n336), .B0(n2517), .C0(n2509), .Y(n2516) );
  AOI31X1 U2194 ( .A0(n2301), .A1(n2302), .A2(n2303), .B0(n269), .Y(N3028) );
  NOR3BX1 U2195 ( .AN(n2304), .B(n2305), .C(n2306), .Y(n2303) );
  AOI21X1 U2196 ( .A0(n2310), .A1(n182), .B0(n728), .Y(n2301) );
  AOI31X1 U2197 ( .A0(n2480), .A1(n2481), .A2(n2482), .B0(n268), .Y(N3010) );
  AOI222X1 U2198 ( .A0(n2486), .A1(n2406), .B0(n2487), .B1(n1389), .C0(n2409), 
        .C1(n47), .Y(n2481) );
  NOR4BX1 U2199 ( .AN(n733), .B(n2483), .C(n2484), .D(n2485), .Y(n2482) );
  AOI31X1 U2200 ( .A0(n2290), .A1(n2291), .A2(n2292), .B0(n269), .Y(N3029) );
  AOI222X1 U2201 ( .A0(n2298), .A1(n1384), .B0(n2247), .B1(n1371), .C0(n2299), 
        .C1(n336), .Y(n2291) );
  NOR3X1 U2202 ( .A(n2293), .B(n2294), .C(n2295), .Y(n2292) );
  AOI31X1 U2203 ( .A0(n2350), .A1(n2351), .A2(n2352), .B0(n269), .Y(N3024) );
  AOI22X1 U2204 ( .A0(n2361), .A1(n1371), .B0(n2261), .B1(n2259), .Y(n2350) );
  NOR3X1 U2205 ( .A(n2353), .B(n2354), .C(n2294), .Y(n2352) );
  AOI211X1 U2206 ( .A0(n2262), .A1(n2358), .B0(n2359), .C0(n2360), .Y(n2351)
         );
  AOI31X1 U2207 ( .A0(n2376), .A1(n2377), .A2(n2378), .B0(n269), .Y(N3022) );
  AOI222X1 U2208 ( .A0(n2259), .A1(n717), .B0(n2355), .B1(n726), .C0(n2381), 
        .C1(n1384), .Y(n2377) );
  AND4X2 U2209 ( .A(n2379), .B(n750), .C(n2282), .D(n739), .Y(n2378) );
  OAI2BB1X1 U2210 ( .A0N(SHA256_result[214]), .A1N(n37), .B0(n552), .Y(
        f2_ABC_32[22]) );
  OAI21XL U2211 ( .A0(SHA256_result[214]), .A1(n37), .B0(SHA256_result[182]), 
        .Y(n552) );
  OAI2BB1X1 U2212 ( .A0N(SHA256_result[212]), .A1N(n163), .B0(n554), .Y(
        f2_ABC_32[20]) );
  OAI21XL U2213 ( .A0(SHA256_result[212]), .A1(n163), .B0(SHA256_result[180]), 
        .Y(n554) );
  OAI2BB1X1 U2214 ( .A0N(SHA256_result[213]), .A1N(n162), .B0(n553), .Y(
        f2_ABC_32[21]) );
  OAI21XL U2215 ( .A0(SHA256_result[213]), .A1(n162), .B0(SHA256_result[181]), 
        .Y(n553) );
  OAI2BB1X1 U2216 ( .A0N(SHA256_result[211]), .A1N(n164), .B0(n555), .Y(
        f2_ABC_32[19]) );
  OAI21XL U2217 ( .A0(SHA256_result[211]), .A1(n164), .B0(SHA256_result[179]), 
        .Y(n555) );
  OAI2BB1X1 U2218 ( .A0N(SHA256_result[208]), .A1N(n167), .B0(n558), .Y(
        f2_ABC_32[16]) );
  OAI21XL U2219 ( .A0(SHA256_result[208]), .A1(n167), .B0(SHA256_result[176]), 
        .Y(n558) );
  OAI2BB1X1 U2220 ( .A0N(SHA256_result[210]), .A1N(n165), .B0(n556), .Y(
        f2_ABC_32[18]) );
  OAI21XL U2221 ( .A0(SHA256_result[210]), .A1(n165), .B0(SHA256_result[178]), 
        .Y(n556) );
  XOR3X2 U2222 ( .A(SHA256_result[127]), .B(SHA256_result[100]), .C(
        SHA256_result[114]), .Y(f4_E_32[25]) );
  XOR3X2 U2223 ( .A(n77), .B(SHA256_result[101]), .C(n147), .Y(f4_E_32[26]) );
  XOR3X2 U2224 ( .A(n154), .B(n74), .C(SHA256_result[116]), .Y(f4_E_32[27]) );
  XOR3X2 U2225 ( .A(SHA256_result[98]), .B(SHA256_result[103]), .C(n146), .Y(
        f4_E_32[28]) );
  MX2X1 U2226 ( .A(SHA256_result[58]), .B(SHA256_result[90]), .S0(
        SHA256_result[122]), .Y(f1_EFG_32[26]) );
  MX2X1 U2227 ( .A(SHA256_result[60]), .B(SHA256_result[92]), .S0(
        SHA256_result[124]), .Y(f1_EFG_32[28]) );
  XOR3X2 U2228 ( .A(n72), .B(n173), .C(n37), .Y(f3_A_32[20]) );
  MX2X1 U2229 ( .A(SHA256_result[59]), .B(SHA256_result[91]), .S0(n73), .Y(
        f1_EFG_32[27]) );
  MX2X1 U2230 ( .A(SHA256_result[57]), .B(SHA256_result[89]), .S0(
        SHA256_result[121]), .Y(f1_EFG_32[25]) );
  NAND2X1 U2231 ( .A(n142), .B(n1976), .Y(N3453) );
  XNOR2X1 U2232 ( .A(read_counter[5]), .B(n704), .Y(n142) );
  NAND2X1 U2233 ( .A(n143), .B(n1976), .Y(N3452) );
  XOR2X1 U2234 ( .A(read_counter[4]), .B(n703), .Y(n143) );
  NAND2BX1 U2235 ( .AN(N3435), .B(n1976), .Y(N3451) );
  NAND2BX1 U2236 ( .AN(N3434), .B(n1976), .Y(N3450) );
  NAND2BX1 U2237 ( .AN(N3433), .B(n1976), .Y(N3449) );
  NAND2X1 U2238 ( .A(read_counter[0]), .B(n1976), .Y(N3448) );
  OAI2BB1X1 U2239 ( .A0N(SHA256_result[217]), .A1N(n159), .B0(n549), .Y(
        f2_ABC_32[25]) );
  OAI21XL U2240 ( .A0(SHA256_result[217]), .A1(n159), .B0(SHA256_result[185]), 
        .Y(n549) );
  OAI2BB1X1 U2241 ( .A0N(SHA256_result[215]), .A1N(n161), .B0(n551), .Y(
        f2_ABC_32[23]) );
  OAI21XL U2242 ( .A0(SHA256_result[215]), .A1(n161), .B0(SHA256_result[183]), 
        .Y(n551) );
  OAI2BB1X1 U2243 ( .A0N(SHA256_result[216]), .A1N(n160), .B0(n550), .Y(
        f2_ABC_32[24]) );
  OAI21XL U2244 ( .A0(SHA256_result[216]), .A1(n160), .B0(SHA256_result[184]), 
        .Y(n550) );
  OAI2BB1X1 U2245 ( .A0N(SHA256_result[218]), .A1N(n158), .B0(n548), .Y(
        f2_ABC_32[26]) );
  OAI21XL U2246 ( .A0(SHA256_result[218]), .A1(n158), .B0(SHA256_result[186]), 
        .Y(n548) );
  XOR3X2 U2247 ( .A(n152), .B(SHA256_result[100]), .C(SHA256_result[119]), .Y(
        f4_E_32[30]) );
  XOR3X2 U2248 ( .A(n153), .B(SHA256_result[99]), .C(SHA256_result[118]), .Y(
        f4_E_32[29]) );
  MX2X1 U2249 ( .A(SHA256_result[61]), .B(SHA256_result[93]), .S0(
        SHA256_result[125]), .Y(f1_EFG_32[29]) );
  XOR3X2 U2250 ( .A(n167), .B(n176), .C(SHA256_result[252]), .Y(f3_A_32[26])
         );
  MX2X1 U2251 ( .A(SHA256_result[62]), .B(SHA256_result[94]), .S0(n145), .Y(
        f1_EFG_32[30]) );
  NOR2X1 U2252 ( .A(n729), .B(n1371), .Y(n2314) );
  AOI211X1 U2253 ( .A0(n708), .A1(n1384), .B0(n2382), .C0(n2370), .Y(n2518) );
  OAI2BB1X1 U2254 ( .A0N(SHA256_result[220]), .A1N(SHA256_result[252]), .B0(
        n546), .Y(f2_ABC_32[28]) );
  OAI21XL U2255 ( .A0(SHA256_result[220]), .A1(SHA256_result[252]), .B0(
        SHA256_result[188]), .Y(n546) );
  OAI2BB1X1 U2256 ( .A0N(SHA256_result[219]), .A1N(n157), .B0(n547), .Y(
        f2_ABC_32[27]) );
  OAI21XL U2257 ( .A0(SHA256_result[219]), .A1(n157), .B0(SHA256_result[187]), 
        .Y(n547) );
  OAI2BB1X1 U2258 ( .A0N(SHA256_result[222]), .A1N(n155), .B0(n544), .Y(
        f2_ABC_32[30]) );
  OAI21XL U2259 ( .A0(SHA256_result[222]), .A1(n155), .B0(SHA256_result[190]), 
        .Y(n544) );
  OAI2BB1X1 U2260 ( .A0N(SHA256_result[221]), .A1N(n156), .B0(n545), .Y(
        f2_ABC_32[29]) );
  OAI21XL U2261 ( .A0(SHA256_result[221]), .A1(n156), .B0(SHA256_result[189]), 
        .Y(n545) );
  INVX1 U2262 ( .A(n2311), .Y(n728) );
  AOI221X1 U2263 ( .A0(n330), .A1(n2312), .B0(n1389), .B1(n2313), .C0(n2314), 
        .Y(n2311) );
  XOR3X2 U2264 ( .A(n164), .B(n173), .C(SHA256_result[255]), .Y(f3_A_32[29])
         );
  INVX1 U2265 ( .A(n1397), .Y(n329) );
  MX2X1 U2266 ( .A(SHA256_result[63]), .B(SHA256_result[95]), .S0(
        SHA256_result[127]), .Y(f1_EFG_32[31]) );
  NOR2X1 U2267 ( .A(n742), .B(n1389), .Y(n2259) );
  NOR2X1 U2268 ( .A(n749), .B(n1389), .Y(n2267) );
  OAI222XL U2269 ( .A0(n718), .A1(n1389), .B0(n2369), .B1(n183), .C0(n735), 
        .C1(n336), .Y(n2368) );
  AOI211X1 U2270 ( .A0(n1384), .A1(n2261), .B0(n2342), .C0(n2370), .Y(n2369)
         );
  OAI222XL U2271 ( .A0(n758), .A1(n140), .B0(n336), .B1(n734), .C0(n1389), 
        .C1(n716), .Y(n2404) );
  OAI221XL U2272 ( .A0(n755), .A1(n330), .B0(n1389), .B1(n717), .C0(n2307), 
        .Y(n2442) );
  NOR2X1 U2273 ( .A(n726), .B(n1389), .Y(n2438) );
  OR2X2 U2274 ( .A(read_counter[1]), .B(read_counter[0]), .Y(n701) );
  NOR2X1 U2275 ( .A(n1384), .B(n335), .Y(n2244) );
  NOR2X1 U2276 ( .A(n738), .B(n1389), .Y(n2325) );
  OAI31X1 U2277 ( .A0(n730), .A1(n752), .A2(n1384), .B0(n2333), .Y(n2407) );
  NOR2X1 U2278 ( .A(n749), .B(n1384), .Y(n2251) );
  NOR2X1 U2279 ( .A(n1384), .B(n332), .Y(n2447) );
  NAND2X1 U2280 ( .A(n743), .B(n1389), .Y(n2256) );
  NAND2X1 U2281 ( .A(n131), .B(n1384), .Y(n2296) );
  NOR2X1 U2282 ( .A(n725), .B(n1384), .Y(n2247) );
  NOR2X1 U2283 ( .A(n2289), .B(n1389), .Y(n2321) );
  NOR2X1 U2284 ( .A(n738), .B(n1384), .Y(n2410) );
  NOR2X1 U2285 ( .A(n140), .B(n1389), .Y(n2308) );
  NAND2X1 U2286 ( .A(n40), .B(n1389), .Y(n2397) );
  NOR2X1 U2287 ( .A(n757), .B(n1371), .Y(n2390) );
  NOR2X1 U2288 ( .A(n726), .B(n1384), .Y(n2425) );
  AOI31X1 U2289 ( .A0(n1389), .A1(n1371), .A2(n2261), .B0(n2354), .Y(n2433) );
  AOI21X1 U2290 ( .A0(n2288), .A1(n719), .B0(n1389), .Y(n2287) );
  AOI21X1 U2291 ( .A0(n714), .A1(n2304), .B0(n1389), .Y(n2418) );
  NAND4X1 U2292 ( .A(n2211), .B(n2212), .C(n2213), .D(n2214), .Y(n2210) );
  NAND4X1 U2293 ( .A(n2173), .B(n2174), .C(n2175), .D(n2176), .Y(n2172) );
  NAND4X1 U2294 ( .A(n2131), .B(n2132), .C(n2133), .D(n2134), .Y(n2130) );
  NAND4X1 U2295 ( .A(n2109), .B(n2110), .C(n2111), .D(n2112), .Y(n2108) );
  NAND4X1 U2296 ( .A(n2089), .B(n2090), .C(n2091), .D(n2092), .Y(n2088) );
  NAND4X1 U2297 ( .A(n2035), .B(n2036), .C(n2037), .D(n2038), .Y(n2034) );
  NAND4X1 U2298 ( .A(n1984), .B(n1985), .C(n1986), .D(n1987), .Y(n1983) );
  NAND4X1 U2299 ( .A(n2225), .B(n2226), .C(n2227), .D(n2228), .Y(n2208) );
  AOI22X1 U2300 ( .A0(n2069), .A1(SHA256_result[184]), .B0(n2070), .B1(
        SHA256_result[188]), .Y(n2225) );
  NAND4X1 U2301 ( .A(n2193), .B(n2194), .C(n2195), .D(n2196), .Y(n2170) );
  AOI22X1 U2302 ( .A0(n2018), .A1(SHA256_result[56]), .B0(n2019), .B1(
        SHA256_result[60]), .Y(n2193) );
  NAND4X1 U2303 ( .A(n2159), .B(n2160), .C(n2161), .D(n2162), .Y(n2148) );
  AOI22X1 U2304 ( .A0(n2069), .A1(SHA256_result[185]), .B0(n2070), .B1(
        SHA256_result[189]), .Y(n2159) );
  NAND4X1 U2305 ( .A(n2139), .B(n2140), .C(n2141), .D(n2142), .Y(n2128) );
  AOI22X1 U2306 ( .A0(n2018), .A1(SHA256_result[57]), .B0(n2019), .B1(
        SHA256_result[61]), .Y(n2139) );
  NAND4X1 U2307 ( .A(n2117), .B(n2118), .C(n2119), .D(n2120), .Y(n2106) );
  AOI22X1 U2308 ( .A0(n2069), .A1(SHA256_result[186]), .B0(n2070), .B1(
        SHA256_result[190]), .Y(n2117) );
  NAND4X1 U2309 ( .A(n2097), .B(n2098), .C(n2099), .D(n2100), .Y(n2086) );
  AOI22X1 U2310 ( .A0(n2018), .A1(SHA256_result[58]), .B0(n2019), .B1(
        SHA256_result[62]), .Y(n2097) );
  NAND4X1 U2311 ( .A(n2059), .B(n2060), .C(n2061), .D(n2062), .Y(n2032) );
  AOI22X1 U2312 ( .A0(n2069), .A1(SHA256_result[187]), .B0(n2070), .B1(
        SHA256_result[191]), .Y(n2059) );
  NAND4X1 U2313 ( .A(n2008), .B(n2009), .C(n2010), .D(n2011), .Y(n1981) );
  AOI22X1 U2314 ( .A0(n2018), .A1(SHA256_result[59]), .B0(n2019), .B1(
        SHA256_result[63]), .Y(n2008) );
  NAND4X1 U2315 ( .A(n2219), .B(n2220), .C(n2221), .D(n2222), .Y(n2209) );
  AOI22X1 U2316 ( .A0(n2057), .A1(SHA256_result[216]), .B0(n2058), .B1(
        SHA256_result[220]), .Y(n2219) );
  NAND4X1 U2317 ( .A(n2183), .B(n2184), .C(n2185), .D(n2186), .Y(n2171) );
  AOI22X1 U2318 ( .A0(n2006), .A1(SHA256_result[88]), .B0(n2007), .B1(
        SHA256_result[92]), .Y(n2183) );
  NAND4X1 U2319 ( .A(n2155), .B(n2156), .C(n2157), .D(n2158), .Y(n2149) );
  AOI22X1 U2320 ( .A0(n2057), .A1(SHA256_result[217]), .B0(n2058), .B1(
        SHA256_result[221]), .Y(n2155) );
  NAND4X1 U2321 ( .A(n2135), .B(n2136), .C(n2137), .D(n2138), .Y(n2129) );
  AOI22X1 U2322 ( .A0(n2006), .A1(SHA256_result[89]), .B0(n2007), .B1(
        SHA256_result[93]), .Y(n2135) );
  NAND4X1 U2323 ( .A(n2113), .B(n2114), .C(n2115), .D(n2116), .Y(n2107) );
  AOI22X1 U2324 ( .A0(n2057), .A1(SHA256_result[218]), .B0(n2058), .B1(
        SHA256_result[222]), .Y(n2113) );
  NAND4X1 U2325 ( .A(n2093), .B(n2094), .C(n2095), .D(n2096), .Y(n2087) );
  AOI22X1 U2326 ( .A0(n2006), .A1(SHA256_result[90]), .B0(n2007), .B1(
        SHA256_result[94]), .Y(n2093) );
  NAND4X1 U2327 ( .A(n2047), .B(n2048), .C(n2049), .D(n2050), .Y(n2033) );
  AOI22X1 U2328 ( .A0(n2057), .A1(SHA256_result[219]), .B0(n2058), .B1(
        SHA256_result[223]), .Y(n2047) );
  NAND4X1 U2329 ( .A(n1996), .B(n1997), .C(n1998), .D(n1999), .Y(n1982) );
  AOI22X1 U2330 ( .A0(n2006), .A1(SHA256_result[91]), .B0(n2007), .B1(
        SHA256_result[95]), .Y(n1996) );
  NAND4X1 U2331 ( .A(n2233), .B(n2234), .C(n2235), .D(n2236), .Y(n2207) );
  AOI22X1 U2332 ( .A0(n2081), .A1(SHA256_result[152]), .B0(n2082), .B1(
        SHA256_result[156]), .Y(n2233) );
  AOI22X1 U2333 ( .A0(n2079), .A1(SHA256_result[144]), .B0(n2080), .B1(
        SHA256_result[148]), .Y(n2234) );
  AOI22X1 U2334 ( .A0(n2077), .A1(SHA256_result[136]), .B0(n2078), .B1(
        SHA256_result[140]), .Y(n2235) );
  NAND4X1 U2335 ( .A(n2163), .B(n2164), .C(n2165), .D(n2166), .Y(n2147) );
  AOI22X1 U2336 ( .A0(n2081), .A1(SHA256_result[153]), .B0(n2082), .B1(
        SHA256_result[157]), .Y(n2163) );
  AOI22X1 U2337 ( .A0(n2079), .A1(SHA256_result[145]), .B0(n2080), .B1(
        SHA256_result[149]), .Y(n2164) );
  AOI22X1 U2338 ( .A0(n2077), .A1(SHA256_result[137]), .B0(n2078), .B1(
        SHA256_result[141]), .Y(n2165) );
  NAND4X1 U2339 ( .A(n2121), .B(n2122), .C(n2123), .D(n2124), .Y(n2105) );
  AOI22X1 U2340 ( .A0(n2081), .A1(SHA256_result[154]), .B0(n2082), .B1(
        SHA256_result[158]), .Y(n2121) );
  AOI22X1 U2341 ( .A0(n2079), .A1(SHA256_result[146]), .B0(n2080), .B1(
        SHA256_result[150]), .Y(n2122) );
  AOI22X1 U2342 ( .A0(n2077), .A1(SHA256_result[138]), .B0(n2078), .B1(
        SHA256_result[142]), .Y(n2123) );
  NAND4X1 U2343 ( .A(n2071), .B(n2072), .C(n2073), .D(n2074), .Y(n2031) );
  AOI22X1 U2344 ( .A0(n2081), .A1(SHA256_result[155]), .B0(n2082), .B1(
        SHA256_result[159]), .Y(n2071) );
  AOI22X1 U2345 ( .A0(n2079), .A1(SHA256_result[147]), .B0(n2080), .B1(
        SHA256_result[151]), .Y(n2072) );
  AOI22X1 U2346 ( .A0(n2077), .A1(SHA256_result[139]), .B0(n2078), .B1(
        SHA256_result[143]), .Y(n2073) );
  NOR2X1 U2347 ( .A(read_counter[5]), .B(read_counter[0]), .Y(n2191) );
  NOR2X1 U2348 ( .A(read_counter[4]), .B(read_counter[1]), .Y(n2205) );
  NOR2X1 U2349 ( .A(n950), .B(read_counter[0]), .Y(n2224) );
  NOR2X1 U2350 ( .A(n948), .B(read_counter[4]), .Y(n2206) );
  AOI22XL U2351 ( .A0(n1988), .A1(n74), .B0(n1989), .B1(SHA256_result[101]), 
        .Y(n2134) );
  AOI22XL U2352 ( .A0(n1988), .A1(SHA256_result[99]), .B0(n1989), .B1(
        SHA256_result[103]), .Y(n1987) );
  AOI22XL U2353 ( .A0(n1988), .A1(SHA256_result[98]), .B0(n1989), .B1(n154), 
        .Y(n2092) );
  AOI22X1 U2354 ( .A0(n2029), .A1(SHA256_result[24]), .B0(n2030), .B1(
        SHA256_result[28]), .Y(n2201) );
  AOI22X1 U2355 ( .A0(n2029), .A1(SHA256_result[25]), .B0(n2030), .B1(
        SHA256_result[29]), .Y(n2143) );
  AOI22X1 U2356 ( .A0(n2029), .A1(SHA256_result[26]), .B0(n2030), .B1(
        SHA256_result[30]), .Y(n2101) );
  AOI22X1 U2357 ( .A0(n2029), .A1(SHA256_result[27]), .B0(n2030), .B1(
        SHA256_result[31]), .Y(n2020) );
  OAI21XL U2358 ( .A0(round[3]), .A1(n2493), .B0(n2494), .Y(n2492) );
  AOI22X1 U2359 ( .A0(n726), .A1(n1371), .B0(n2258), .B1(n182), .Y(n2493) );
  OAI21XL U2360 ( .A0(n2306), .A1(n2449), .B0(n332), .Y(n2494) );
  BUFX3 U2361 ( .A(n334), .Y(n182) );
  OAI2BB1X1 U2362 ( .A0N(SHA256_result[223]), .A1N(SHA256_result[255]), .B0(
        n543), .Y(f2_ABC_32[31]) );
  OAI21XL U2363 ( .A0(SHA256_result[223]), .A1(SHA256_result[255]), .B0(
        SHA256_result[191]), .Y(n543) );
  INVX1 U2364 ( .A(read_counter[2]), .Y(n949) );
  INVX1 U2365 ( .A(read_counter[1]), .Y(n948) );
  INVX1 U2366 ( .A(read_counter[5]), .Y(n950) );
  NOR2X1 U2367 ( .A(n1389), .B(n332), .Y(n2486) );
  NOR3X1 U2368 ( .A(n717), .B(n1384), .C(n1371), .Y(n2360) );
  INVX1 U2369 ( .A(SHA256_result[218]), .Y(n786) );
  INVX1 U2370 ( .A(SHA256_result[184]), .Y(n811) );
  INVX1 U2371 ( .A(SHA256_result[90]), .Y(n885) );
  INVX1 U2372 ( .A(SHA256_result[214]), .Y(n782) );
  INVX1 U2373 ( .A(SHA256_result[219]), .Y(n787) );
  INVX1 U2374 ( .A(SHA256_result[222]), .Y(n790) );
  INVX1 U2375 ( .A(SHA256_result[215]), .Y(n783) );
  INVX1 U2376 ( .A(SHA256_result[212]), .Y(n780) );
  INVX1 U2377 ( .A(SHA256_result[221]), .Y(n789) );
  INVX1 U2378 ( .A(SHA256_result[220]), .Y(n788) );
  INVX1 U2379 ( .A(SHA256_result[213]), .Y(n781) );
  INVX1 U2380 ( .A(SHA256_result[155]), .Y(n847) );
  INVX1 U2381 ( .A(SHA256_result[156]), .Y(n848) );
  INVXL U2382 ( .A(SHA256_result[103]), .Y(n479) );
  INVX1 U2383 ( .A(SHA256_result[185]), .Y(n812) );
  INVX1 U2384 ( .A(SHA256_result[186]), .Y(n813) );
  INVX1 U2385 ( .A(SHA256_result[190]), .Y(n817) );
  INVX1 U2386 ( .A(SHA256_result[183]), .Y(n810) );
  INVX1 U2387 ( .A(SHA256_result[180]), .Y(n807) );
  INVX1 U2388 ( .A(SHA256_result[189]), .Y(n816) );
  INVX1 U2389 ( .A(SHA256_result[182]), .Y(n809) );
  INVX1 U2390 ( .A(SHA256_result[59]), .Y(n911) );
  INVX1 U2391 ( .A(SHA256_result[57]), .Y(n909) );
  INVX1 U2392 ( .A(SHA256_result[56]), .Y(n908) );
  INVX1 U2393 ( .A(SHA256_result[148]), .Y(n840) );
  INVX1 U2394 ( .A(SHA256_result[63]), .Y(n915) );
  INVX1 U2395 ( .A(SHA256_result[61]), .Y(n913) );
  INVX1 U2396 ( .A(SHA256_result[60]), .Y(n912) );
  INVX1 U2397 ( .A(SHA256_result[88]), .Y(n883) );
  INVX1 U2398 ( .A(SHA256_result[94]), .Y(n889) );
  INVX1 U2399 ( .A(SHA256_result[93]), .Y(n888) );
  INVX1 U2400 ( .A(SHA256_result[149]), .Y(n841) );
  INVX1 U2401 ( .A(SHA256_result[26]), .Y(n943) );
  INVX1 U2402 ( .A(SHA256_result[29]), .Y(n946) );
  INVX1 U2403 ( .A(SHA256_result[158]), .Y(n850) );
  INVX1 U2404 ( .A(SHA256_result[151]), .Y(n843) );
  INVX1 U2405 ( .A(SHA256_result[135]), .Y(n827) );
  INVX1 U2406 ( .A(SHA256_result[134]), .Y(n826) );
  INVX1 U2407 ( .A(SHA256_result[31]), .Y(n916) );
  INVX1 U2408 ( .A(SHA256_result[153]), .Y(n845) );
  INVX1 U2409 ( .A(SHA256_result[139]), .Y(n831) );
  INVX1 U2410 ( .A(SHA256_result[137]), .Y(n829) );
  INVX1 U2411 ( .A(SHA256_result[217]), .Y(n785) );
  INVX1 U2412 ( .A(SHA256_result[216]), .Y(n784) );
  INVXL U2413 ( .A(SHA256_result[99]), .Y(n495) );
  INVXL U2414 ( .A(n74), .Y(n502) );
  INVX1 U2415 ( .A(SHA256_result[154]), .Y(n846) );
  INVX1 U2416 ( .A(SHA256_result[223]), .Y(n759) );
  INVX1 U2417 ( .A(SHA256_result[187]), .Y(n814) );
  INVX1 U2418 ( .A(SHA256_result[188]), .Y(n815) );
  INVX1 U2419 ( .A(SHA256_result[181]), .Y(n808) );
  INVX1 U2420 ( .A(SHA256_result[143]), .Y(n835) );
  INVX1 U2421 ( .A(SHA256_result[91]), .Y(n886) );
  INVX1 U2422 ( .A(SHA256_result[89]), .Y(n884) );
  INVX1 U2423 ( .A(SHA256_result[58]), .Y(n910) );
  INVX1 U2424 ( .A(SHA256_result[92]), .Y(n887) );
  INVX1 U2425 ( .A(SHA256_result[152]), .Y(n844) );
  INVX1 U2426 ( .A(SHA256_result[27]), .Y(n944) );
  INVX1 U2427 ( .A(SHA256_result[25]), .Y(n942) );
  INVX1 U2428 ( .A(SHA256_result[24]), .Y(n941) );
  INVX1 U2429 ( .A(SHA256_result[145]), .Y(n837) );
  INVX1 U2430 ( .A(SHA256_result[144]), .Y(n836) );
  INVX1 U2431 ( .A(SHA256_result[138]), .Y(n830) );
  INVX1 U2432 ( .A(SHA256_result[136]), .Y(n828) );
  INVX1 U2433 ( .A(SHA256_result[28]), .Y(n945) );
  INVX1 U2434 ( .A(SHA256_result[157]), .Y(n849) );
  INVX1 U2435 ( .A(SHA256_result[150]), .Y(n842) );
  INVX1 U2436 ( .A(SHA256_result[142]), .Y(n834) );
  INVX1 U2437 ( .A(SHA256_result[140]), .Y(n832) );
  INVX1 U2438 ( .A(SHA256_result[133]), .Y(n825) );
  INVX1 U2439 ( .A(SHA256_result[132]), .Y(n824) );
  INVX1 U2440 ( .A(SHA256_result[159]), .Y(n819) );
  INVX1 U2441 ( .A(SHA256_result[147]), .Y(n839) );
  INVX1 U2442 ( .A(SHA256_result[146]), .Y(n838) );
  INVX1 U2443 ( .A(SHA256_result[141]), .Y(n833) );
  AOI21XL U2444 ( .A0(next_A[28]), .A1(n10), .B0(n583), .Y(n584) );
  AOI21XL U2445 ( .A0(next_E[25]), .A1(n10), .B0(n427), .Y(n428) );
  NAND2XL U2446 ( .A(next_E[28]), .B(n10), .Y(n415) );
  AOI21XL U2447 ( .A0(n52), .A1(n10), .B0(n432), .Y(n433) );
  AOI21XL U2448 ( .A0(next_E[29]), .A1(n11), .B0(n411), .Y(n412) );
  NAND2XL U2449 ( .A(next_A[29]), .B(n11), .Y(n581) );
  AOI21XL U2450 ( .A0(next_A[23]), .A1(n11), .B0(n602), .Y(n603) );
  AOI2BB2XL U2451 ( .B0(n193), .B1(n149), .A0N(n14), .A1N(n451), .Y(n452) );
  OAI2BB1X1 U2452 ( .A0N(N994), .A1N(n245), .B0(n452), .Y(n2842) );
  INVXL U2453 ( .A(next_A[13]), .Y(n630) );
  INVXL U2454 ( .A(next_E[15]), .Y(n451) );
  INVXL U2455 ( .A(next_A[15]), .Y(n624) );
  AOI21XL U2456 ( .A0(next_E[26]), .A1(n11), .B0(n423), .Y(n424) );
  NAND2XL U2457 ( .A(next_A[27]), .B(n11), .Y(n586) );
  AOI21XL U2458 ( .A0(next_A[26]), .A1(n11), .B0(n590), .Y(n591) );
  NAND2XL U2459 ( .A(next_A[25]), .B(n10), .Y(n594) );
  OAI2BB1X1 U2460 ( .A0N(read_counter[0]), .A1N(read_counter[1]), .B0(n701), 
        .Y(N3433) );
  OR2X1 U2461 ( .A(n701), .B(read_counter[2]), .Y(n702) );
  OAI2BB1X1 U2462 ( .A0N(n701), .A1N(read_counter[2]), .B0(n702), .Y(N3434) );
  OR2X1 U2463 ( .A(n702), .B(read_counter[3]), .Y(n703) );
  OAI2BB1X1 U2464 ( .A0N(n702), .A1N(read_counter[3]), .B0(n703), .Y(N3435) );
  NOR2X1 U2465 ( .A(read_counter[4]), .B(n703), .Y(n704) );
endmodule


module controller_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module controller_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module controller ( clk, reset, first_block, last_block, output_enable, busy, 
        inner_busy, first_block_core );
  input clk, reset, first_block, last_block;
  output output_enable, busy, inner_busy, first_block_core;
  wire   N13, N14, N24, N25, N26, N27, N28, N29, N30, N45, N46, N47, N48, N49,
         N50, N51, N52, n25, n26, n29, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n27, n28, n30, n31, n32, n33;
  wire   [1:0] state;
  wire   [7:0] counter2;
  wire   [6:0] counter1;

  CLKINVX4 U29 ( .A(reset), .Y(n26) );
  controller_DW01_inc_0 add_97 ( .A(counter2), .SUM({N52, N51, N50, N49, N48, 
        N47, N46, N45}) );
  controller_DW01_inc_1 add_83 ( .A(counter1), .SUM({N30, N29, N28, N27, N26, 
        N25, N24}) );
  DFFTRX1 counter2_reg_0_ ( .D(N45), .RN(n29), .CK(clk), .Q(counter2[0]), .QN(
        n10) );
  DFFTRX1 counter1_reg_1_ ( .D(N25), .RN(n33), .CK(clk), .Q(counter1[1]) );
  DFFTRX1 counter1_reg_0_ ( .D(N24), .RN(n33), .CK(clk), .Q(counter1[0]), .QN(
        n25) );
  DFFTRX1 counter1_reg_3_ ( .D(N27), .RN(n33), .CK(clk), .Q(counter1[3]), .QN(
        n1) );
  DFFTRX1 counter1_reg_5_ ( .D(N29), .RN(n33), .CK(clk), .Q(counter1[5]), .QN(
        n12) );
  DFFTRX1 counter1_reg_6_ ( .D(N30), .RN(n33), .CK(clk), .Q(counter1[6]), .QN(
        n11) );
  DFFTRX1 counter1_reg_2_ ( .D(N26), .RN(n33), .CK(clk), .Q(counter1[2]), .QN(
        n2) );
  DFFTRX1 counter1_reg_4_ ( .D(N28), .RN(n33), .CK(clk), .Q(counter1[4]), .QN(
        n13) );
  DFFHQX1 state_reg_0_ ( .D(N13), .CK(clk), .Q(state[0]) );
  DFFTRX1 counter2_reg_2_ ( .D(N47), .RN(n29), .CK(clk), .Q(counter2[2]), .QN(
        n8) );
  DFFTRX1 counter2_reg_3_ ( .D(N48), .RN(n29), .CK(clk), .Q(counter2[3]), .QN(
        n7) );
  DFFTRX1 counter2_reg_4_ ( .D(N49), .RN(n29), .CK(clk), .Q(counter2[4]), .QN(
        n6) );
  DFFTRX1 counter2_reg_5_ ( .D(N50), .RN(n29), .CK(clk), .Q(counter2[5]), .QN(
        n5) );
  DFFTRX1 counter2_reg_7_ ( .D(N52), .RN(n29), .CK(clk), .Q(counter2[7]), .QN(
        n3) );
  DFFTRX1 counter2_reg_6_ ( .D(N51), .RN(n29), .CK(clk), .Q(counter2[6]), .QN(
        n4) );
  DFFTRX1 counter2_reg_1_ ( .D(N46), .RN(n29), .CK(clk), .Q(counter2[1]), .QN(
        n9) );
  DFFXL state_reg_1_ ( .D(N14), .CK(clk), .Q(state[1]), .QN(n30) );
  NAND3X1 U3 ( .A(n9), .B(n16), .C(n4), .Y(n20) );
  AND4X2 U4 ( .A(n8), .B(n7), .C(n6), .D(n5), .Y(n16) );
  NOR3X1 U5 ( .A(n14), .B(n3), .C(n15), .Y(output_enable) );
  AOI21XL U6 ( .A0(n9), .A1(n16), .B0(n4), .Y(n15) );
  NOR2X1 U7 ( .A(n30), .B(state[0]), .Y(inner_busy) );
  NOR2XL U8 ( .A(state[1]), .B(state[0]), .Y(n22) );
  MXI2XL U9 ( .A(n18), .B(n19), .S0(n3), .Y(n17) );
  NAND4BBXL U10 ( .AN(n4), .BN(n9), .C(n10), .D(n16), .Y(n18) );
  NAND3BXL U11 ( .AN(last_block), .B(n10), .C(n14), .Y(n19) );
  NOR3XL U12 ( .A(n20), .B(n10), .C(n3), .Y(n24) );
  INVXL U13 ( .A(inner_busy), .Y(n23) );
  NAND3XL U14 ( .A(n26), .B(n30), .C(state[0]), .Y(n28) );
  NOR2X1 U15 ( .A(reset), .B(n17), .Y(n29) );
  INVX1 U16 ( .A(n20), .Y(n14) );
  NOR4BBX1 U17 ( .AN(n12), .BN(n13), .C(n21), .D(counter1[1]), .Y(
        first_block_core) );
  NAND4BBX1 U18 ( .AN(n25), .BN(n11), .C(n2), .D(n1), .Y(n21) );
  INVX1 U19 ( .A(n22), .Y(busy) );
  OAI32X1 U20 ( .A0(n23), .A1(reset), .A2(n24), .B0(n27), .B1(n28), .Y(N14) );
  OAI2BB1X1 U21 ( .A0N(n27), .A1N(n33), .B0(n31), .Y(N13) );
  NAND3X1 U22 ( .A(n26), .B(n22), .C(first_block), .Y(n31) );
  INVX1 U23 ( .A(n28), .Y(n33) );
  NAND4X1 U24 ( .A(n13), .B(n12), .C(n25), .D(n32), .Y(n27) );
  NOR4BBX1 U25 ( .AN(n1), .BN(n2), .C(counter1[1]), .D(n11), .Y(n32) );
endmodule


module top ( clk, reset, data, write_enable, last_block, first_block, busy, 
        digest, output_valid );
  input [7:0] data;
  output [3:0] digest;
  input clk, reset, write_enable, last_block, first_block;
  output busy, output_valid;
  wire   inner_busy, first_block_core, output_enable;
  wire   [31:0] Wt;

  message_schedule our_message_schedule ( .clk(clk), .reset(reset), .data(data), .write_enable(write_enable), .inner_busy(inner_busy), .Wt(Wt) );
  hash_core our_hash_core ( .clk(clk), .reset(reset), .Wt(Wt), .inner_busy(
        inner_busy), .first_block_core(first_block_core), .output_enable(
        output_enable), .digest(digest), .output_valid(output_valid) );
  controller our_controller ( .clk(clk), .reset(reset), .first_block(
        first_block), .last_block(last_block), .output_enable(output_enable), 
        .busy(busy), .inner_busy(inner_busy), .first_block_core(
        first_block_core) );
endmodule


module sha256_chip ( clk, reset, data, write_enable, last_block, first_block, 
        busy, digest, output_valid );
  input [7:0] data;
  output [3:0] digest;
  input clk, reset, write_enable, last_block, first_block;
  output busy, output_valid;
  wire   net_clk, net_reset, net_write_enable, net_last_block, net_first_block,
         net_busy, net_output_valid;
  wire   [7:0] net_data;
  wire   [3:0] net_digest;

  PIW PIW_clk ( .PAD(clk), .C(net_clk) );
  PIW PIW_reset ( .PAD(reset), .C(net_reset) );
  PIW PIW_data0 ( .PAD(data[0]), .C(net_data[0]) );
  PIW PIW_data1 ( .PAD(data[1]), .C(net_data[1]) );
  PIW PIW_data2 ( .PAD(data[2]), .C(net_data[2]) );
  PIW PIW_data3 ( .PAD(data[3]), .C(net_data[3]) );
  PIW PIW_data4 ( .PAD(data[4]), .C(net_data[4]) );
  PIW PIW_data5 ( .PAD(data[5]), .C(net_data[5]) );
  PIW PIW_data6 ( .PAD(data[6]), .C(net_data[6]) );
  PIW PIW_data7 ( .PAD(data[7]), .C(net_data[7]) );
  PIW PIW_write_enable ( .PAD(write_enable), .C(net_write_enable) );
  PIW PIW_last_block ( .PAD(last_block), .C(net_last_block) );
  PIW PIW_first_block ( .PAD(first_block), .C(net_first_block) );
  PO8W PO8W_busy ( .I(net_busy), .PAD(busy) );
  PO8W PO8W_digest0 ( .I(net_digest[0]), .PAD(digest[0]) );
  PO8W PO8W_digest1 ( .I(net_digest[1]), .PAD(digest[1]) );
  PO8W PO8W_digest2 ( .I(net_digest[2]), .PAD(digest[2]) );
  PO8W PO8W_digest3 ( .I(net_digest[3]), .PAD(digest[3]) );
  PO8W PO8W_output_valid ( .I(net_output_valid), .PAD(output_valid) );
  top inst_top ( .clk(net_clk), .reset(net_reset), .data(net_data), 
        .write_enable(net_write_enable), .last_block(net_last_block), 
        .first_block(net_first_block), .busy(net_busy), .digest(net_digest), 
        .output_valid(net_output_valid) );
endmodule



module message_schedule_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module message_schedule_DW01_add_2 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1;
  wire   [31:1] carry;

  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX4 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFHX4 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX4 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX4 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX4 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX4 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  INVX4 U1 ( .A(n1), .Y(carry[1]) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X4 U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module message_schedule_DW01_add_4 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215;

  OAI21XL U2 ( .A0(n151), .A1(n13), .B0(n152), .Y(n150) );
  OAI21XL U3 ( .A0(n9), .A1(n157), .B0(n158), .Y(n154) );
  NAND2X2 U4 ( .A(n145), .B(n146), .Y(n122) );
  OAI21X1 U5 ( .A0(n160), .A1(n5), .B0(n149), .Y(n145) );
  INVX1 U6 ( .A(n150), .Y(n149) );
  NAND2X1 U7 ( .A(n94), .B(n95), .Y(n74) );
  OR2X2 U8 ( .A(A[5]), .B(B[5]), .Y(n36) );
  NAND2X1 U9 ( .A(B[4]), .B(A[4]), .Y(n39) );
  INVX1 U10 ( .A(n165), .Y(n203) );
  NOR2X1 U11 ( .A(A[9]), .B(B[9]), .Y(n8) );
  INVX1 U12 ( .A(n189), .Y(n194) );
  NAND2X1 U13 ( .A(n142), .B(n132), .Y(n140) );
  NAND2X1 U14 ( .A(n115), .B(n110), .Y(n113) );
  OAI21XL U15 ( .A0(n58), .A1(n59), .B0(n60), .Y(n56) );
  OAI21X4 U16 ( .A0(n204), .A1(n205), .B0(n26), .Y(n165) );
  NAND3BX4 U17 ( .AN(n170), .B(n48), .C(n168), .Y(n38) );
  NAND3X2 U18 ( .A(n210), .B(n64), .C(n211), .Y(n168) );
  BUFX3 U19 ( .A(n118), .Y(n1) );
  OAI21X4 U20 ( .A0(n10), .A1(n184), .B0(n23), .Y(n18) );
  INVX4 U21 ( .A(n21), .Y(n184) );
  NOR2XL U22 ( .A(n40), .B(n45), .Y(n214) );
  OR2X1 U23 ( .A(A[6]), .B(B[6]), .Y(n206) );
  NAND2XL U24 ( .A(B[9]), .B(A[9]), .Y(n20) );
  OR2XL U25 ( .A(A[4]), .B(B[4]), .Y(n37) );
  XOR2X1 U26 ( .A(n67), .B(n59), .Y(SUM[29]) );
  OR2X1 U27 ( .A(A[1]), .B(B[1]), .Y(n64) );
  XOR2X2 U28 ( .A(n56), .B(n6), .Y(SUM[30]) );
  NOR2BXL U29 ( .AN(n48), .B(n49), .Y(n47) );
  NAND2X1 U30 ( .A(B[1]), .B(A[1]), .Y(n65) );
  NAND2X1 U31 ( .A(B[6]), .B(A[6]), .Y(n30) );
  NAND2XL U32 ( .A(B[2]), .B(A[2]), .Y(n52) );
  NAND2XL U33 ( .A(B[13]), .B(A[13]), .Y(n158) );
  OAI21XL U34 ( .A0(n139), .A1(n128), .B0(n127), .Y(n137) );
  OAI21XL U35 ( .A0(n50), .A1(n51), .B0(n52), .Y(n46) );
  NOR2XL U36 ( .A(n39), .B(n40), .Y(n33) );
  INVX1 U37 ( .A(n156), .Y(n155) );
  XOR2X1 U38 ( .A(n113), .B(n7), .Y(SUM[22]) );
  NOR2X1 U39 ( .A(n49), .B(n51), .Y(n210) );
  NOR2X1 U40 ( .A(A[13]), .B(B[13]), .Y(n9) );
  NAND2XL U41 ( .A(B[5]), .B(A[5]), .Y(n34) );
  NAND2X1 U42 ( .A(B[8]), .B(A[8]), .Y(n23) );
  OAI2BB1X2 U43 ( .A0N(n202), .A1N(n38), .B0(n203), .Y(n21) );
  CLKINVX3 U44 ( .A(n159), .Y(n202) );
  OAI21X2 U45 ( .A0(n12), .A1(n181), .B0(n157), .Y(n179) );
  INVX2 U46 ( .A(n182), .Y(n181) );
  OAI21X2 U47 ( .A0(n8), .A1(n201), .B0(n20), .Y(n199) );
  INVX2 U48 ( .A(n18), .Y(n201) );
  OAI21X2 U49 ( .A0(n178), .A1(n9), .B0(n158), .Y(n176) );
  INVX2 U50 ( .A(n179), .Y(n178) );
  NAND2XL U51 ( .A(n206), .B(n207), .Y(n205) );
  NOR2BXL U52 ( .AN(n156), .B(n173), .Y(n177) );
  XOR2X2 U53 ( .A(n174), .B(n175), .Y(SUM[15]) );
  NOR2BXL U54 ( .AN(n152), .B(n13), .Y(n175) );
  INVXL U55 ( .A(n212), .Y(n49) );
  NOR2BX1 U56 ( .AN(n133), .B(n125), .Y(n124) );
  XNOR2X1 U57 ( .A(n89), .B(n2), .Y(SUM[26]) );
  NAND2X1 U58 ( .A(n82), .B(n77), .Y(n2) );
  NOR2BXL U59 ( .AN(n39), .B(n45), .Y(n44) );
  NOR2BXL U60 ( .AN(n30), .B(n29), .Y(n32) );
  NOR2BXL U61 ( .AN(n132), .B(n130), .Y(n144) );
  NOR2BXL U62 ( .AN(n23), .B(n10), .Y(n22) );
  INVXL U63 ( .A(n161), .Y(n166) );
  AOI21XL U64 ( .A0(n167), .A1(n168), .B0(n159), .Y(n164) );
  NOR2XL U65 ( .A(n169), .B(n170), .Y(n167) );
  NAND3XL U66 ( .A(n36), .B(n37), .C(n38), .Y(n35) );
  NAND2X2 U67 ( .A(n1), .B(n119), .Y(n98) );
  XNOR2X1 U68 ( .A(n94), .B(n3), .Y(SUM[24]) );
  NAND2X1 U69 ( .A(n85), .B(n95), .Y(n3) );
  XNOR2X1 U70 ( .A(n68), .B(n4), .Y(SUM[28]) );
  NAND2X1 U71 ( .A(n71), .B(n69), .Y(n4) );
  NAND2XL U72 ( .A(n52), .B(n66), .Y(n62) );
  NAND2XL U73 ( .A(n56), .B(n57), .Y(n55) );
  NAND2XL U74 ( .A(B[3]), .B(A[3]), .Y(n48) );
  NAND2XL U75 ( .A(B[7]), .B(A[7]), .Y(n26) );
  NAND2XL U76 ( .A(B[10]), .B(A[10]), .Y(n191) );
  NAND2XL U77 ( .A(B[11]), .B(A[11]), .Y(n188) );
  NOR2XL U78 ( .A(A[0]), .B(B[0]), .Y(n15) );
  AND2X1 U79 ( .A(B[0]), .B(A[0]), .Y(n16) );
  NOR2XL U80 ( .A(A[12]), .B(B[12]), .Y(n12) );
  NAND2XL U81 ( .A(B[0]), .B(A[0]), .Y(n17) );
  NAND2XL U82 ( .A(B[17]), .B(A[17]), .Y(n132) );
  NAND2XL U83 ( .A(B[15]), .B(A[15]), .Y(n152) );
  NAND3XL U84 ( .A(A[0]), .B(B[0]), .C(n64), .Y(n63) );
  AND2X1 U85 ( .A(n65), .B(n63), .Y(n50) );
  OAI21XL U86 ( .A0(n184), .A1(n161), .B0(n162), .Y(n182) );
  NAND2X1 U87 ( .A(n214), .B(n215), .Y(n159) );
  NOR2X1 U88 ( .A(n27), .B(n29), .Y(n215) );
  AND2X2 U89 ( .A(n162), .B(n163), .Y(n5) );
  INVX1 U90 ( .A(n36), .Y(n40) );
  INVX1 U91 ( .A(n206), .Y(n29) );
  AOI21X1 U92 ( .A0(n185), .A1(n186), .B0(n187), .Y(n162) );
  INVX1 U93 ( .A(n188), .Y(n187) );
  OAI2BB1X1 U94 ( .A0N(n189), .A1N(n190), .B0(n191), .Y(n186) );
  OAI21XL U95 ( .A0(n8), .A1(n23), .B0(n20), .Y(n190) );
  NOR2X1 U96 ( .A(n208), .B(n209), .Y(n204) );
  NAND2X1 U97 ( .A(n30), .B(n34), .Y(n209) );
  INVX1 U98 ( .A(n37), .Y(n45) );
  INVX1 U99 ( .A(n66), .Y(n51) );
  INVX1 U100 ( .A(n207), .Y(n27) );
  XOR2X1 U101 ( .A(n199), .B(n200), .Y(SUM[10]) );
  NOR2BX1 U102 ( .AN(n191), .B(n194), .Y(n200) );
  XOR2X1 U103 ( .A(n18), .B(n19), .Y(SUM[9]) );
  NOR2BX1 U104 ( .AN(n20), .B(n8), .Y(n19) );
  XOR2X1 U105 ( .A(n179), .B(n180), .Y(SUM[13]) );
  NOR2BX1 U106 ( .AN(n158), .B(n9), .Y(n180) );
  XOR2X1 U107 ( .A(n176), .B(n177), .Y(SUM[14]) );
  XOR2X1 U108 ( .A(n24), .B(n25), .Y(SUM[7]) );
  NOR2BX1 U109 ( .AN(n26), .B(n27), .Y(n25) );
  OAI21XL U110 ( .A0(n28), .A1(n29), .B0(n30), .Y(n24) );
  INVX1 U111 ( .A(n31), .Y(n28) );
  XOR2X1 U112 ( .A(n196), .B(n197), .Y(SUM[11]) );
  NOR2BX1 U113 ( .AN(n188), .B(n195), .Y(n197) );
  OAI21XL U114 ( .A0(n198), .A1(n194), .B0(n191), .Y(n196) );
  INVX1 U115 ( .A(n199), .Y(n198) );
  OAI2BB1X1 U116 ( .A0N(n153), .A1N(n176), .B0(n156), .Y(n174) );
  NAND3BX1 U117 ( .AN(n33), .B(n34), .C(n35), .Y(n31) );
  NOR2X1 U118 ( .A(n40), .B(n39), .Y(n208) );
  INVX1 U119 ( .A(n213), .Y(n170) );
  NAND2BX1 U120 ( .AN(n52), .B(n212), .Y(n213) );
  AND2X2 U121 ( .A(n54), .B(n57), .Y(n6) );
  AOI21X1 U122 ( .A0(n68), .A1(n69), .B0(n70), .Y(n59) );
  INVX1 U123 ( .A(n71), .Y(n70) );
  OAI21XL U124 ( .A0(n122), .A1(n123), .B0(n124), .Y(n118) );
  NAND3BX1 U125 ( .AN(n11), .B(n134), .C(n135), .Y(n123) );
  INVX1 U126 ( .A(n61), .Y(n58) );
  INVX1 U127 ( .A(n134), .Y(n128) );
  XOR2X1 U128 ( .A(n92), .B(n93), .Y(SUM[25]) );
  NOR2BX1 U129 ( .AN(n86), .B(n84), .Y(n93) );
  NAND2X1 U130 ( .A(n60), .B(n61), .Y(n67) );
  XOR2X1 U131 ( .A(n41), .B(n42), .Y(SUM[5]) );
  NAND2X1 U132 ( .A(n36), .B(n34), .Y(n41) );
  AOI21X1 U133 ( .A0(n38), .A1(n37), .B0(n43), .Y(n42) );
  INVX1 U134 ( .A(n39), .Y(n43) );
  INVX1 U135 ( .A(n135), .Y(n130) );
  INVX1 U136 ( .A(n153), .Y(n173) );
  INVX1 U137 ( .A(n185), .Y(n195) );
  XOR2X1 U138 ( .A(n46), .B(n47), .Y(SUM[3]) );
  XOR2X1 U139 ( .A(n38), .B(n44), .Y(SUM[4]) );
  AOI21X1 U140 ( .A0(n126), .A1(n127), .B0(n11), .Y(n125) );
  NAND2BX1 U141 ( .AN(n128), .B(n129), .Y(n126) );
  OAI21XL U142 ( .A0(n130), .A1(n131), .B0(n132), .Y(n129) );
  XOR2X1 U143 ( .A(n1), .B(n120), .Y(SUM[20]) );
  NOR2BX1 U144 ( .AN(n109), .B(n121), .Y(n120) );
  INVX1 U145 ( .A(n119), .Y(n121) );
  XOR2X1 U146 ( .A(n182), .B(n183), .Y(SUM[12]) );
  NOR2BX1 U147 ( .AN(n157), .B(n12), .Y(n183) );
  XOR2X1 U148 ( .A(n31), .B(n32), .Y(SUM[6]) );
  XOR2X1 U149 ( .A(n137), .B(n138), .Y(SUM[19]) );
  NOR2BX1 U150 ( .AN(n133), .B(n11), .Y(n138) );
  INVX1 U151 ( .A(n140), .Y(n139) );
  XOR2X1 U152 ( .A(n143), .B(n144), .Y(SUM[17]) );
  XOR2X1 U153 ( .A(n116), .B(n117), .Y(SUM[21]) );
  NOR2BX1 U154 ( .AN(n110), .B(n108), .Y(n117) );
  XOR2X1 U155 ( .A(n62), .B(n50), .Y(SUM[2]) );
  XOR2X1 U156 ( .A(n111), .B(n112), .Y(SUM[23]) );
  NAND2X1 U157 ( .A(n104), .B(n100), .Y(n111) );
  AOI21X1 U158 ( .A0(n101), .A1(n113), .B0(n114), .Y(n112) );
  INVX1 U159 ( .A(n106), .Y(n114) );
  XOR2X1 U160 ( .A(n87), .B(n88), .Y(SUM[27]) );
  NAND2X1 U161 ( .A(n80), .B(n76), .Y(n87) );
  AOI21X1 U162 ( .A0(n77), .A1(n89), .B0(n90), .Y(n88) );
  INVX1 U163 ( .A(n82), .Y(n90) );
  XOR2X1 U164 ( .A(n21), .B(n22), .Y(SUM[8]) );
  XOR2X1 U165 ( .A(n140), .B(n141), .Y(SUM[18]) );
  NOR2BX1 U166 ( .AN(n127), .B(n128), .Y(n141) );
  XOR2X1 U167 ( .A(n145), .B(n147), .Y(SUM[16]) );
  NOR2BX1 U168 ( .AN(n131), .B(n148), .Y(n147) );
  INVX1 U169 ( .A(n146), .Y(n148) );
  AND2X2 U170 ( .A(n106), .B(n101), .Y(n7) );
  NAND2X1 U171 ( .A(n74), .B(n85), .Y(n92) );
  NAND2X1 U172 ( .A(n122), .B(n131), .Y(n143) );
  NAND2X1 U173 ( .A(n98), .B(n109), .Y(n116) );
  OAI21XL U174 ( .A0(n164), .A1(n165), .B0(n166), .Y(n163) );
  AOI21X1 U175 ( .A0(n153), .A1(n154), .B0(n155), .Y(n151) );
  NAND2X1 U176 ( .A(n99), .B(n116), .Y(n115) );
  NAND2X1 U177 ( .A(n91), .B(n86), .Y(n89) );
  NAND2X1 U178 ( .A(n75), .B(n92), .Y(n91) );
  NAND2X1 U179 ( .A(n72), .B(n73), .Y(n68) );
  AOI21X1 U180 ( .A0(n78), .A1(n76), .B0(n79), .Y(n72) );
  NAND4BXL U181 ( .AN(n74), .B(n75), .C(n76), .D(n77), .Y(n73) );
  INVX1 U182 ( .A(n80), .Y(n79) );
  NAND2X1 U183 ( .A(n96), .B(n97), .Y(n94) );
  AOI21X1 U184 ( .A0(n102), .A1(n100), .B0(n103), .Y(n96) );
  NAND4BXL U185 ( .AN(n98), .B(n99), .C(n100), .D(n101), .Y(n97) );
  INVX1 U186 ( .A(n104), .Y(n103) );
  NAND2X1 U187 ( .A(n192), .B(n193), .Y(n161) );
  NOR2X1 U188 ( .A(n194), .B(n195), .Y(n192) );
  NOR2X1 U189 ( .A(n10), .B(n8), .Y(n193) );
  INVX1 U190 ( .A(n48), .Y(n169) );
  NAND2X1 U191 ( .A(n135), .B(n143), .Y(n142) );
  NAND2X1 U192 ( .A(n65), .B(n64), .Y(n136) );
  NAND2X1 U193 ( .A(n171), .B(n172), .Y(n160) );
  NOR2X1 U194 ( .A(n13), .B(n173), .Y(n172) );
  NOR2X1 U195 ( .A(n9), .B(n12), .Y(n171) );
  INVX1 U196 ( .A(n99), .Y(n108) );
  NAND2X1 U197 ( .A(n105), .B(n106), .Y(n102) );
  NAND2X1 U198 ( .A(n101), .B(n107), .Y(n105) );
  OAI21XL U199 ( .A0(n108), .A1(n109), .B0(n110), .Y(n107) );
  INVX1 U200 ( .A(n75), .Y(n84) );
  NAND2X1 U201 ( .A(n81), .B(n82), .Y(n78) );
  NAND2X1 U202 ( .A(n77), .B(n83), .Y(n81) );
  OAI21XL U203 ( .A0(n84), .A1(n85), .B0(n86), .Y(n83) );
  OAI2BB1X1 U204 ( .A0N(B[0]), .A1N(A[0]), .B0(n65), .Y(n211) );
  OR2X2 U205 ( .A(A[3]), .B(B[3]), .Y(n212) );
  OR2X2 U206 ( .A(A[2]), .B(B[2]), .Y(n66) );
  OR2X2 U207 ( .A(A[7]), .B(B[7]), .Y(n207) );
  NOR2X1 U208 ( .A(A[8]), .B(B[8]), .Y(n10) );
  NOR2X1 U209 ( .A(A[19]), .B(B[19]), .Y(n11) );
  NAND2X1 U210 ( .A(B[16]), .B(A[16]), .Y(n131) );
  NAND2X1 U211 ( .A(B[12]), .B(A[12]), .Y(n157) );
  NAND2X1 U212 ( .A(B[14]), .B(A[14]), .Y(n156) );
  OR2X2 U213 ( .A(A[17]), .B(B[17]), .Y(n135) );
  OR2X2 U214 ( .A(A[14]), .B(B[14]), .Y(n153) );
  OR2X2 U215 ( .A(A[11]), .B(B[11]), .Y(n185) );
  OR2X2 U216 ( .A(A[18]), .B(B[18]), .Y(n134) );
  XOR2X1 U217 ( .A(n17), .B(n136), .Y(SUM[1]) );
  OR2X2 U218 ( .A(A[10]), .B(B[10]), .Y(n189) );
  NOR2X1 U219 ( .A(A[15]), .B(B[15]), .Y(n13) );
  OR2X2 U220 ( .A(A[22]), .B(B[22]), .Y(n101) );
  NAND2X1 U221 ( .A(B[20]), .B(A[20]), .Y(n109) );
  NAND2X1 U222 ( .A(B[18]), .B(A[18]), .Y(n127) );
  NAND2X1 U223 ( .A(B[22]), .B(A[22]), .Y(n106) );
  OR2X2 U224 ( .A(A[23]), .B(B[23]), .Y(n100) );
  NAND2X1 U225 ( .A(B[21]), .B(A[21]), .Y(n110) );
  OR2X2 U226 ( .A(A[21]), .B(B[21]), .Y(n99) );
  NOR2X1 U227 ( .A(n15), .B(n16), .Y(SUM[0]) );
  NAND2X1 U228 ( .A(B[23]), .B(A[23]), .Y(n104) );
  NAND2X1 U229 ( .A(B[19]), .B(A[19]), .Y(n133) );
  OR2X2 U230 ( .A(A[16]), .B(B[16]), .Y(n146) );
  OR2X2 U231 ( .A(A[20]), .B(B[20]), .Y(n119) );
  OR2X2 U232 ( .A(A[26]), .B(B[26]), .Y(n77) );
  NAND2X1 U233 ( .A(B[24]), .B(A[24]), .Y(n85) );
  NAND2X1 U234 ( .A(B[26]), .B(A[26]), .Y(n82) );
  OR2X2 U235 ( .A(A[27]), .B(B[27]), .Y(n76) );
  NAND2X1 U236 ( .A(B[25]), .B(A[25]), .Y(n86) );
  OR2X2 U237 ( .A(A[25]), .B(B[25]), .Y(n75) );
  NAND2X1 U238 ( .A(B[27]), .B(A[27]), .Y(n80) );
  OR2X2 U239 ( .A(A[24]), .B(B[24]), .Y(n95) );
  NAND2X1 U240 ( .A(B[30]), .B(A[30]), .Y(n54) );
  NAND2X1 U241 ( .A(B[29]), .B(A[29]), .Y(n60) );
  NAND2X1 U242 ( .A(B[28]), .B(A[28]), .Y(n71) );
  OR2X2 U243 ( .A(A[28]), .B(B[28]), .Y(n69) );
  OR2X2 U244 ( .A(A[30]), .B(B[30]), .Y(n57) );
  OR2X2 U245 ( .A(A[29]), .B(B[29]), .Y(n61) );
  XOR3X2 U246 ( .A(B[31]), .B(A[31]), .C(n53), .Y(SUM[31]) );
  NAND2X1 U247 ( .A(n54), .B(n55), .Y(n53) );
endmodule


module message_schedule_DW01_add_5 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217;

  OAI21X1 U2 ( .A0(n184), .A1(n6), .B0(n163), .Y(n182) );
  XOR2X4 U3 ( .A(n85), .B(n86), .Y(SUM[27]) );
  OAI21X2 U4 ( .A0(n87), .A1(n82), .B0(n88), .Y(n85) );
  NAND2X2 U5 ( .A(n1), .B(n2), .Y(n3) );
  NAND2X2 U6 ( .A(n123), .B(n124), .Y(n100) );
  OR2X2 U7 ( .A(A[28]), .B(B[28]), .Y(n68) );
  INVX1 U8 ( .A(n206), .Y(n199) );
  NAND2X1 U9 ( .A(n91), .B(n79), .Y(n89) );
  NAND2X2 U10 ( .A(n70), .B(n95), .Y(n93) );
  OAI211X1 U11 ( .A0(n77), .A1(n78), .B0(n79), .C0(n80), .Y(n74) );
  OAI21X2 U12 ( .A0(n48), .A1(n49), .B0(n50), .Y(n47) );
  OAI21X1 U13 ( .A0(n33), .A1(n175), .B0(n210), .Y(n15) );
  OR2X2 U14 ( .A(A[25]), .B(B[25]), .Y(n92) );
  NOR2X1 U15 ( .A(A[25]), .B(B[25]), .Y(n77) );
  NOR2BX2 U16 ( .AN(n52), .B(n51), .Y(n45) );
  XNOR2X4 U17 ( .A(B[31]), .B(A[31]), .Y(n43) );
  NAND2X1 U18 ( .A(n52), .B(n56), .Y(n66) );
  NAND2X1 U19 ( .A(B[27]), .B(A[27]), .Y(n76) );
  NAND3BX1 U20 ( .AN(n77), .B(n83), .C(n84), .Y(n71) );
  XOR2X4 U21 ( .A(n43), .B(n44), .Y(SUM[31]) );
  NAND2X2 U22 ( .A(B[28]), .B(A[28]), .Y(n59) );
  NAND2X2 U23 ( .A(B[30]), .B(A[30]), .Y(n50) );
  NAND2X1 U24 ( .A(B[29]), .B(A[29]), .Y(n56) );
  XOR2X2 U25 ( .A(n66), .B(n67), .Y(SUM[29]) );
  AOI21X4 U26 ( .A0(n45), .A1(n46), .B0(n47), .Y(n44) );
  OAI21X4 U27 ( .A0(n57), .A1(n58), .B0(n59), .Y(n46) );
  INVX3 U28 ( .A(n76), .Y(n75) );
  INVX4 U29 ( .A(n60), .Y(n58) );
  OAI2BB1X2 U30 ( .A0N(n60), .A1N(n68), .B0(n59), .Y(n4) );
  AOI21X4 U31 ( .A0(n73), .A1(n74), .B0(n75), .Y(n72) );
  NOR2X2 U32 ( .A(n81), .B(n82), .Y(n73) );
  AOI21X2 U33 ( .A0(n52), .A1(n46), .B0(n55), .Y(n54) );
  NAND2X4 U34 ( .A(n3), .B(n102), .Y(n96) );
  CLKINVX2 U35 ( .A(n100), .Y(n1) );
  INVX1 U36 ( .A(n101), .Y(n2) );
  AOI21X2 U37 ( .A0(n103), .A1(n104), .B0(n105), .Y(n102) );
  NAND2X4 U38 ( .A(n96), .B(n97), .Y(n70) );
  OAI21X4 U39 ( .A0(n70), .A1(n71), .B0(n72), .Y(n60) );
  NAND2XL U40 ( .A(B[9]), .B(A[9]), .Y(n14) );
  OAI21XL U41 ( .A0(n193), .A1(n194), .B0(n195), .Y(n192) );
  INVX2 U42 ( .A(n4), .Y(n67) );
  OR2X2 U43 ( .A(A[10]), .B(B[10]), .Y(n201) );
  NAND2X1 U44 ( .A(B[13]), .B(A[13]), .Y(n163) );
  NAND2X1 U45 ( .A(B[14]), .B(A[14]), .Y(n164) );
  NOR2X1 U46 ( .A(A[13]), .B(B[13]), .Y(n6) );
  NOR2X2 U47 ( .A(A[30]), .B(B[30]), .Y(n51) );
  NAND2X2 U48 ( .A(n156), .B(n157), .Y(n130) );
  OAI21X1 U49 ( .A0(n171), .A1(n167), .B0(n172), .Y(n170) );
  OAI2BB1XL U50 ( .A0N(n191), .A1N(n15), .B0(n172), .Y(n189) );
  INVXL U51 ( .A(n174), .Y(n210) );
  NAND3BXL U52 ( .AN(n107), .B(n113), .C(n114), .Y(n101) );
  INVX2 U53 ( .A(n177), .Y(n166) );
  NAND4BBXL U54 ( .AN(n18), .BN(n7), .C(n201), .D(n196), .Y(n167) );
  INVXL U55 ( .A(n56), .Y(n55) );
  NAND4BBXL U56 ( .AN(n8), .BN(n9), .C(n28), .D(n212), .Y(n175) );
  NAND2XL U57 ( .A(n130), .B(n133), .Y(n154) );
  NAND2XL U58 ( .A(n100), .B(n108), .Y(n121) );
  NAND2XL U59 ( .A(n209), .B(n17), .Y(n12) );
  NAND2XL U60 ( .A(n15), .B(n202), .Y(n209) );
  AOI21XL U61 ( .A0(n201), .A1(n205), .B0(n199), .Y(n204) );
  NOR2BXL U62 ( .AN(n161), .B(n165), .Y(n180) );
  NAND2XL U63 ( .A(n133), .B(n134), .Y(n129) );
  NOR2BXL U64 ( .AN(n142), .B(n132), .Y(n150) );
  NOR2BXL U65 ( .AN(n164), .B(n166), .Y(n183) );
  NOR2BXL U66 ( .AN(n206), .B(n200), .Y(n207) );
  INVXL U67 ( .A(n176), .Y(n187) );
  NAND2XL U68 ( .A(n195), .B(n196), .Y(n203) );
  INVXL U69 ( .A(n97), .Y(n99) );
  NOR2BXL U70 ( .AN(n14), .B(n7), .Y(n13) );
  NOR2BXL U71 ( .AN(n141), .B(n139), .Y(n153) );
  NOR2BXL U72 ( .AN(n21), .B(n22), .Y(n20) );
  INVXL U73 ( .A(n124), .Y(n126) );
  AND2X1 U74 ( .A(n140), .B(n133), .Y(n155) );
  NOR2BXL U75 ( .AN(n30), .B(n8), .Y(n32) );
  INVXL U76 ( .A(n28), .Y(n24) );
  NOR2BXL U77 ( .AN(n38), .B(n10), .Y(n37) );
  NOR2BXL U78 ( .AN(n65), .B(n144), .Y(n143) );
  NAND2XL U79 ( .A(B[11]), .B(A[11]), .Y(n195) );
  NAND2XL U80 ( .A(B[15]), .B(A[15]), .Y(n161) );
  NAND2XL U81 ( .A(B[18]), .B(A[18]), .Y(n142) );
  NAND2XL U82 ( .A(B[22]), .B(A[22]), .Y(n110) );
  NAND2XL U83 ( .A(B[19]), .B(A[19]), .Y(n138) );
  NAND2XL U84 ( .A(B[23]), .B(A[23]), .Y(n106) );
  NAND2XL U85 ( .A(B[7]), .B(A[7]), .Y(n21) );
  NAND2XL U86 ( .A(B[24]), .B(A[24]), .Y(n95) );
  NAND2XL U87 ( .A(B[3]), .B(A[3]), .Y(n38) );
  OR2XL U88 ( .A(A[2]), .B(B[2]), .Y(n62) );
  XOR2X2 U89 ( .A(n53), .B(n54), .Y(SUM[30]) );
  XNOR2X1 U90 ( .A(B[30]), .B(A[30]), .Y(n53) );
  NOR2BXL U91 ( .AN(n138), .B(n5), .Y(n147) );
  NOR2BXL U92 ( .AN(n79), .B(n77), .Y(n94) );
  NOR2BXL U93 ( .AN(n106), .B(n111), .Y(n116) );
  NOR2BXL U94 ( .AN(n110), .B(n112), .Y(n119) );
  NOR2BXL U95 ( .AN(n109), .B(n107), .Y(n122) );
  INVX1 U96 ( .A(n173), .Y(n33) );
  NOR2X1 U97 ( .A(n111), .B(n112), .Y(n103) );
  NAND2BX1 U98 ( .AN(n169), .B(n170), .Y(n156) );
  AOI21X1 U99 ( .A0(n158), .A1(n159), .B0(n160), .Y(n157) );
  NOR2X1 U100 ( .A(n165), .B(n166), .Y(n158) );
  AOI21X1 U101 ( .A0(n168), .A1(n173), .B0(n174), .Y(n171) );
  INVX1 U102 ( .A(n175), .Y(n168) );
  INVX1 U103 ( .A(n167), .Y(n191) );
  OAI211X1 U104 ( .A0(n107), .A1(n108), .B0(n109), .C0(n110), .Y(n104) );
  INVX1 U105 ( .A(n113), .Y(n112) );
  INVX1 U106 ( .A(n106), .Y(n105) );
  INVX1 U107 ( .A(n120), .Y(n107) );
  INVX1 U108 ( .A(n114), .Y(n111) );
  INVX1 U109 ( .A(n89), .Y(n87) );
  NAND2X1 U110 ( .A(n127), .B(n128), .Y(n123) );
  AOI21X1 U111 ( .A0(n135), .A1(n136), .B0(n137), .Y(n127) );
  NAND3BX1 U112 ( .AN(n129), .B(n130), .C(n131), .Y(n128) );
  INVX1 U113 ( .A(n138), .Y(n137) );
  NAND2X1 U114 ( .A(n92), .B(n93), .Y(n91) );
  NOR2X1 U115 ( .A(n132), .B(n5), .Y(n131) );
  OAI211X1 U116 ( .A0(n6), .A1(n162), .B0(n163), .C0(n164), .Y(n159) );
  OAI211X1 U117 ( .A0(n139), .A1(n140), .B0(n141), .C0(n142), .Y(n136) );
  INVX1 U118 ( .A(n148), .Y(n132) );
  INVX1 U119 ( .A(n134), .Y(n139) );
  INVX1 U120 ( .A(n178), .Y(n165) );
  OAI21XL U121 ( .A0(n117), .A1(n112), .B0(n110), .Y(n115) );
  INVX1 U122 ( .A(n118), .Y(n117) );
  NOR2X1 U123 ( .A(n5), .B(n132), .Y(n135) );
  OAI2BB1X1 U124 ( .A0N(n120), .A1N(n121), .B0(n109), .Y(n118) );
  NAND4BXL U125 ( .AN(n6), .B(n176), .C(n177), .D(n178), .Y(n169) );
  OAI21XL U126 ( .A0(n211), .A1(n22), .B0(n21), .Y(n174) );
  AOI21X1 U127 ( .A0(n28), .A1(n213), .B0(n214), .Y(n211) );
  INVX1 U128 ( .A(n25), .Y(n214) );
  OAI21XL U129 ( .A0(n8), .A1(n34), .B0(n30), .Y(n213) );
  OAI21XL U130 ( .A0(n151), .A1(n139), .B0(n141), .Y(n149) );
  INVX1 U131 ( .A(n152), .Y(n151) );
  INVX1 U132 ( .A(n201), .Y(n200) );
  INVX1 U133 ( .A(n212), .Y(n22) );
  INVX1 U134 ( .A(n192), .Y(n172) );
  INVX1 U135 ( .A(n196), .Y(n194) );
  AOI21X1 U136 ( .A0(n197), .A1(n198), .B0(n199), .Y(n193) );
  NOR2X1 U137 ( .A(n7), .B(n200), .Y(n197) );
  NAND2X1 U138 ( .A(n154), .B(n140), .Y(n152) );
  NAND2X1 U139 ( .A(n17), .B(n14), .Y(n198) );
  OAI2BB1X1 U140 ( .A0N(n148), .A1N(n149), .B0(n142), .Y(n146) );
  INVX1 U141 ( .A(n161), .Y(n160) );
  INVX1 U142 ( .A(n185), .Y(n184) );
  OAI21XL U143 ( .A0(n215), .A1(n10), .B0(n38), .Y(n173) );
  AOI21X1 U144 ( .A0(n62), .A1(n216), .B0(n217), .Y(n215) );
  INVX1 U145 ( .A(n41), .Y(n217) );
  OAI21XL U146 ( .A0(n144), .A1(n145), .B0(n65), .Y(n216) );
  OAI21XL U147 ( .A0(n187), .A1(n188), .B0(n162), .Y(n185) );
  INVX1 U148 ( .A(n189), .Y(n188) );
  INVX1 U149 ( .A(n63), .Y(n144) );
  OAI21XL U150 ( .A0(n181), .A1(n166), .B0(n164), .Y(n179) );
  INVX1 U151 ( .A(n182), .Y(n181) );
  INVX1 U152 ( .A(n202), .Y(n18) );
  OAI21XL U153 ( .A0(n208), .A1(n7), .B0(n14), .Y(n205) );
  INVX1 U154 ( .A(n12), .Y(n208) );
  OAI21XL U155 ( .A0(n29), .A1(n8), .B0(n30), .Y(n26) );
  INVX1 U156 ( .A(n31), .Y(n29) );
  OAI21XL U157 ( .A0(n9), .A1(n33), .B0(n34), .Y(n31) );
  NOR2BX1 U158 ( .AN(n163), .B(n6), .Y(n186) );
  NOR2BX1 U159 ( .AN(n162), .B(n187), .Y(n190) );
  OAI21XL U160 ( .A0(n23), .A1(n24), .B0(n25), .Y(n19) );
  INVX1 U161 ( .A(n26), .Y(n23) );
  INVX1 U162 ( .A(n62), .Y(n40) );
  NOR2BX1 U163 ( .AN(n34), .B(n9), .Y(n35) );
  NOR2BX1 U164 ( .AN(n25), .B(n24), .Y(n27) );
  NOR2BX1 U165 ( .AN(n41), .B(n40), .Y(n61) );
  NOR2BX1 U166 ( .AN(n17), .B(n18), .Y(n16) );
  OAI21XL U167 ( .A0(n39), .A1(n40), .B0(n41), .Y(n36) );
  INVX1 U168 ( .A(n42), .Y(n39) );
  OAI2BB1X1 U169 ( .A0N(n63), .A1N(n64), .B0(n65), .Y(n42) );
  INVX1 U170 ( .A(n145), .Y(n64) );
  NOR2X1 U171 ( .A(A[19]), .B(B[19]), .Y(n5) );
  NAND2XL U172 ( .A(A[29]), .B(B[29]), .Y(n49) );
  NAND2X1 U173 ( .A(B[25]), .B(A[25]), .Y(n79) );
  NAND2XL U174 ( .A(B[26]), .B(A[26]), .Y(n88) );
  OR2X2 U175 ( .A(A[24]), .B(B[24]), .Y(n97) );
  OR2X2 U176 ( .A(A[23]), .B(B[23]), .Y(n114) );
  OR2X2 U177 ( .A(A[22]), .B(B[22]), .Y(n113) );
  NAND2XL U178 ( .A(B[26]), .B(A[26]), .Y(n80) );
  NAND2X1 U179 ( .A(A[24]), .B(B[24]), .Y(n78) );
  OR2X2 U180 ( .A(A[21]), .B(B[21]), .Y(n120) );
  NAND2X1 U181 ( .A(B[16]), .B(A[16]), .Y(n140) );
  NAND2X1 U182 ( .A(B[20]), .B(A[20]), .Y(n108) );
  NAND2X1 U183 ( .A(B[17]), .B(A[17]), .Y(n141) );
  NAND2X1 U184 ( .A(B[21]), .B(A[21]), .Y(n109) );
  OR2X2 U185 ( .A(A[16]), .B(B[16]), .Y(n133) );
  OR2X2 U186 ( .A(A[15]), .B(B[15]), .Y(n178) );
  OR2X2 U187 ( .A(A[14]), .B(B[14]), .Y(n177) );
  OR2X2 U188 ( .A(A[17]), .B(B[17]), .Y(n134) );
  OR2X2 U189 ( .A(A[20]), .B(B[20]), .Y(n124) );
  OR2X2 U190 ( .A(A[18]), .B(B[18]), .Y(n148) );
  NOR2X1 U191 ( .A(A[9]), .B(B[9]), .Y(n7) );
  NAND2X1 U192 ( .A(B[12]), .B(A[12]), .Y(n162) );
  OR2X2 U193 ( .A(A[11]), .B(B[11]), .Y(n196) );
  NAND2X1 U194 ( .A(B[10]), .B(A[10]), .Y(n206) );
  OR2X2 U195 ( .A(A[7]), .B(B[7]), .Y(n212) );
  OR2X2 U196 ( .A(A[12]), .B(B[12]), .Y(n176) );
  NOR2X1 U197 ( .A(A[5]), .B(B[5]), .Y(n8) );
  NOR2X1 U198 ( .A(A[4]), .B(B[4]), .Y(n9) );
  NAND2X1 U199 ( .A(B[4]), .B(A[4]), .Y(n34) );
  NAND2X1 U200 ( .A(B[8]), .B(A[8]), .Y(n17) );
  NAND2X1 U201 ( .A(B[5]), .B(A[5]), .Y(n30) );
  NAND2X1 U202 ( .A(B[6]), .B(A[6]), .Y(n25) );
  NAND2X1 U203 ( .A(B[2]), .B(A[2]), .Y(n41) );
  OR2X2 U204 ( .A(A[6]), .B(B[6]), .Y(n28) );
  NOR2X1 U205 ( .A(A[3]), .B(B[3]), .Y(n10) );
  OR2X2 U206 ( .A(A[8]), .B(B[8]), .Y(n202) );
  OR2X2 U207 ( .A(A[1]), .B(B[1]), .Y(n63) );
  NAND2X1 U208 ( .A(B[1]), .B(A[1]), .Y(n65) );
  NAND2X1 U209 ( .A(B[0]), .B(A[0]), .Y(n145) );
  NOR2X1 U210 ( .A(A[0]), .B(B[0]), .Y(n11) );
  XOR2X1 U211 ( .A(n60), .B(n69), .Y(SUM[28]) );
  NOR2BX1 U212 ( .AN(n59), .B(n57), .Y(n69) );
  XOR2X1 U213 ( .A(n93), .B(n94), .Y(SUM[25]) );
  XOR2X1 U214 ( .A(n89), .B(n90), .Y(SUM[26]) );
  NOR2BXL U215 ( .AN(n88), .B(n82), .Y(n90) );
  NOR2BXL U216 ( .AN(n76), .B(n81), .Y(n86) );
  XOR2X1 U217 ( .A(n118), .B(n119), .Y(SUM[22]) );
  XOR2X1 U218 ( .A(n115), .B(n116), .Y(SUM[23]) );
  XOR2X1 U219 ( .A(n96), .B(n98), .Y(SUM[24]) );
  NOR2BX1 U220 ( .AN(n95), .B(n99), .Y(n98) );
  XOR2X1 U221 ( .A(n36), .B(n37), .Y(SUM[3]) );
  NOR2BX1 U222 ( .AN(n145), .B(n11), .Y(SUM[0]) );
  XOR2X1 U223 ( .A(n64), .B(n143), .Y(SUM[1]) );
  XOR2X1 U224 ( .A(n42), .B(n61), .Y(SUM[2]) );
  XOR2X1 U225 ( .A(n173), .B(n35), .Y(SUM[4]) );
  XOR2X1 U226 ( .A(n31), .B(n32), .Y(SUM[5]) );
  XOR2X1 U227 ( .A(n26), .B(n27), .Y(SUM[6]) );
  XOR2X1 U228 ( .A(n19), .B(n20), .Y(SUM[7]) );
  XOR2X1 U229 ( .A(n15), .B(n16), .Y(SUM[8]) );
  XOR2X1 U230 ( .A(n12), .B(n13), .Y(SUM[9]) );
  XOR2X1 U231 ( .A(n205), .B(n207), .Y(SUM[10]) );
  XOR2X1 U232 ( .A(n203), .B(n204), .Y(SUM[11]) );
  XOR2X1 U233 ( .A(n189), .B(n190), .Y(SUM[12]) );
  XOR2X1 U234 ( .A(n185), .B(n186), .Y(SUM[13]) );
  XOR2X1 U235 ( .A(n182), .B(n183), .Y(SUM[14]) );
  XOR2X1 U236 ( .A(n179), .B(n180), .Y(SUM[15]) );
  XOR2X1 U237 ( .A(n130), .B(n155), .Y(SUM[16]) );
  XOR2X1 U238 ( .A(n152), .B(n153), .Y(SUM[17]) );
  XOR2X1 U239 ( .A(n149), .B(n150), .Y(SUM[18]) );
  XOR2X1 U240 ( .A(n146), .B(n147), .Y(SUM[19]) );
  XOR2X1 U241 ( .A(n123), .B(n125), .Y(SUM[20]) );
  NOR2BX1 U242 ( .AN(n108), .B(n126), .Y(n125) );
  XOR2X1 U243 ( .A(n121), .B(n122), .Y(SUM[21]) );
  NOR2X4 U244 ( .A(B[30]), .B(A[30]), .Y(n48) );
  OR2X4 U245 ( .A(A[29]), .B(B[29]), .Y(n52) );
  CLKINVX3 U246 ( .A(n68), .Y(n57) );
  CLKINVX3 U247 ( .A(n84), .Y(n81) );
  OR2X4 U248 ( .A(A[27]), .B(B[27]), .Y(n84) );
  CLKINVX3 U249 ( .A(n83), .Y(n82) );
  OR2X4 U250 ( .A(A[26]), .B(B[26]), .Y(n83) );
endmodule


module message_schedule ( clk, reset, data, write_enable, inner_busy, Wt );
  input [31:0] data;
  output [31:0] Wt;
  input clk, reset, write_enable, inner_busy;
  wire   n647, N622, N623, N624, N625, N626, N627, N628, n578, n613, n614,
         n615, N9, N8, N7, N67, N66, N65, N64, N63, N62, N61, N60, N6, N59,
         N58, N57, N56, N55, N54, N53, N52, N51, N50, N5, N49, N48, N47, N46,
         N45, N44, N43, N42, N41, N40, N4, N39, N38, N37, N36, N35, N34, N33,
         N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, n14, n17, n21, n23, n24,
         n377, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643;
  wire   [31:0] R14;
  wire   [31:0] sigma0;
  wire   [31:0] R1;
  wire   [31:0] sigma1;
  wire   [31:0] R15;
  wire   [31:0] R6;
  wire   [31:0] logic_result;
  wire   [6:0] counter;
  wire   [31:0] R2;
  wire   [31:0] R3;
  wire   [31:0] R4;
  wire   [31:0] R5;
  wire   [31:0] R7;
  wire   [31:0] R8;
  wire   [31:0] R9;
  wire   [31:0] R10;
  wire   [31:0] R11;
  wire   [31:0] R12;
  wire   [31:0] R13;

  DFFHQX4 Wt_reg_15_ ( .D(n627), .CK(clk), .Q(Wt[15]) );
  DFFHQX4 Wt_reg_14_ ( .D(n628), .CK(clk), .Q(Wt[14]) );
  DFFHQX4 Wt_reg_13_ ( .D(n629), .CK(clk), .Q(Wt[13]) );
  DFFHQX4 Wt_reg_12_ ( .D(n630), .CK(clk), .Q(Wt[12]) );
  DFFHQX4 Wt_reg_11_ ( .D(n631), .CK(clk), .Q(Wt[11]) );
  DFFHQX4 Wt_reg_10_ ( .D(n632), .CK(clk), .Q(Wt[10]) );
  DFFHQX4 Wt_reg_9_ ( .D(n633), .CK(clk), .Q(Wt[9]) );
  DFFHQX4 Wt_reg_8_ ( .D(n634), .CK(clk), .Q(Wt[8]) );
  DFFHQX4 Wt_reg_7_ ( .D(n635), .CK(clk), .Q(Wt[7]) );
  DFFHQX4 Wt_reg_6_ ( .D(n636), .CK(clk), .Q(Wt[6]) );
  DFFHQX4 Wt_reg_5_ ( .D(n637), .CK(clk), .Q(Wt[5]) );
  DFFHQX4 Wt_reg_4_ ( .D(n638), .CK(clk), .Q(Wt[4]) );
  DFFHQX4 Wt_reg_3_ ( .D(n639), .CK(clk), .Q(Wt[3]) );
  DFFHQX4 Wt_reg_2_ ( .D(n640), .CK(clk), .Q(Wt[2]) );
  DFFTRX4 R6_reg_1_ ( .D(R5[1]), .RN(n503), .CK(clk), .Q(R6[1]) );
  DFFTRX4 R15_reg_1_ ( .D(R14[1]), .RN(n502), .CK(clk), .Q(R15[1]) );
  DFFHQX4 Wt_reg_0_ ( .D(n642), .CK(clk), .Q(n647) );
  DFFTRX4 R6_reg_0_ ( .D(R5[0]), .RN(n501), .CK(clk), .Q(R6[0]) );
  DFFTRX4 R15_reg_0_ ( .D(R14[0]), .RN(n501), .CK(clk), .Q(R15[0]) );
  message_schedule_DW01_inc_0 add_110 ( .A(counter), .SUM({N628, N627, N626, 
        N625, N624, N623, N622}) );
  message_schedule_DW01_add_2 add_2_root_add_0_root_add_34_3 ( .A(R15), .B(R6), 
        .SUM({N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, 
        N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, 
        N40, N39, N38, N37, N36}) );
  message_schedule_DW01_add_4 add_1_root_add_0_root_add_34_3 ( .A(sigma1), .B(
        sigma0), .SUM({N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4}) );
  message_schedule_DW01_add_5 add_0_root_add_0_root_add_34_3 ( .A({N67, N66, 
        N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, 
        N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, 
        N37, N36}), .B({N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4}), .SUM(logic_result) );
  DFFTRX1 R15_reg_31_ ( .D(R14[31]), .RN(n539), .CK(clk), .Q(R15[31]) );
  DFFTRX1 R15_reg_29_ ( .D(R14[29]), .RN(n537), .CK(clk), .Q(R15[29]) );
  DFFTRX1 R15_reg_30_ ( .D(R14[30]), .RN(n538), .CK(clk), .Q(R15[30]) );
  DFFTRX1 counter_reg_6_ ( .D(N628), .RN(n539), .CK(clk), .Q(counter[6]) );
  DFFTRX1 R6_reg_31_ ( .D(R5[31]), .RN(n540), .CK(clk), .Q(R6[31]) );
  DFFTRX1 R6_reg_29_ ( .D(R5[29]), .RN(n538), .CK(clk), .Q(R6[29]) );
  DFFTRX1 R6_reg_30_ ( .D(R5[30]), .RN(n539), .CK(clk), .Q(R6[30]) );
  DFFTRX1 counter_reg_1_ ( .D(N623), .RN(n536), .CK(clk), .Q(counter[1]) );
  DFFTRX1 counter_reg_0_ ( .D(N622), .RN(n537), .CK(clk), .Q(counter[0]) );
  DFFTRX1 R15_reg_28_ ( .D(R14[28]), .RN(n536), .CK(clk), .Q(R15[28]) );
  DFFTRX1 R15_reg_27_ ( .D(R14[27]), .RN(n534), .CK(clk), .Q(R15[27]) );
  DFFTRX1 R15_reg_26_ ( .D(R14[26]), .RN(n533), .CK(clk), .Q(R15[26]) );
  DFFTRX1 R6_reg_28_ ( .D(R5[28]), .RN(n536), .CK(clk), .Q(R6[28]) );
  DFFTRX1 R6_reg_27_ ( .D(R5[27]), .RN(n535), .CK(clk), .Q(R6[27]) );
  DFFTRX1 R6_reg_26_ ( .D(R5[26]), .RN(n534), .CK(clk), .Q(R6[26]) );
  DFFTRX1 counter_reg_5_ ( .D(N627), .RN(n540), .CK(clk), .Q(counter[5]) );
  DFFTRX1 counter_reg_3_ ( .D(N625), .RN(n540), .CK(clk), .Q(counter[3]) );
  DFFTRX1 counter_reg_4_ ( .D(N626), .RN(n539), .CK(clk), .Q(counter[4]) );
  DFFTRX1 counter_reg_2_ ( .D(N624), .RN(n538), .CK(clk), .Q(counter[2]) );
  DFFTRX1 R15_reg_25_ ( .D(R14[25]), .RN(n532), .CK(clk), .Q(R15[25]) );
  DFFTRX1 R15_reg_24_ ( .D(R14[24]), .RN(n531), .CK(clk), .Q(R15[24]) );
  DFFTRX1 R15_reg_23_ ( .D(R14[23]), .RN(n529), .CK(clk), .Q(R15[23]) );
  DFFTRX1 R15_reg_22_ ( .D(R14[22]), .RN(n528), .CK(clk), .Q(R15[22]) );
  DFFTRX1 R6_reg_25_ ( .D(R5[25]), .RN(n533), .CK(clk), .Q(R6[25]) );
  DFFTRX1 R6_reg_24_ ( .D(R5[24]), .RN(n531), .CK(clk), .Q(R6[24]) );
  DFFTRX1 R6_reg_23_ ( .D(R5[23]), .RN(n530), .CK(clk), .Q(R6[23]) );
  DFFTRX1 R6_reg_22_ ( .D(R5[22]), .RN(n529), .CK(clk), .Q(R6[22]) );
  DFFTRX1 R6_reg_21_ ( .D(R5[21]), .RN(n528), .CK(clk), .Q(R6[21]) );
  DFFHQXL Wt_reg_31_ ( .D(n608), .CK(clk), .Q(Wt[31]) );
  DFFTRX1 R15_reg_21_ ( .D(R14[21]), .RN(n527), .CK(clk), .Q(R15[21]) );
  DFFTRX1 R15_reg_20_ ( .D(R14[20]), .RN(n526), .CK(clk), .Q(R15[20]) );
  DFFTRX1 R15_reg_19_ ( .D(R14[19]), .RN(n524), .CK(clk), .Q(R15[19]) );
  DFFTRX1 R15_reg_18_ ( .D(R14[18]), .RN(n523), .CK(clk), .Q(R15[18]) );
  DFFTRX1 R6_reg_20_ ( .D(R5[20]), .RN(n526), .CK(clk), .Q(R6[20]) );
  DFFTRX1 R6_reg_19_ ( .D(R5[19]), .RN(n525), .CK(clk), .Q(R6[19]) );
  DFFTRX1 R6_reg_18_ ( .D(R5[18]), .RN(n524), .CK(clk), .Q(R6[18]) );
  DFFTRX1 R14_reg_2_ ( .D(R13[2]), .RN(n503), .CK(clk), .Q(R14[2]) );
  DFFTRX1 R1_reg_9_ ( .D(Wt[9]), .RN(n513), .CK(clk), .Q(R1[9]) );
  DFFTRX1 R1_reg_6_ ( .D(Wt[6]), .RN(n509), .CK(clk), .Q(R1[6]) );
  DFFTRX1 R1_reg_5_ ( .D(Wt[5]), .RN(n508), .CK(clk), .Q(R1[5]) );
  DFFTRX1 R1_reg_8_ ( .D(Wt[8]), .RN(n512), .CK(clk), .Q(R1[8]) );
  DFFTRX1 R1_reg_7_ ( .D(Wt[7]), .RN(n510), .CK(clk), .Q(R1[7]) );
  DFFHQXL Wt_reg_30_ ( .D(n609), .CK(clk), .Q(Wt[30]) );
  DFFHQX1 Wt_reg_29_ ( .D(n610), .CK(clk), .Q(Wt[29]) );
  DFFTRX1 R15_reg_17_ ( .D(R14[17]), .RN(n522), .CK(clk), .Q(R15[17]) );
  DFFTRX1 R15_reg_16_ ( .D(R14[16]), .RN(n521), .CK(clk), .Q(R15[16]) );
  DFFTRX1 R15_reg_15_ ( .D(R14[15]), .RN(n519), .CK(clk), .Q(R15[15]) );
  DFFTRX1 R15_reg_14_ ( .D(R14[14]), .RN(n518), .CK(clk), .Q(R15[14]) );
  DFFTRX1 R6_reg_17_ ( .D(R5[17]), .RN(n523), .CK(clk), .Q(R6[17]) );
  DFFTRX1 R6_reg_16_ ( .D(R5[16]), .RN(n521), .CK(clk), .Q(R6[16]) );
  DFFTRX1 R6_reg_15_ ( .D(R5[15]), .RN(n520), .CK(clk), .Q(R6[15]) );
  DFFTRX1 R6_reg_14_ ( .D(R5[14]), .RN(n519), .CK(clk), .Q(R6[14]) );
  DFFTRX1 R14_reg_1_ ( .D(R13[1]), .RN(n502), .CK(clk), .Q(R14[1]) );
  DFFTRX1 R14_reg_0_ ( .D(R13[0]), .RN(n501), .CK(clk), .Q(R14[0]) );
  DFFTRX1 R1_reg_4_ ( .D(Wt[4]), .RN(n507), .CK(clk), .Q(R1[4]) );
  DFFHQX1 Wt_reg_28_ ( .D(n611), .CK(clk), .Q(Wt[28]) );
  DFFTRX1 R1_reg_29_ ( .D(Wt[29]), .RN(n538), .CK(clk), .Q(R1[29]) );
  DFFTRX1 R1_reg_27_ ( .D(Wt[27]), .RN(n535), .CK(clk), .Q(R1[27]) );
  DFFTRX1 R14_reg_26_ ( .D(R13[26]), .RN(n533), .CK(clk), .Q(R14[26]) );
  DFFTRX1 R1_reg_31_ ( .D(Wt[31]), .RN(n540), .CK(clk), .Q(R1[31]) );
  DFFTRX1 R1_reg_30_ ( .D(Wt[30]), .RN(n539), .CK(clk), .Q(R1[30]) );
  DFFTRX1 R14_reg_28_ ( .D(R13[28]), .RN(n536), .CK(clk), .Q(R14[28]) );
  DFFTRX1 R14_reg_15_ ( .D(R13[15]), .RN(n519), .CK(clk), .Q(R14[15]) );
  DFFTRX1 R14_reg_17_ ( .D(R13[17]), .RN(n522), .CK(clk), .Q(R14[17]) );
  DFFTRX1 R14_reg_31_ ( .D(R13[31]), .RN(n539), .CK(clk), .Q(R14[31]) );
  DFFTRX1 R14_reg_30_ ( .D(R13[30]), .RN(n538), .CK(clk), .Q(R14[30]) );
  DFFTRX1 R14_reg_29_ ( .D(R13[29]), .RN(n537), .CK(clk), .Q(R14[29]) );
  DFFTRX1 R1_reg_0_ ( .D(Wt[0]), .RN(n502), .CK(clk), .Q(R1[0]) );
  DFFTRX1 R1_reg_3_ ( .D(Wt[3]), .RN(n505), .CK(clk), .Q(R1[3]) );
  DFFTRX1 R1_reg_2_ ( .D(Wt[2]), .RN(n504), .CK(clk), .Q(R1[2]) );
  DFFTRX1 R15_reg_13_ ( .D(R14[13]), .RN(n517), .CK(clk), .Q(R15[13]) );
  DFFTRX1 R15_reg_12_ ( .D(R14[12]), .RN(n516), .CK(clk), .Q(R15[12]) );
  DFFTRX1 R15_reg_11_ ( .D(R14[11]), .RN(n514), .CK(clk), .Q(R15[11]) );
  DFFTRX1 R15_reg_10_ ( .D(R14[10]), .RN(n513), .CK(clk), .Q(R15[10]) );
  DFFTRX1 R6_reg_13_ ( .D(R5[13]), .RN(n518), .CK(clk), .Q(R6[13]) );
  DFFTRX1 R6_reg_12_ ( .D(R5[12]), .RN(n516), .CK(clk), .Q(R6[12]) );
  DFFTRX1 R6_reg_11_ ( .D(R5[11]), .RN(n515), .CK(clk), .Q(R6[11]) );
  DFFTRX1 R6_reg_10_ ( .D(R5[10]), .RN(n514), .CK(clk), .Q(R6[10]) );
  DFFTRX1 R14_reg_19_ ( .D(R13[19]), .RN(n524), .CK(clk), .Q(R14[19]) );
  DFFTRX1 R14_reg_18_ ( .D(R13[18]), .RN(n523), .CK(clk), .Q(R14[18]) );
  DFFTRX1 R1_reg_19_ ( .D(Wt[19]), .RN(n525), .CK(clk), .Q(R1[19]) );
  DFFTRX1 R14_reg_3_ ( .D(R13[3]), .RN(n504), .CK(clk), .Q(R14[3]) );
  DFFTRX1 R14_reg_6_ ( .D(R13[6]), .RN(n508), .CK(clk), .Q(R14[6]) );
  DFFTRX1 R14_reg_5_ ( .D(R13[5]), .RN(n507), .CK(clk), .Q(R14[5]) );
  DFFTRX1 R14_reg_4_ ( .D(R13[4]), .RN(n506), .CK(clk), .Q(R14[4]) );
  DFFTRX1 R1_reg_28_ ( .D(Wt[28]), .RN(n537), .CK(clk), .Q(R1[28]) );
  DFFTRX1 R14_reg_27_ ( .D(R13[27]), .RN(n534), .CK(clk), .Q(R14[27]) );
  DFFTRX1 R1_reg_26_ ( .D(Wt[26]), .RN(n534), .CK(clk), .Q(R1[26]) );
  DFFTRX1 R1_reg_25_ ( .D(Wt[25]), .RN(n533), .CK(clk), .Q(R1[25]) );
  DFFTRX1 R14_reg_25_ ( .D(R13[25]), .RN(n532), .CK(clk), .Q(R14[25]) );
  DFFTRX1 R1_reg_24_ ( .D(Wt[24]), .RN(n532), .CK(clk), .Q(R1[24]) );
  DFFTRX1 R14_reg_24_ ( .D(R13[24]), .RN(n531), .CK(clk), .Q(R14[24]) );
  DFFTRX1 R1_reg_22_ ( .D(Wt[22]), .RN(n529), .CK(clk), .Q(R1[22]) );
  DFFTRX1 R14_reg_14_ ( .D(R13[14]), .RN(n518), .CK(clk), .Q(R14[14]) );
  DFFTRX1 R14_reg_13_ ( .D(R13[13]), .RN(n517), .CK(clk), .Q(R14[13]) );
  DFFTRX1 R1_reg_16_ ( .D(Wt[16]), .RN(n522), .CK(clk), .Q(R1[16]) );
  DFFTRX1 R1_reg_15_ ( .D(Wt[15]), .RN(n520), .CK(clk), .Q(R1[15]) );
  DFFTRX1 R1_reg_14_ ( .D(Wt[14]), .RN(n519), .CK(clk), .Q(R1[14]) );
  DFFTRX1 R1_reg_13_ ( .D(Wt[13]), .RN(n518), .CK(clk), .Q(R1[13]) );
  DFFTRX1 R1_reg_12_ ( .D(Wt[12]), .RN(n517), .CK(clk), .Q(R1[12]) );
  DFFTRX1 R1_reg_11_ ( .D(Wt[11]), .RN(n515), .CK(clk), .Q(R1[11]) );
  DFFTRX1 R1_reg_10_ ( .D(Wt[10]), .RN(n514), .CK(clk), .Q(R1[10]) );
  DFFTRX1 R14_reg_10_ ( .D(R13[10]), .RN(n513), .CK(clk), .Q(R14[10]) );
  DFFTRX1 R14_reg_9_ ( .D(R13[9]), .RN(n512), .CK(clk), .Q(R14[9]) );
  DFFTRX1 R14_reg_8_ ( .D(R13[8]), .RN(n511), .CK(clk), .Q(R14[8]) );
  DFFTRX1 R14_reg_7_ ( .D(R13[7]), .RN(n509), .CK(clk), .Q(R14[7]) );
  DFFTRX1 R14_reg_16_ ( .D(R13[16]), .RN(n521), .CK(clk), .Q(R14[16]) );
  DFFTRX1 R15_reg_9_ ( .D(R14[9]), .RN(n512), .CK(clk), .Q(R15[9]) );
  DFFTRX1 R15_reg_8_ ( .D(R14[8]), .RN(n511), .CK(clk), .Q(R15[8]) );
  DFFTRX1 R15_reg_7_ ( .D(R14[7]), .RN(n509), .CK(clk), .Q(R15[7]) );
  DFFTRX1 R15_reg_6_ ( .D(R14[6]), .RN(n508), .CK(clk), .Q(R15[6]) );
  DFFTRX1 R6_reg_9_ ( .D(R5[9]), .RN(n513), .CK(clk), .Q(R6[9]) );
  DFFTRX1 R6_reg_8_ ( .D(R5[8]), .RN(n511), .CK(clk), .Q(R6[8]) );
  DFFTRX1 R6_reg_7_ ( .D(R5[7]), .RN(n510), .CK(clk), .Q(R6[7]) );
  DFFTRX1 R6_reg_6_ ( .D(R5[6]), .RN(n509), .CK(clk), .Q(R6[6]) );
  DFFHQX1 Wt_reg_22_ ( .D(n620), .CK(clk), .Q(Wt[22]) );
  DFFTRX1 R15_reg_5_ ( .D(R14[5]), .RN(n507), .CK(clk), .Q(R15[5]) );
  DFFTRX1 R15_reg_4_ ( .D(R14[4]), .RN(n506), .CK(clk), .Q(R15[4]) );
  DFFTRX1 R15_reg_3_ ( .D(R14[3]), .RN(n504), .CK(clk), .Q(R15[3]) );
  DFFTRX1 R6_reg_5_ ( .D(R5[5]), .RN(n508), .CK(clk), .Q(R6[5]) );
  DFFTRX1 R6_reg_4_ ( .D(R5[4]), .RN(n506), .CK(clk), .Q(R6[4]) );
  DFFTRX1 R6_reg_3_ ( .D(R5[3]), .RN(n505), .CK(clk), .Q(R6[3]) );
  DFFHQX1 Wt_reg_19_ ( .D(n623), .CK(clk), .Q(Wt[19]) );
  DFFHQX1 Wt_reg_16_ ( .D(n626), .CK(clk), .Q(Wt[16]) );
  DFFTRX1 R2_reg_31_ ( .D(R1[31]), .RN(n540), .CK(clk), .Q(R2[31]) );
  DFFTRX1 R3_reg_31_ ( .D(R2[31]), .RN(n540), .CK(clk), .Q(R3[31]) );
  DFFTRX1 R4_reg_31_ ( .D(R3[31]), .RN(n540), .CK(clk), .Q(R4[31]) );
  DFFTRX1 R5_reg_31_ ( .D(R4[31]), .RN(n540), .CK(clk), .Q(R5[31]) );
  DFFTRX1 R7_reg_31_ ( .D(R6[31]), .RN(n540), .CK(clk), .Q(R7[31]) );
  DFFTRX1 R8_reg_31_ ( .D(R7[31]), .RN(n540), .CK(clk), .Q(R8[31]) );
  DFFTRX1 R9_reg_31_ ( .D(R8[31]), .RN(n540), .CK(clk), .Q(R9[31]) );
  DFFTRX1 R10_reg_31_ ( .D(R9[31]), .RN(n540), .CK(clk), .Q(R10[31]) );
  DFFTRX1 R11_reg_31_ ( .D(R10[31]), .RN(n540), .CK(clk), .Q(R11[31]) );
  DFFTRX1 R12_reg_31_ ( .D(R11[31]), .RN(n540), .CK(clk), .Q(R12[31]) );
  DFFTRX1 R13_reg_31_ ( .D(R12[31]), .RN(n539), .CK(clk), .Q(R13[31]) );
  DFFTRX1 R2_reg_30_ ( .D(R1[30]), .RN(n539), .CK(clk), .Q(R2[30]) );
  DFFTRX1 R3_reg_30_ ( .D(R2[30]), .RN(n539), .CK(clk), .Q(R3[30]) );
  DFFTRX1 R4_reg_30_ ( .D(R3[30]), .RN(n539), .CK(clk), .Q(R4[30]) );
  DFFTRX1 R5_reg_30_ ( .D(R4[30]), .RN(n539), .CK(clk), .Q(R5[30]) );
  DFFTRX1 R7_reg_30_ ( .D(R6[30]), .RN(n539), .CK(clk), .Q(R7[30]) );
  DFFTRX1 R8_reg_30_ ( .D(R7[30]), .RN(n539), .CK(clk), .Q(R8[30]) );
  DFFTRX1 R9_reg_30_ ( .D(R8[30]), .RN(n539), .CK(clk), .Q(R9[30]) );
  DFFTRX1 R10_reg_30_ ( .D(R9[30]), .RN(n538), .CK(clk), .Q(R10[30]) );
  DFFTRX1 R11_reg_30_ ( .D(R10[30]), .RN(n538), .CK(clk), .Q(R11[30]) );
  DFFTRX1 R12_reg_30_ ( .D(R11[30]), .RN(n538), .CK(clk), .Q(R12[30]) );
  DFFTRX1 R13_reg_30_ ( .D(R12[30]), .RN(n538), .CK(clk), .Q(R13[30]) );
  DFFTRX1 R2_reg_29_ ( .D(R1[29]), .RN(n538), .CK(clk), .Q(R2[29]) );
  DFFTRX1 R3_reg_29_ ( .D(R2[29]), .RN(n538), .CK(clk), .Q(R3[29]) );
  DFFTRX1 R4_reg_29_ ( .D(R3[29]), .RN(n538), .CK(clk), .Q(R4[29]) );
  DFFTRX1 R5_reg_29_ ( .D(R4[29]), .RN(n538), .CK(clk), .Q(R5[29]) );
  DFFTRX1 R7_reg_29_ ( .D(R6[29]), .RN(n537), .CK(clk), .Q(R7[29]) );
  DFFTRX1 R8_reg_29_ ( .D(R7[29]), .RN(n537), .CK(clk), .Q(R8[29]) );
  DFFTRX1 R9_reg_29_ ( .D(R8[29]), .RN(n537), .CK(clk), .Q(R9[29]) );
  DFFTRX1 R10_reg_29_ ( .D(R9[29]), .RN(n537), .CK(clk), .Q(R10[29]) );
  DFFTRX1 R11_reg_29_ ( .D(R10[29]), .RN(n537), .CK(clk), .Q(R11[29]) );
  DFFTRX1 R12_reg_29_ ( .D(R11[29]), .RN(n537), .CK(clk), .Q(R12[29]) );
  DFFTRX1 R13_reg_29_ ( .D(R12[29]), .RN(n537), .CK(clk), .Q(R13[29]) );
  DFFTRX1 R2_reg_28_ ( .D(R1[28]), .RN(n537), .CK(clk), .Q(R2[28]) );
  DFFTRX1 R3_reg_28_ ( .D(R2[28]), .RN(n537), .CK(clk), .Q(R3[28]) );
  DFFTRX1 R4_reg_28_ ( .D(R3[28]), .RN(n536), .CK(clk), .Q(R4[28]) );
  DFFTRX1 R5_reg_28_ ( .D(R4[28]), .RN(n536), .CK(clk), .Q(R5[28]) );
  DFFTRX1 R7_reg_28_ ( .D(R6[28]), .RN(n536), .CK(clk), .Q(R7[28]) );
  DFFTRX1 R8_reg_28_ ( .D(R7[28]), .RN(n536), .CK(clk), .Q(R8[28]) );
  DFFTRX1 R9_reg_28_ ( .D(R8[28]), .RN(n536), .CK(clk), .Q(R9[28]) );
  DFFTRX1 R10_reg_28_ ( .D(R9[28]), .RN(n536), .CK(clk), .Q(R10[28]) );
  DFFTRX1 R11_reg_28_ ( .D(R10[28]), .RN(n536), .CK(clk), .Q(R11[28]) );
  DFFTRX1 R12_reg_28_ ( .D(R11[28]), .RN(n536), .CK(clk), .Q(R12[28]) );
  DFFTRX1 R13_reg_28_ ( .D(R12[28]), .RN(n536), .CK(clk), .Q(R13[28]) );
  DFFTRX1 R4_reg_0_ ( .D(R3[0]), .RN(n501), .CK(clk), .Q(R4[0]) );
  DFFTRX1 R5_reg_0_ ( .D(R4[0]), .RN(n501), .CK(clk), .Q(R5[0]) );
  DFFTRX1 R8_reg_0_ ( .D(R7[0]), .RN(n501), .CK(clk), .Q(R8[0]) );
  DFFTRX1 R9_reg_0_ ( .D(R8[0]), .RN(n501), .CK(clk), .Q(R9[0]) );
  DFFTRX1 R10_reg_0_ ( .D(R9[0]), .RN(n501), .CK(clk), .Q(R10[0]) );
  DFFTRX1 R11_reg_0_ ( .D(R10[0]), .RN(n501), .CK(clk), .Q(R11[0]) );
  DFFTRX1 R12_reg_0_ ( .D(R11[0]), .RN(n501), .CK(clk), .Q(R12[0]) );
  DFFTRX1 R13_reg_0_ ( .D(R12[0]), .RN(n501), .CK(clk), .Q(R13[0]) );
  DFFTRX1 R2_reg_27_ ( .D(R1[27]), .RN(n535), .CK(clk), .Q(R2[27]) );
  DFFTRX1 R3_reg_27_ ( .D(R2[27]), .RN(n535), .CK(clk), .Q(R3[27]) );
  DFFTRX1 R4_reg_27_ ( .D(R3[27]), .RN(n535), .CK(clk), .Q(R4[27]) );
  DFFTRX1 R5_reg_27_ ( .D(R4[27]), .RN(n535), .CK(clk), .Q(R5[27]) );
  DFFTRX1 R7_reg_27_ ( .D(R6[27]), .RN(n535), .CK(clk), .Q(R7[27]) );
  DFFTRX1 R8_reg_27_ ( .D(R7[27]), .RN(n535), .CK(clk), .Q(R8[27]) );
  DFFTRX1 R9_reg_27_ ( .D(R8[27]), .RN(n535), .CK(clk), .Q(R9[27]) );
  DFFTRX1 R10_reg_27_ ( .D(R9[27]), .RN(n535), .CK(clk), .Q(R10[27]) );
  DFFTRX1 R11_reg_27_ ( .D(R10[27]), .RN(n535), .CK(clk), .Q(R11[27]) );
  DFFTRX1 R12_reg_27_ ( .D(R11[27]), .RN(n535), .CK(clk), .Q(R12[27]) );
  DFFTRX1 R13_reg_27_ ( .D(R12[27]), .RN(n534), .CK(clk), .Q(R13[27]) );
  DFFTRX1 R2_reg_26_ ( .D(R1[26]), .RN(n534), .CK(clk), .Q(R2[26]) );
  DFFTRX1 R3_reg_26_ ( .D(R2[26]), .RN(n534), .CK(clk), .Q(R3[26]) );
  DFFTRX1 R4_reg_26_ ( .D(R3[26]), .RN(n534), .CK(clk), .Q(R4[26]) );
  DFFTRX1 R5_reg_26_ ( .D(R4[26]), .RN(n534), .CK(clk), .Q(R5[26]) );
  DFFTRX1 R7_reg_26_ ( .D(R6[26]), .RN(n534), .CK(clk), .Q(R7[26]) );
  DFFTRX1 R8_reg_26_ ( .D(R7[26]), .RN(n534), .CK(clk), .Q(R8[26]) );
  DFFTRX1 R9_reg_26_ ( .D(R8[26]), .RN(n534), .CK(clk), .Q(R9[26]) );
  DFFTRX1 R10_reg_26_ ( .D(R9[26]), .RN(n533), .CK(clk), .Q(R10[26]) );
  DFFTRX1 R11_reg_26_ ( .D(R10[26]), .RN(n533), .CK(clk), .Q(R11[26]) );
  DFFTRX1 R12_reg_26_ ( .D(R11[26]), .RN(n533), .CK(clk), .Q(R12[26]) );
  DFFTRX1 R13_reg_26_ ( .D(R12[26]), .RN(n533), .CK(clk), .Q(R13[26]) );
  DFFTRX1 R2_reg_25_ ( .D(R1[25]), .RN(n533), .CK(clk), .Q(R2[25]) );
  DFFTRX1 R3_reg_25_ ( .D(R2[25]), .RN(n533), .CK(clk), .Q(R3[25]) );
  DFFTRX1 R4_reg_25_ ( .D(R3[25]), .RN(n533), .CK(clk), .Q(R4[25]) );
  DFFTRX1 R5_reg_25_ ( .D(R4[25]), .RN(n533), .CK(clk), .Q(R5[25]) );
  DFFTRX1 R7_reg_25_ ( .D(R6[25]), .RN(n532), .CK(clk), .Q(R7[25]) );
  DFFTRX1 R8_reg_25_ ( .D(R7[25]), .RN(n532), .CK(clk), .Q(R8[25]) );
  DFFTRX1 R9_reg_25_ ( .D(R8[25]), .RN(n532), .CK(clk), .Q(R9[25]) );
  DFFTRX1 R10_reg_25_ ( .D(R9[25]), .RN(n532), .CK(clk), .Q(R10[25]) );
  DFFTRX1 R11_reg_25_ ( .D(R10[25]), .RN(n532), .CK(clk), .Q(R11[25]) );
  DFFTRX1 R12_reg_25_ ( .D(R11[25]), .RN(n532), .CK(clk), .Q(R12[25]) );
  DFFTRX1 R13_reg_25_ ( .D(R12[25]), .RN(n532), .CK(clk), .Q(R13[25]) );
  DFFTRX1 R2_reg_24_ ( .D(R1[24]), .RN(n532), .CK(clk), .Q(R2[24]) );
  DFFTRX1 R3_reg_24_ ( .D(R2[24]), .RN(n532), .CK(clk), .Q(R3[24]) );
  DFFTRX1 R4_reg_24_ ( .D(R3[24]), .RN(n531), .CK(clk), .Q(R4[24]) );
  DFFTRX1 R5_reg_24_ ( .D(R4[24]), .RN(n531), .CK(clk), .Q(R5[24]) );
  DFFTRX1 R7_reg_24_ ( .D(R6[24]), .RN(n531), .CK(clk), .Q(R7[24]) );
  DFFTRX1 R8_reg_24_ ( .D(R7[24]), .RN(n531), .CK(clk), .Q(R8[24]) );
  DFFTRX1 R9_reg_24_ ( .D(R8[24]), .RN(n531), .CK(clk), .Q(R9[24]) );
  DFFTRX1 R10_reg_24_ ( .D(R9[24]), .RN(n531), .CK(clk), .Q(R10[24]) );
  DFFTRX1 R11_reg_24_ ( .D(R10[24]), .RN(n531), .CK(clk), .Q(R11[24]) );
  DFFTRX1 R12_reg_24_ ( .D(R11[24]), .RN(n531), .CK(clk), .Q(R12[24]) );
  DFFTRX1 R13_reg_24_ ( .D(R12[24]), .RN(n531), .CK(clk), .Q(R13[24]) );
  DFFTRX1 R2_reg_23_ ( .D(R1[23]), .RN(n530), .CK(clk), .Q(R2[23]) );
  DFFTRX1 R3_reg_23_ ( .D(R2[23]), .RN(n530), .CK(clk), .Q(R3[23]) );
  DFFTRX1 R4_reg_23_ ( .D(R3[23]), .RN(n530), .CK(clk), .Q(R4[23]) );
  DFFTRX1 R5_reg_23_ ( .D(R4[23]), .RN(n530), .CK(clk), .Q(R5[23]) );
  DFFTRX1 R7_reg_23_ ( .D(R6[23]), .RN(n530), .CK(clk), .Q(R7[23]) );
  DFFTRX1 R8_reg_23_ ( .D(R7[23]), .RN(n530), .CK(clk), .Q(R8[23]) );
  DFFTRX1 R9_reg_23_ ( .D(R8[23]), .RN(n530), .CK(clk), .Q(R9[23]) );
  DFFTRX1 R10_reg_23_ ( .D(R9[23]), .RN(n530), .CK(clk), .Q(R10[23]) );
  DFFTRX1 R11_reg_23_ ( .D(R10[23]), .RN(n530), .CK(clk), .Q(R11[23]) );
  DFFTRX1 R12_reg_23_ ( .D(R11[23]), .RN(n530), .CK(clk), .Q(R12[23]) );
  DFFTRX1 R13_reg_23_ ( .D(R12[23]), .RN(n529), .CK(clk), .Q(R13[23]) );
  DFFTRX1 R2_reg_22_ ( .D(R1[22]), .RN(n529), .CK(clk), .Q(R2[22]) );
  DFFTRX1 R3_reg_22_ ( .D(R2[22]), .RN(n529), .CK(clk), .Q(R3[22]) );
  DFFTRX1 R4_reg_22_ ( .D(R3[22]), .RN(n529), .CK(clk), .Q(R4[22]) );
  DFFTRX1 R5_reg_22_ ( .D(R4[22]), .RN(n529), .CK(clk), .Q(R5[22]) );
  DFFTRX1 R7_reg_22_ ( .D(R6[22]), .RN(n529), .CK(clk), .Q(R7[22]) );
  DFFTRX1 R8_reg_22_ ( .D(R7[22]), .RN(n529), .CK(clk), .Q(R8[22]) );
  DFFTRX1 R9_reg_22_ ( .D(R8[22]), .RN(n529), .CK(clk), .Q(R9[22]) );
  DFFTRX1 R10_reg_22_ ( .D(R9[22]), .RN(n528), .CK(clk), .Q(R10[22]) );
  DFFTRX1 R11_reg_22_ ( .D(R10[22]), .RN(n528), .CK(clk), .Q(R11[22]) );
  DFFTRX1 R12_reg_22_ ( .D(R11[22]), .RN(n528), .CK(clk), .Q(R12[22]) );
  DFFTRX1 R13_reg_22_ ( .D(R12[22]), .RN(n528), .CK(clk), .Q(R13[22]) );
  DFFTRX1 R2_reg_21_ ( .D(R1[21]), .RN(n528), .CK(clk), .Q(R2[21]) );
  DFFTRX1 R3_reg_21_ ( .D(R2[21]), .RN(n528), .CK(clk), .Q(R3[21]) );
  DFFTRX1 R4_reg_21_ ( .D(R3[21]), .RN(n528), .CK(clk), .Q(R4[21]) );
  DFFTRX1 R5_reg_21_ ( .D(R4[21]), .RN(n528), .CK(clk), .Q(R5[21]) );
  DFFTRX1 R7_reg_21_ ( .D(R6[21]), .RN(n527), .CK(clk), .Q(R7[21]) );
  DFFTRX1 R8_reg_21_ ( .D(R7[21]), .RN(n527), .CK(clk), .Q(R8[21]) );
  DFFTRX1 R9_reg_21_ ( .D(R8[21]), .RN(n527), .CK(clk), .Q(R9[21]) );
  DFFTRX1 R10_reg_21_ ( .D(R9[21]), .RN(n527), .CK(clk), .Q(R10[21]) );
  DFFTRX1 R11_reg_21_ ( .D(R10[21]), .RN(n527), .CK(clk), .Q(R11[21]) );
  DFFTRX1 R12_reg_21_ ( .D(R11[21]), .RN(n527), .CK(clk), .Q(R12[21]) );
  DFFTRX1 R13_reg_21_ ( .D(R12[21]), .RN(n527), .CK(clk), .Q(R13[21]) );
  DFFTRX1 R2_reg_20_ ( .D(R1[20]), .RN(n527), .CK(clk), .Q(R2[20]) );
  DFFTRX1 R3_reg_20_ ( .D(R2[20]), .RN(n527), .CK(clk), .Q(R3[20]) );
  DFFTRX1 R4_reg_20_ ( .D(R3[20]), .RN(n526), .CK(clk), .Q(R4[20]) );
  DFFTRX1 R5_reg_20_ ( .D(R4[20]), .RN(n526), .CK(clk), .Q(R5[20]) );
  DFFTRX1 R7_reg_20_ ( .D(R6[20]), .RN(n526), .CK(clk), .Q(R7[20]) );
  DFFTRX1 R8_reg_20_ ( .D(R7[20]), .RN(n526), .CK(clk), .Q(R8[20]) );
  DFFTRX1 R9_reg_20_ ( .D(R8[20]), .RN(n526), .CK(clk), .Q(R9[20]) );
  DFFTRX1 R10_reg_20_ ( .D(R9[20]), .RN(n526), .CK(clk), .Q(R10[20]) );
  DFFTRX1 R11_reg_20_ ( .D(R10[20]), .RN(n526), .CK(clk), .Q(R11[20]) );
  DFFTRX1 R12_reg_20_ ( .D(R11[20]), .RN(n526), .CK(clk), .Q(R12[20]) );
  DFFTRX1 R13_reg_20_ ( .D(R12[20]), .RN(n526), .CK(clk), .Q(R13[20]) );
  DFFTRX1 R2_reg_19_ ( .D(R1[19]), .RN(n525), .CK(clk), .Q(R2[19]) );
  DFFTRX1 R3_reg_19_ ( .D(R2[19]), .RN(n525), .CK(clk), .Q(R3[19]) );
  DFFTRX1 R4_reg_19_ ( .D(R3[19]), .RN(n525), .CK(clk), .Q(R4[19]) );
  DFFTRX1 R5_reg_19_ ( .D(R4[19]), .RN(n525), .CK(clk), .Q(R5[19]) );
  DFFTRX1 R7_reg_19_ ( .D(R6[19]), .RN(n525), .CK(clk), .Q(R7[19]) );
  DFFTRX1 R8_reg_19_ ( .D(R7[19]), .RN(n525), .CK(clk), .Q(R8[19]) );
  DFFTRX1 R9_reg_19_ ( .D(R8[19]), .RN(n525), .CK(clk), .Q(R9[19]) );
  DFFTRX1 R10_reg_19_ ( .D(R9[19]), .RN(n525), .CK(clk), .Q(R10[19]) );
  DFFTRX1 R11_reg_19_ ( .D(R10[19]), .RN(n525), .CK(clk), .Q(R11[19]) );
  DFFTRX1 R12_reg_19_ ( .D(R11[19]), .RN(n525), .CK(clk), .Q(R12[19]) );
  DFFTRX1 R13_reg_19_ ( .D(R12[19]), .RN(n524), .CK(clk), .Q(R13[19]) );
  DFFTRX1 R2_reg_18_ ( .D(R1[18]), .RN(n524), .CK(clk), .Q(R2[18]) );
  DFFTRX1 R3_reg_18_ ( .D(R2[18]), .RN(n524), .CK(clk), .Q(R3[18]) );
  DFFTRX1 R4_reg_18_ ( .D(R3[18]), .RN(n524), .CK(clk), .Q(R4[18]) );
  DFFTRX1 R5_reg_18_ ( .D(R4[18]), .RN(n524), .CK(clk), .Q(R5[18]) );
  DFFTRX1 R7_reg_18_ ( .D(R6[18]), .RN(n524), .CK(clk), .Q(R7[18]) );
  DFFTRX1 R8_reg_18_ ( .D(R7[18]), .RN(n524), .CK(clk), .Q(R8[18]) );
  DFFTRX1 R9_reg_18_ ( .D(R8[18]), .RN(n524), .CK(clk), .Q(R9[18]) );
  DFFTRX1 R10_reg_18_ ( .D(R9[18]), .RN(n523), .CK(clk), .Q(R10[18]) );
  DFFTRX1 R11_reg_18_ ( .D(R10[18]), .RN(n523), .CK(clk), .Q(R11[18]) );
  DFFTRX1 R12_reg_18_ ( .D(R11[18]), .RN(n523), .CK(clk), .Q(R12[18]) );
  DFFTRX1 R13_reg_18_ ( .D(R12[18]), .RN(n523), .CK(clk), .Q(R13[18]) );
  DFFTRX1 R2_reg_17_ ( .D(R1[17]), .RN(n523), .CK(clk), .Q(R2[17]) );
  DFFTRX1 R3_reg_17_ ( .D(R2[17]), .RN(n523), .CK(clk), .Q(R3[17]) );
  DFFTRX1 R4_reg_17_ ( .D(R3[17]), .RN(n523), .CK(clk), .Q(R4[17]) );
  DFFTRX1 R5_reg_17_ ( .D(R4[17]), .RN(n523), .CK(clk), .Q(R5[17]) );
  DFFTRX1 R7_reg_17_ ( .D(R6[17]), .RN(n522), .CK(clk), .Q(R7[17]) );
  DFFTRX1 R8_reg_17_ ( .D(R7[17]), .RN(n522), .CK(clk), .Q(R8[17]) );
  DFFTRX1 R9_reg_17_ ( .D(R8[17]), .RN(n522), .CK(clk), .Q(R9[17]) );
  DFFTRX1 R10_reg_17_ ( .D(R9[17]), .RN(n522), .CK(clk), .Q(R10[17]) );
  DFFTRX1 R11_reg_17_ ( .D(R10[17]), .RN(n522), .CK(clk), .Q(R11[17]) );
  DFFTRX1 R12_reg_17_ ( .D(R11[17]), .RN(n522), .CK(clk), .Q(R12[17]) );
  DFFTRX1 R13_reg_17_ ( .D(R12[17]), .RN(n522), .CK(clk), .Q(R13[17]) );
  DFFTRX1 R2_reg_16_ ( .D(R1[16]), .RN(n522), .CK(clk), .Q(R2[16]) );
  DFFTRX1 R3_reg_16_ ( .D(R2[16]), .RN(n522), .CK(clk), .Q(R3[16]) );
  DFFTRX1 R4_reg_16_ ( .D(R3[16]), .RN(n521), .CK(clk), .Q(R4[16]) );
  DFFTRX1 R5_reg_16_ ( .D(R4[16]), .RN(n521), .CK(clk), .Q(R5[16]) );
  DFFTRX1 R7_reg_16_ ( .D(R6[16]), .RN(n521), .CK(clk), .Q(R7[16]) );
  DFFTRX1 R8_reg_16_ ( .D(R7[16]), .RN(n521), .CK(clk), .Q(R8[16]) );
  DFFTRX1 R9_reg_16_ ( .D(R8[16]), .RN(n521), .CK(clk), .Q(R9[16]) );
  DFFTRX1 R10_reg_16_ ( .D(R9[16]), .RN(n521), .CK(clk), .Q(R10[16]) );
  DFFTRX1 R11_reg_16_ ( .D(R10[16]), .RN(n521), .CK(clk), .Q(R11[16]) );
  DFFTRX1 R12_reg_16_ ( .D(R11[16]), .RN(n521), .CK(clk), .Q(R12[16]) );
  DFFTRX1 R13_reg_16_ ( .D(R12[16]), .RN(n521), .CK(clk), .Q(R13[16]) );
  DFFTRX1 R2_reg_15_ ( .D(R1[15]), .RN(n520), .CK(clk), .Q(R2[15]) );
  DFFTRX1 R3_reg_15_ ( .D(R2[15]), .RN(n520), .CK(clk), .Q(R3[15]) );
  DFFTRX1 R4_reg_15_ ( .D(R3[15]), .RN(n520), .CK(clk), .Q(R4[15]) );
  DFFTRX1 R5_reg_15_ ( .D(R4[15]), .RN(n520), .CK(clk), .Q(R5[15]) );
  DFFTRX1 R7_reg_15_ ( .D(R6[15]), .RN(n520), .CK(clk), .Q(R7[15]) );
  DFFTRX1 R8_reg_15_ ( .D(R7[15]), .RN(n520), .CK(clk), .Q(R8[15]) );
  DFFTRX1 R9_reg_15_ ( .D(R8[15]), .RN(n520), .CK(clk), .Q(R9[15]) );
  DFFTRX1 R10_reg_15_ ( .D(R9[15]), .RN(n520), .CK(clk), .Q(R10[15]) );
  DFFTRX1 R11_reg_15_ ( .D(R10[15]), .RN(n520), .CK(clk), .Q(R11[15]) );
  DFFTRX1 R12_reg_15_ ( .D(R11[15]), .RN(n520), .CK(clk), .Q(R12[15]) );
  DFFTRX1 R13_reg_15_ ( .D(R12[15]), .RN(n519), .CK(clk), .Q(R13[15]) );
  DFFTRX1 R2_reg_14_ ( .D(R1[14]), .RN(n519), .CK(clk), .Q(R2[14]) );
  DFFTRX1 R3_reg_14_ ( .D(R2[14]), .RN(n519), .CK(clk), .Q(R3[14]) );
  DFFTRX1 R4_reg_14_ ( .D(R3[14]), .RN(n519), .CK(clk), .Q(R4[14]) );
  DFFTRX1 R5_reg_14_ ( .D(R4[14]), .RN(n519), .CK(clk), .Q(R5[14]) );
  DFFTRX1 R7_reg_14_ ( .D(R6[14]), .RN(n519), .CK(clk), .Q(R7[14]) );
  DFFTRX1 R8_reg_14_ ( .D(R7[14]), .RN(n519), .CK(clk), .Q(R8[14]) );
  DFFTRX1 R9_reg_14_ ( .D(R8[14]), .RN(n519), .CK(clk), .Q(R9[14]) );
  DFFTRX1 R10_reg_14_ ( .D(R9[14]), .RN(n518), .CK(clk), .Q(R10[14]) );
  DFFTRX1 R11_reg_14_ ( .D(R10[14]), .RN(n518), .CK(clk), .Q(R11[14]) );
  DFFTRX1 R12_reg_14_ ( .D(R11[14]), .RN(n518), .CK(clk), .Q(R12[14]) );
  DFFTRX1 R13_reg_14_ ( .D(R12[14]), .RN(n518), .CK(clk), .Q(R13[14]) );
  DFFTRX1 R2_reg_13_ ( .D(R1[13]), .RN(n518), .CK(clk), .Q(R2[13]) );
  DFFTRX1 R3_reg_13_ ( .D(R2[13]), .RN(n518), .CK(clk), .Q(R3[13]) );
  DFFTRX1 R4_reg_13_ ( .D(R3[13]), .RN(n518), .CK(clk), .Q(R4[13]) );
  DFFTRX1 R5_reg_13_ ( .D(R4[13]), .RN(n518), .CK(clk), .Q(R5[13]) );
  DFFTRX1 R7_reg_13_ ( .D(R6[13]), .RN(n517), .CK(clk), .Q(R7[13]) );
  DFFTRX1 R8_reg_13_ ( .D(R7[13]), .RN(n517), .CK(clk), .Q(R8[13]) );
  DFFTRX1 R9_reg_13_ ( .D(R8[13]), .RN(n517), .CK(clk), .Q(R9[13]) );
  DFFTRX1 R10_reg_13_ ( .D(R9[13]), .RN(n517), .CK(clk), .Q(R10[13]) );
  DFFTRX1 R11_reg_13_ ( .D(R10[13]), .RN(n517), .CK(clk), .Q(R11[13]) );
  DFFTRX1 R12_reg_13_ ( .D(R11[13]), .RN(n517), .CK(clk), .Q(R12[13]) );
  DFFTRX1 R13_reg_13_ ( .D(R12[13]), .RN(n517), .CK(clk), .Q(R13[13]) );
  DFFTRX1 R2_reg_12_ ( .D(R1[12]), .RN(n517), .CK(clk), .Q(R2[12]) );
  DFFTRX1 R3_reg_12_ ( .D(R2[12]), .RN(n517), .CK(clk), .Q(R3[12]) );
  DFFTRX1 R4_reg_12_ ( .D(R3[12]), .RN(n516), .CK(clk), .Q(R4[12]) );
  DFFTRX1 R5_reg_12_ ( .D(R4[12]), .RN(n516), .CK(clk), .Q(R5[12]) );
  DFFTRX1 R7_reg_12_ ( .D(R6[12]), .RN(n516), .CK(clk), .Q(R7[12]) );
  DFFTRX1 R8_reg_12_ ( .D(R7[12]), .RN(n516), .CK(clk), .Q(R8[12]) );
  DFFTRX1 R9_reg_12_ ( .D(R8[12]), .RN(n516), .CK(clk), .Q(R9[12]) );
  DFFTRX1 R10_reg_12_ ( .D(R9[12]), .RN(n516), .CK(clk), .Q(R10[12]) );
  DFFTRX1 R11_reg_12_ ( .D(R10[12]), .RN(n516), .CK(clk), .Q(R11[12]) );
  DFFTRX1 R12_reg_12_ ( .D(R11[12]), .RN(n516), .CK(clk), .Q(R12[12]) );
  DFFTRX1 R13_reg_12_ ( .D(R12[12]), .RN(n516), .CK(clk), .Q(R13[12]) );
  DFFTRX1 R2_reg_11_ ( .D(R1[11]), .RN(n515), .CK(clk), .Q(R2[11]) );
  DFFTRX1 R3_reg_11_ ( .D(R2[11]), .RN(n515), .CK(clk), .Q(R3[11]) );
  DFFTRX1 R4_reg_11_ ( .D(R3[11]), .RN(n515), .CK(clk), .Q(R4[11]) );
  DFFTRX1 R5_reg_11_ ( .D(R4[11]), .RN(n515), .CK(clk), .Q(R5[11]) );
  DFFTRX1 R7_reg_11_ ( .D(R6[11]), .RN(n515), .CK(clk), .Q(R7[11]) );
  DFFTRX1 R8_reg_11_ ( .D(R7[11]), .RN(n515), .CK(clk), .Q(R8[11]) );
  DFFTRX1 R9_reg_11_ ( .D(R8[11]), .RN(n515), .CK(clk), .Q(R9[11]) );
  DFFTRX1 R10_reg_11_ ( .D(R9[11]), .RN(n515), .CK(clk), .Q(R10[11]) );
  DFFTRX1 R11_reg_11_ ( .D(R10[11]), .RN(n515), .CK(clk), .Q(R11[11]) );
  DFFTRX1 R12_reg_11_ ( .D(R11[11]), .RN(n515), .CK(clk), .Q(R12[11]) );
  DFFTRX1 R13_reg_11_ ( .D(R12[11]), .RN(n514), .CK(clk), .Q(R13[11]) );
  DFFTRX1 R2_reg_10_ ( .D(R1[10]), .RN(n514), .CK(clk), .Q(R2[10]) );
  DFFTRX1 R3_reg_10_ ( .D(R2[10]), .RN(n514), .CK(clk), .Q(R3[10]) );
  DFFTRX1 R4_reg_10_ ( .D(R3[10]), .RN(n514), .CK(clk), .Q(R4[10]) );
  DFFTRX1 R5_reg_10_ ( .D(R4[10]), .RN(n514), .CK(clk), .Q(R5[10]) );
  DFFTRX1 R7_reg_10_ ( .D(R6[10]), .RN(n514), .CK(clk), .Q(R7[10]) );
  DFFTRX1 R8_reg_10_ ( .D(R7[10]), .RN(n514), .CK(clk), .Q(R8[10]) );
  DFFTRX1 R9_reg_10_ ( .D(R8[10]), .RN(n514), .CK(clk), .Q(R9[10]) );
  DFFTRX1 R10_reg_10_ ( .D(R9[10]), .RN(n513), .CK(clk), .Q(R10[10]) );
  DFFTRX1 R11_reg_10_ ( .D(R10[10]), .RN(n513), .CK(clk), .Q(R11[10]) );
  DFFTRX1 R12_reg_10_ ( .D(R11[10]), .RN(n513), .CK(clk), .Q(R12[10]) );
  DFFTRX1 R13_reg_10_ ( .D(R12[10]), .RN(n513), .CK(clk), .Q(R13[10]) );
  DFFTRX1 R2_reg_9_ ( .D(R1[9]), .RN(n513), .CK(clk), .Q(R2[9]) );
  DFFTRX1 R3_reg_9_ ( .D(R2[9]), .RN(n513), .CK(clk), .Q(R3[9]) );
  DFFTRX1 R4_reg_9_ ( .D(R3[9]), .RN(n513), .CK(clk), .Q(R4[9]) );
  DFFTRX1 R5_reg_9_ ( .D(R4[9]), .RN(n513), .CK(clk), .Q(R5[9]) );
  DFFTRX1 R7_reg_9_ ( .D(R6[9]), .RN(n512), .CK(clk), .Q(R7[9]) );
  DFFTRX1 R8_reg_9_ ( .D(R7[9]), .RN(n512), .CK(clk), .Q(R8[9]) );
  DFFTRX1 R9_reg_9_ ( .D(R8[9]), .RN(n512), .CK(clk), .Q(R9[9]) );
  DFFTRX1 R10_reg_9_ ( .D(R9[9]), .RN(n512), .CK(clk), .Q(R10[9]) );
  DFFTRX1 R11_reg_9_ ( .D(R10[9]), .RN(n512), .CK(clk), .Q(R11[9]) );
  DFFTRX1 R12_reg_9_ ( .D(R11[9]), .RN(n512), .CK(clk), .Q(R12[9]) );
  DFFTRX1 R13_reg_9_ ( .D(R12[9]), .RN(n512), .CK(clk), .Q(R13[9]) );
  DFFTRX1 R2_reg_8_ ( .D(R1[8]), .RN(n512), .CK(clk), .Q(R2[8]) );
  DFFTRX1 R3_reg_8_ ( .D(R2[8]), .RN(n512), .CK(clk), .Q(R3[8]) );
  DFFTRX1 R4_reg_8_ ( .D(R3[8]), .RN(n511), .CK(clk), .Q(R4[8]) );
  DFFTRX1 R5_reg_8_ ( .D(R4[8]), .RN(n511), .CK(clk), .Q(R5[8]) );
  DFFTRX1 R7_reg_8_ ( .D(R6[8]), .RN(n511), .CK(clk), .Q(R7[8]) );
  DFFTRX1 R8_reg_8_ ( .D(R7[8]), .RN(n511), .CK(clk), .Q(R8[8]) );
  DFFTRX1 R9_reg_8_ ( .D(R8[8]), .RN(n511), .CK(clk), .Q(R9[8]) );
  DFFTRX1 R10_reg_8_ ( .D(R9[8]), .RN(n511), .CK(clk), .Q(R10[8]) );
  DFFTRX1 R11_reg_8_ ( .D(R10[8]), .RN(n511), .CK(clk), .Q(R11[8]) );
  DFFTRX1 R12_reg_8_ ( .D(R11[8]), .RN(n511), .CK(clk), .Q(R12[8]) );
  DFFTRX1 R13_reg_8_ ( .D(R12[8]), .RN(n511), .CK(clk), .Q(R13[8]) );
  DFFTRX1 R2_reg_7_ ( .D(R1[7]), .RN(n510), .CK(clk), .Q(R2[7]) );
  DFFTRX1 R3_reg_7_ ( .D(R2[7]), .RN(n510), .CK(clk), .Q(R3[7]) );
  DFFTRX1 R4_reg_7_ ( .D(R3[7]), .RN(n510), .CK(clk), .Q(R4[7]) );
  DFFTRX1 R5_reg_7_ ( .D(R4[7]), .RN(n510), .CK(clk), .Q(R5[7]) );
  DFFTRX1 R7_reg_7_ ( .D(R6[7]), .RN(n510), .CK(clk), .Q(R7[7]) );
  DFFTRX1 R8_reg_7_ ( .D(R7[7]), .RN(n510), .CK(clk), .Q(R8[7]) );
  DFFTRX1 R9_reg_7_ ( .D(R8[7]), .RN(n510), .CK(clk), .Q(R9[7]) );
  DFFTRX1 R10_reg_7_ ( .D(R9[7]), .RN(n510), .CK(clk), .Q(R10[7]) );
  DFFTRX1 R11_reg_7_ ( .D(R10[7]), .RN(n510), .CK(clk), .Q(R11[7]) );
  DFFTRX1 R12_reg_7_ ( .D(R11[7]), .RN(n510), .CK(clk), .Q(R12[7]) );
  DFFTRX1 R13_reg_7_ ( .D(R12[7]), .RN(n509), .CK(clk), .Q(R13[7]) );
  DFFTRX1 R2_reg_6_ ( .D(R1[6]), .RN(n509), .CK(clk), .Q(R2[6]) );
  DFFTRX1 R3_reg_6_ ( .D(R2[6]), .RN(n509), .CK(clk), .Q(R3[6]) );
  DFFTRX1 R4_reg_6_ ( .D(R3[6]), .RN(n509), .CK(clk), .Q(R4[6]) );
  DFFTRX1 R5_reg_6_ ( .D(R4[6]), .RN(n509), .CK(clk), .Q(R5[6]) );
  DFFTRX1 R7_reg_6_ ( .D(R6[6]), .RN(n509), .CK(clk), .Q(R7[6]) );
  DFFTRX1 R8_reg_6_ ( .D(R7[6]), .RN(n509), .CK(clk), .Q(R8[6]) );
  DFFTRX1 R9_reg_6_ ( .D(R8[6]), .RN(n509), .CK(clk), .Q(R9[6]) );
  DFFTRX1 R10_reg_6_ ( .D(R9[6]), .RN(n508), .CK(clk), .Q(R10[6]) );
  DFFTRX1 R11_reg_6_ ( .D(R10[6]), .RN(n508), .CK(clk), .Q(R11[6]) );
  DFFTRX1 R12_reg_6_ ( .D(R11[6]), .RN(n508), .CK(clk), .Q(R12[6]) );
  DFFTRX1 R13_reg_6_ ( .D(R12[6]), .RN(n508), .CK(clk), .Q(R13[6]) );
  DFFTRX1 R2_reg_5_ ( .D(R1[5]), .RN(n508), .CK(clk), .Q(R2[5]) );
  DFFTRX1 R3_reg_5_ ( .D(R2[5]), .RN(n508), .CK(clk), .Q(R3[5]) );
  DFFTRX1 R4_reg_5_ ( .D(R3[5]), .RN(n508), .CK(clk), .Q(R4[5]) );
  DFFTRX1 R5_reg_5_ ( .D(R4[5]), .RN(n508), .CK(clk), .Q(R5[5]) );
  DFFTRX1 R7_reg_5_ ( .D(R6[5]), .RN(n507), .CK(clk), .Q(R7[5]) );
  DFFTRX1 R8_reg_5_ ( .D(R7[5]), .RN(n507), .CK(clk), .Q(R8[5]) );
  DFFTRX1 R9_reg_5_ ( .D(R8[5]), .RN(n507), .CK(clk), .Q(R9[5]) );
  DFFTRX1 R10_reg_5_ ( .D(R9[5]), .RN(n507), .CK(clk), .Q(R10[5]) );
  DFFTRX1 R11_reg_5_ ( .D(R10[5]), .RN(n507), .CK(clk), .Q(R11[5]) );
  DFFTRX1 R12_reg_5_ ( .D(R11[5]), .RN(n507), .CK(clk), .Q(R12[5]) );
  DFFTRX1 R13_reg_5_ ( .D(R12[5]), .RN(n507), .CK(clk), .Q(R13[5]) );
  DFFTRX1 R2_reg_4_ ( .D(R1[4]), .RN(n507), .CK(clk), .Q(R2[4]) );
  DFFTRX1 R3_reg_4_ ( .D(R2[4]), .RN(n507), .CK(clk), .Q(R3[4]) );
  DFFTRX1 R4_reg_4_ ( .D(R3[4]), .RN(n506), .CK(clk), .Q(R4[4]) );
  DFFTRX1 R5_reg_4_ ( .D(R4[4]), .RN(n506), .CK(clk), .Q(R5[4]) );
  DFFTRX1 R7_reg_4_ ( .D(R6[4]), .RN(n506), .CK(clk), .Q(R7[4]) );
  DFFTRX1 R8_reg_4_ ( .D(R7[4]), .RN(n506), .CK(clk), .Q(R8[4]) );
  DFFTRX1 R9_reg_4_ ( .D(R8[4]), .RN(n506), .CK(clk), .Q(R9[4]) );
  DFFTRX1 R10_reg_4_ ( .D(R9[4]), .RN(n506), .CK(clk), .Q(R10[4]) );
  DFFTRX1 R11_reg_4_ ( .D(R10[4]), .RN(n506), .CK(clk), .Q(R11[4]) );
  DFFTRX1 R12_reg_4_ ( .D(R11[4]), .RN(n506), .CK(clk), .Q(R12[4]) );
  DFFTRX1 R13_reg_4_ ( .D(R12[4]), .RN(n506), .CK(clk), .Q(R13[4]) );
  DFFTRX1 R2_reg_3_ ( .D(R1[3]), .RN(n505), .CK(clk), .Q(R2[3]) );
  DFFTRX1 R3_reg_3_ ( .D(R2[3]), .RN(n505), .CK(clk), .Q(R3[3]) );
  DFFTRX1 R4_reg_3_ ( .D(R3[3]), .RN(n505), .CK(clk), .Q(R4[3]) );
  DFFTRX1 R5_reg_3_ ( .D(R4[3]), .RN(n505), .CK(clk), .Q(R5[3]) );
  DFFTRX1 R7_reg_3_ ( .D(R6[3]), .RN(n505), .CK(clk), .Q(R7[3]) );
  DFFTRX1 R8_reg_3_ ( .D(R7[3]), .RN(n505), .CK(clk), .Q(R8[3]) );
  DFFTRX1 R9_reg_3_ ( .D(R8[3]), .RN(n505), .CK(clk), .Q(R9[3]) );
  DFFTRX1 R10_reg_3_ ( .D(R9[3]), .RN(n505), .CK(clk), .Q(R10[3]) );
  DFFTRX1 R11_reg_3_ ( .D(R10[3]), .RN(n505), .CK(clk), .Q(R11[3]) );
  DFFTRX1 R12_reg_3_ ( .D(R11[3]), .RN(n505), .CK(clk), .Q(R12[3]) );
  DFFTRX1 R13_reg_3_ ( .D(R12[3]), .RN(n504), .CK(clk), .Q(R13[3]) );
  DFFTRX1 R2_reg_2_ ( .D(R1[2]), .RN(n504), .CK(clk), .Q(R2[2]) );
  DFFTRX1 R3_reg_2_ ( .D(R2[2]), .RN(n504), .CK(clk), .Q(R3[2]) );
  DFFTRX1 R4_reg_2_ ( .D(R3[2]), .RN(n504), .CK(clk), .Q(R4[2]) );
  DFFTRX1 R5_reg_2_ ( .D(R4[2]), .RN(n504), .CK(clk), .Q(R5[2]) );
  DFFTRX1 R7_reg_2_ ( .D(R6[2]), .RN(n504), .CK(clk), .Q(R7[2]) );
  DFFTRX1 R8_reg_2_ ( .D(R7[2]), .RN(n504), .CK(clk), .Q(R8[2]) );
  DFFTRX1 R9_reg_2_ ( .D(R8[2]), .RN(n504), .CK(clk), .Q(R9[2]) );
  DFFTRX1 R10_reg_2_ ( .D(R9[2]), .RN(n503), .CK(clk), .Q(R10[2]) );
  DFFTRX1 R11_reg_2_ ( .D(R10[2]), .RN(n503), .CK(clk), .Q(R11[2]) );
  DFFTRX1 R12_reg_2_ ( .D(R11[2]), .RN(n503), .CK(clk), .Q(R12[2]) );
  DFFTRX1 R13_reg_2_ ( .D(R12[2]), .RN(n503), .CK(clk), .Q(R13[2]) );
  DFFTRX1 R2_reg_1_ ( .D(R1[1]), .RN(n503), .CK(clk), .Q(R2[1]) );
  DFFTRX1 R3_reg_1_ ( .D(R2[1]), .RN(n503), .CK(clk), .Q(R3[1]) );
  DFFTRX1 R4_reg_1_ ( .D(R3[1]), .RN(n503), .CK(clk), .Q(R4[1]) );
  DFFTRX1 R5_reg_1_ ( .D(R4[1]), .RN(n503), .CK(clk), .Q(R5[1]) );
  DFFTRX1 R7_reg_1_ ( .D(R6[1]), .RN(n502), .CK(clk), .Q(R7[1]) );
  DFFTRX1 R8_reg_1_ ( .D(R7[1]), .RN(n502), .CK(clk), .Q(R8[1]) );
  DFFTRX1 R9_reg_1_ ( .D(R8[1]), .RN(n502), .CK(clk), .Q(R9[1]) );
  DFFTRX1 R10_reg_1_ ( .D(R9[1]), .RN(n502), .CK(clk), .Q(R10[1]) );
  DFFTRX1 R11_reg_1_ ( .D(R10[1]), .RN(n502), .CK(clk), .Q(R11[1]) );
  DFFTRX1 R12_reg_1_ ( .D(R11[1]), .RN(n502), .CK(clk), .Q(R12[1]) );
  DFFTRX1 R13_reg_1_ ( .D(R12[1]), .RN(n502), .CK(clk), .Q(R13[1]) );
  DFFTRX1 R2_reg_0_ ( .D(R1[0]), .RN(n502), .CK(clk), .Q(R2[0]) );
  DFFTRX1 R3_reg_0_ ( .D(R2[0]), .RN(n502), .CK(clk), .Q(R3[0]) );
  DFFHQXL Wt_reg_25_ ( .D(n617), .CK(clk), .Q(Wt[25]) );
  DFFHQXL Wt_reg_27_ ( .D(n612), .CK(clk), .Q(Wt[27]) );
  DFFHQXL Wt_reg_26_ ( .D(n616), .CK(clk), .Q(Wt[26]) );
  DFFHQX1 Wt_reg_24_ ( .D(n618), .CK(clk), .Q(Wt[24]) );
  DFFTRX1 R15_reg_2_ ( .D(R14[2]), .RN(n503), .CK(clk), .Q(R15[2]) );
  DFFTRX1 R6_reg_2_ ( .D(R5[2]), .RN(n504), .CK(clk), .Q(R6[2]) );
  DFFHQX2 Wt_reg_18_ ( .D(n624), .CK(clk), .Q(Wt[18]) );
  DFFHQX2 Wt_reg_17_ ( .D(n625), .CK(clk), .Q(Wt[17]) );
  DFFTRX2 R14_reg_22_ ( .D(R13[22]), .RN(n528), .CK(clk), .Q(R14[22]) );
  DFFX4 Wt_reg_1_ ( .D(n641), .CK(clk), .Q(Wt[1]), .QN(n14) );
  DFFTRX1 R14_reg_12_ ( .D(R13[12]), .RN(n516), .CK(clk), .Q(R14[12]) );
  DFFTRX1 R1_reg_18_ ( .D(Wt[18]), .RN(n524), .CK(clk), .Q(R1[18]) );
  DFFTRX1 R1_reg_17_ ( .D(Wt[17]), .RN(n523), .CK(clk), .Q(R1[17]) );
  DFFTRX2 R1_reg_21_ ( .D(Wt[21]), .RN(n528), .CK(clk), .Q(R1[21]) );
  DFFHQX1 Wt_reg_21_ ( .D(n621), .CK(clk), .Q(Wt[21]) );
  DFFTRX1 R14_reg_21_ ( .D(R13[21]), .RN(n527), .CK(clk), .Q(R14[21]) );
  DFFTRX1 R1_reg_20_ ( .D(Wt[20]), .RN(n527), .CK(clk), .Q(R1[20]) );
  DFFHQX1 Wt_reg_20_ ( .D(n622), .CK(clk), .Q(Wt[20]) );
  DFFTRX1 R1_reg_1_ ( .D(n17), .RN(n503), .CK(clk), .Q(R1[1]) );
  DFFTRX1 R14_reg_20_ ( .D(R13[20]), .RN(n526), .CK(clk), .Q(R14[20]) );
  DFFTRX1 R14_reg_23_ ( .D(R13[23]), .RN(n529), .CK(clk), .Q(R14[23]) );
  DFFTRX2 R7_reg_0_ ( .D(R6[0]), .RN(n501), .CK(clk), .Q(R7[0]) );
  DFFTRX2 R14_reg_11_ ( .D(R13[11]), .RN(n514), .CK(clk), .Q(R14[11]) );
  DFFTRX2 R1_reg_23_ ( .D(Wt[23]), .RN(n530), .CK(clk), .Q(R1[23]) );
  DFFHQXL Wt_reg_23_ ( .D(n619), .CK(clk), .Q(Wt[23]) );
  XOR3X4 U3 ( .A(R14[22]), .B(R14[11]), .C(R14[7]), .Y(sigma0[4]) );
  XOR3X2 U4 ( .A(R14[23]), .B(R14[12]), .C(R14[8]), .Y(sigma0[5]) );
  XOR3X2 U5 ( .A(R14[26]), .B(R14[15]), .C(R14[11]), .Y(sigma0[8]) );
  OAI2BB1X2 U6 ( .A0N(logic_result[27]), .A1N(n496), .B0(n602), .Y(n612) );
  INVX1 U7 ( .A(logic_result[15]), .Y(n585) );
  OAI22X1 U8 ( .A0(n21), .A1(n586), .B0(n594), .B1(n585), .Y(n627) );
  BUFX16 U9 ( .A(n647), .Y(Wt[0]) );
  INVX1 U10 ( .A(n14), .Y(n17) );
  CLKINVX3 U11 ( .A(n377), .Y(n594) );
  XOR2X1 U12 ( .A(R1[13]), .B(R1[15]), .Y(sigma1[28]) );
  OAI2BB1X4 U13 ( .A0N(logic_result[31]), .A1N(n496), .B0(n607), .Y(n608) );
  OAI2BB1X4 U14 ( .A0N(logic_result[30]), .A1N(n496), .B0(n605), .Y(n609) );
  OAI2BB1X2 U15 ( .A0N(logic_result[29]), .A1N(n496), .B0(n604), .Y(n610) );
  NAND2XL U16 ( .A(inner_busy), .B(n613), .Y(n578) );
  XOR2XL U17 ( .A(R1[16]), .B(R1[18]), .Y(sigma1[31]) );
  NAND2XL U18 ( .A(write_enable), .B(n553), .Y(n21) );
  NAND2XL U19 ( .A(write_enable), .B(n553), .Y(n23) );
  NAND2XL U20 ( .A(write_enable), .B(n553), .Y(n24) );
  XOR2XL U21 ( .A(R1[10]), .B(R1[12]), .Y(sigma1[25]) );
  XOR2XL U22 ( .A(R1[8]), .B(R1[10]), .Y(sigma1[23]) );
  XOR2XL U23 ( .A(R1[9]), .B(R1[11]), .Y(sigma1[24]) );
  XOR2XL U24 ( .A(R1[11]), .B(R1[13]), .Y(sigma1[26]) );
  INVX1 U25 ( .A(n541), .Y(n503) );
  INVX1 U26 ( .A(n551), .Y(n506) );
  INVX1 U27 ( .A(n551), .Y(n507) );
  INVX1 U28 ( .A(n550), .Y(n508) );
  INVX1 U29 ( .A(n550), .Y(n509) );
  INVX1 U30 ( .A(n549), .Y(n510) );
  INVX1 U31 ( .A(n549), .Y(n511) );
  INVX1 U32 ( .A(n548), .Y(n512) );
  INVX1 U33 ( .A(n548), .Y(n513) );
  INVX1 U34 ( .A(n547), .Y(n514) );
  INVX1 U35 ( .A(n547), .Y(n515) );
  INVX1 U36 ( .A(n546), .Y(n516) );
  INVX1 U37 ( .A(n546), .Y(n517) );
  INVX1 U38 ( .A(n545), .Y(n518) );
  INVX1 U39 ( .A(n545), .Y(n519) );
  INVX1 U40 ( .A(n545), .Y(n520) );
  INVX1 U41 ( .A(n545), .Y(n521) );
  INVX1 U42 ( .A(n541), .Y(n522) );
  INVX1 U43 ( .A(n542), .Y(n523) );
  INVX1 U44 ( .A(n544), .Y(n524) );
  INVX1 U45 ( .A(n544), .Y(n525) );
  INVX1 U46 ( .A(n543), .Y(n526) );
  INVX1 U47 ( .A(n544), .Y(n527) );
  INVX1 U48 ( .A(n542), .Y(n528) );
  INVX1 U49 ( .A(n541), .Y(n529) );
  INVX1 U50 ( .A(n543), .Y(n530) );
  INVX1 U51 ( .A(n543), .Y(n531) );
  INVX1 U52 ( .A(n541), .Y(n532) );
  INVX1 U53 ( .A(n543), .Y(n533) );
  INVX1 U54 ( .A(n542), .Y(n534) );
  INVX1 U55 ( .A(n541), .Y(n535) );
  INVX1 U56 ( .A(n542), .Y(n502) );
  INVX1 U57 ( .A(n541), .Y(n504) );
  INVX1 U58 ( .A(n542), .Y(n505) );
  INVX1 U59 ( .A(n552), .Y(n501) );
  INVX1 U60 ( .A(n499), .Y(n552) );
  INVX1 U61 ( .A(n542), .Y(n536) );
  INVX1 U62 ( .A(n542), .Y(n537) );
  INVX1 U63 ( .A(n542), .Y(n538) );
  INVX1 U64 ( .A(n541), .Y(n539) );
  INVX1 U65 ( .A(n541), .Y(n540) );
  INVX1 U66 ( .A(n499), .Y(n551) );
  INVX1 U67 ( .A(n499), .Y(n550) );
  INVX1 U68 ( .A(n499), .Y(n549) );
  INVX1 U69 ( .A(n498), .Y(n548) );
  INVX1 U70 ( .A(n498), .Y(n547) );
  INVX1 U71 ( .A(n498), .Y(n546) );
  INVX1 U72 ( .A(n498), .Y(n545) );
  INVX1 U73 ( .A(n497), .Y(n544) );
  INVX1 U74 ( .A(n497), .Y(n543) );
  INVX1 U75 ( .A(n500), .Y(n499) );
  INVX1 U76 ( .A(n500), .Y(n498) );
  INVX1 U77 ( .A(n500), .Y(n497) );
  INVX1 U78 ( .A(n643), .Y(n542) );
  INVX1 U79 ( .A(n643), .Y(n541) );
  INVX1 U80 ( .A(n643), .Y(n500) );
  INVX1 U81 ( .A(n578), .Y(n553) );
  INVX1 U82 ( .A(n578), .Y(n643) );
  INVX1 U83 ( .A(n21), .Y(n606) );
  BUFX3 U84 ( .A(n377), .Y(n496) );
  OAI2BB1X1 U85 ( .A0N(logic_result[28]), .A1N(n496), .B0(n603), .Y(n611) );
  NAND2X1 U86 ( .A(data[28]), .B(n606), .Y(n603) );
  NAND2X1 U87 ( .A(data[29]), .B(n606), .Y(n604) );
  NAND2X1 U88 ( .A(data[30]), .B(n606), .Y(n605) );
  NAND2X1 U89 ( .A(data[31]), .B(n606), .Y(n607) );
  OAI2BB1X1 U90 ( .A0N(logic_result[25]), .A1N(n496), .B0(n600), .Y(n617) );
  NAND2X1 U91 ( .A(data[25]), .B(n606), .Y(n600) );
  OAI2BB1X1 U92 ( .A0N(logic_result[26]), .A1N(n496), .B0(n601), .Y(n616) );
  NAND2X1 U93 ( .A(data[26]), .B(n606), .Y(n601) );
  NAND2X1 U94 ( .A(data[27]), .B(n606), .Y(n602) );
  OAI2BB1X1 U95 ( .A0N(logic_result[22]), .A1N(n496), .B0(n597), .Y(n620) );
  NAND2X1 U96 ( .A(data[22]), .B(n606), .Y(n597) );
  OAI2BB1X1 U97 ( .A0N(logic_result[23]), .A1N(n496), .B0(n598), .Y(n619) );
  NAND2X1 U98 ( .A(data[23]), .B(n606), .Y(n598) );
  OAI2BB1X1 U99 ( .A0N(logic_result[24]), .A1N(n496), .B0(n599), .Y(n618) );
  NAND2X1 U100 ( .A(data[24]), .B(n606), .Y(n599) );
  INVX1 U101 ( .A(logic_result[3]), .Y(n560) );
  INVX1 U102 ( .A(data[3]), .Y(n561) );
  XOR3X2 U103 ( .A(R14[18]), .B(R14[7]), .C(R14[3]), .Y(sigma0[0]) );
  XOR3X2 U104 ( .A(R1[19]), .B(R1[17]), .C(R1[10]), .Y(sigma1[0]) );
  AOI31X1 U105 ( .A0(n614), .A1(counter[6]), .A2(n615), .B0(reset), .Y(n613)
         );
  NOR2X1 U106 ( .A(counter[1]), .B(counter[0]), .Y(n614) );
  NOR4X1 U107 ( .A(counter[5]), .B(counter[4]), .C(counter[3]), .D(counter[2]), 
        .Y(n615) );
  OAI22XL U108 ( .A0(n24), .A1(n555), .B0(n594), .B1(n554), .Y(n642) );
  INVX1 U109 ( .A(logic_result[0]), .Y(n554) );
  INVX1 U110 ( .A(data[0]), .Y(n555) );
  OAI22XL U111 ( .A0(n21), .A1(n557), .B0(n594), .B1(n556), .Y(n641) );
  INVX1 U112 ( .A(logic_result[1]), .Y(n556) );
  INVX1 U113 ( .A(data[1]), .Y(n557) );
  OAI22XL U114 ( .A0(n23), .A1(n559), .B0(n594), .B1(n558), .Y(n640) );
  INVX1 U115 ( .A(logic_result[2]), .Y(n558) );
  INVX1 U116 ( .A(data[2]), .Y(n559) );
  OAI22XL U117 ( .A0(n24), .A1(n563), .B0(n594), .B1(n562), .Y(n638) );
  INVX1 U118 ( .A(logic_result[4]), .Y(n562) );
  INVX1 U119 ( .A(data[4]), .Y(n563) );
  OAI22XL U120 ( .A0(n21), .A1(n565), .B0(n594), .B1(n564), .Y(n637) );
  INVX1 U121 ( .A(logic_result[5]), .Y(n564) );
  INVX1 U122 ( .A(data[5]), .Y(n565) );
  OAI22XL U123 ( .A0(n21), .A1(n567), .B0(n594), .B1(n566), .Y(n636) );
  INVX1 U124 ( .A(logic_result[6]), .Y(n566) );
  INVX1 U125 ( .A(data[6]), .Y(n567) );
  OAI22XL U126 ( .A0(n23), .A1(n569), .B0(n594), .B1(n568), .Y(n635) );
  INVX1 U127 ( .A(logic_result[7]), .Y(n568) );
  INVX1 U128 ( .A(data[7]), .Y(n569) );
  OAI22XL U129 ( .A0(n24), .A1(n571), .B0(n594), .B1(n570), .Y(n634) );
  INVX1 U130 ( .A(logic_result[8]), .Y(n570) );
  INVX1 U131 ( .A(data[8]), .Y(n571) );
  OAI22XL U132 ( .A0(n24), .A1(n573), .B0(n594), .B1(n572), .Y(n633) );
  INVX1 U133 ( .A(logic_result[9]), .Y(n572) );
  INVX1 U134 ( .A(data[9]), .Y(n573) );
  OAI22XL U135 ( .A0(n21), .A1(n575), .B0(n594), .B1(n574), .Y(n632) );
  INVX1 U136 ( .A(logic_result[10]), .Y(n574) );
  INVX1 U137 ( .A(data[10]), .Y(n575) );
  OAI22XL U138 ( .A0(n23), .A1(n577), .B0(n594), .B1(n576), .Y(n631) );
  INVX1 U139 ( .A(logic_result[11]), .Y(n576) );
  INVX1 U140 ( .A(data[11]), .Y(n577) );
  OAI22XL U141 ( .A0(n23), .A1(n580), .B0(n594), .B1(n579), .Y(n630) );
  INVX1 U142 ( .A(logic_result[12]), .Y(n579) );
  INVX1 U143 ( .A(data[12]), .Y(n580) );
  OAI22XL U144 ( .A0(n24), .A1(n582), .B0(n594), .B1(n581), .Y(n629) );
  INVX1 U145 ( .A(logic_result[13]), .Y(n581) );
  INVX1 U146 ( .A(data[13]), .Y(n582) );
  OAI22XL U147 ( .A0(n21), .A1(n584), .B0(n594), .B1(n583), .Y(n628) );
  INVX1 U148 ( .A(logic_result[14]), .Y(n583) );
  INVX1 U149 ( .A(data[14]), .Y(n584) );
  INVX1 U150 ( .A(data[15]), .Y(n586) );
  OAI22XL U151 ( .A0(n23), .A1(n588), .B0(n594), .B1(n587), .Y(n626) );
  INVX1 U152 ( .A(logic_result[16]), .Y(n587) );
  INVX1 U153 ( .A(data[16]), .Y(n588) );
  OAI22XL U154 ( .A0(n24), .A1(n590), .B0(n594), .B1(n589), .Y(n625) );
  INVX1 U155 ( .A(logic_result[17]), .Y(n589) );
  INVX1 U156 ( .A(data[17]), .Y(n590) );
  OAI22XL U157 ( .A0(n24), .A1(n592), .B0(n594), .B1(n591), .Y(n624) );
  INVX1 U158 ( .A(data[18]), .Y(n592) );
  INVX1 U159 ( .A(logic_result[18]), .Y(n591) );
  NOR2BX1 U160 ( .AN(n553), .B(write_enable), .Y(n377) );
  XOR3X2 U161 ( .A(R14[27]), .B(R14[16]), .C(R14[12]), .Y(sigma0[9]) );
  XOR3X2 U162 ( .A(R14[21]), .B(R14[10]), .C(R14[6]), .Y(sigma0[3]) );
  XOR3X2 U163 ( .A(R14[20]), .B(R14[9]), .C(R14[5]), .Y(sigma0[2]) );
  XOR3X2 U164 ( .A(R14[19]), .B(R14[8]), .C(R14[4]), .Y(sigma0[1]) );
  XOR3X2 U165 ( .A(R14[25]), .B(R14[14]), .C(R14[10]), .Y(sigma0[7]) );
  XOR3X2 U166 ( .A(R14[24]), .B(R14[13]), .C(R14[9]), .Y(sigma0[6]) );
  XOR3X2 U167 ( .A(R1[20]), .B(R1[18]), .C(R1[11]), .Y(sigma1[1]) );
  XOR3X2 U168 ( .A(R1[20]), .B(R1[22]), .C(R1[13]), .Y(sigma1[3]) );
  XOR3X2 U169 ( .A(R1[19]), .B(R1[21]), .C(R1[12]), .Y(sigma1[2]) );
  XOR3X2 U170 ( .A(R1[22]), .B(R1[24]), .C(R1[15]), .Y(sigma1[5]) );
  XOR3X2 U171 ( .A(R1[24]), .B(R1[26]), .C(R1[17]), .Y(sigma1[7]) );
  XOR3X2 U172 ( .A(R1[26]), .B(R1[28]), .C(R1[19]), .Y(sigma1[9]) );
  XOR3X2 U173 ( .A(R1[23]), .B(R1[25]), .C(R1[16]), .Y(sigma1[6]) );
  XOR3X2 U174 ( .A(R1[21]), .B(R1[23]), .C(R1[14]), .Y(sigma1[4]) );
  OAI2BB2X1 U175 ( .B0(n594), .B1(n593), .A0N(data[19]), .A1N(n606), .Y(n623)
         );
  INVX1 U176 ( .A(logic_result[19]), .Y(n593) );
  OAI2BB1X1 U177 ( .A0N(logic_result[20]), .A1N(n496), .B0(n595), .Y(n622) );
  NAND2X1 U178 ( .A(data[20]), .B(n606), .Y(n595) );
  OAI2BB1X1 U179 ( .A0N(logic_result[21]), .A1N(n496), .B0(n596), .Y(n621) );
  NAND2X1 U180 ( .A(data[21]), .B(n606), .Y(n596) );
  XOR3X2 U181 ( .A(R14[18]), .B(R14[29]), .C(R14[14]), .Y(sigma0[11]) );
  XOR3X2 U182 ( .A(R14[19]), .B(R14[30]), .C(R14[15]), .Y(sigma0[12]) );
  XOR3X2 U183 ( .A(R14[20]), .B(R14[31]), .C(R14[16]), .Y(sigma0[13]) );
  XOR3X2 U184 ( .A(R14[21]), .B(R14[17]), .C(R14[0]), .Y(sigma0[14]) );
  XOR3X2 U185 ( .A(R14[28]), .B(R14[17]), .C(R14[13]), .Y(sigma0[10]) );
  XOR3X2 U186 ( .A(R1[25]), .B(R1[2]), .C(R1[0]), .Y(sigma1[15]) );
  XOR3X2 U187 ( .A(R1[26]), .B(R1[3]), .C(R1[1]), .Y(sigma1[16]) );
  XOR3X2 U188 ( .A(R14[18]), .B(R14[22]), .C(R14[1]), .Y(sigma0[15]) );
  XOR3X2 U189 ( .A(R14[20]), .B(R14[24]), .C(R14[3]), .Y(sigma0[17]) );
  XOR3X2 U190 ( .A(R14[22]), .B(R14[26]), .C(R14[5]), .Y(sigma0[19]) );
  XOR3X2 U191 ( .A(R14[21]), .B(R14[25]), .C(R14[4]), .Y(sigma0[18]) );
  XOR3X2 U192 ( .A(R1[28]), .B(R1[30]), .C(R1[21]), .Y(sigma1[11]) );
  XOR3X2 U193 ( .A(R1[24]), .B(R1[31]), .C(R1[1]), .Y(sigma1[14]) );
  XOR3X2 U194 ( .A(R1[29]), .B(R1[31]), .C(R1[22]), .Y(sigma1[12]) );
  XOR3X2 U195 ( .A(R1[23]), .B(R1[30]), .C(R1[0]), .Y(sigma1[13]) );
  XOR3X2 U196 ( .A(R1[25]), .B(R1[27]), .C(R1[18]), .Y(sigma1[8]) );
  XOR3X2 U197 ( .A(R1[27]), .B(R1[29]), .C(R1[20]), .Y(sigma1[10]) );
  XOR3X2 U198 ( .A(R1[27]), .B(R1[4]), .C(R1[2]), .Y(sigma1[17]) );
  XOR3X2 U199 ( .A(R1[29]), .B(R1[6]), .C(R1[4]), .Y(sigma1[19]) );
  XOR3X2 U200 ( .A(R1[28]), .B(R1[5]), .C(R1[3]), .Y(sigma1[18]) );
  XOR2X1 U201 ( .A(R14[6]), .B(R14[17]), .Y(sigma0[31]) );
  XOR3X2 U202 ( .A(R14[26]), .B(R14[30]), .C(R14[9]), .Y(sigma0[23]) );
  XOR3X2 U203 ( .A(R14[25]), .B(R14[29]), .C(R14[8]), .Y(sigma0[22]) );
  XOR3X2 U204 ( .A(R14[24]), .B(R14[28]), .C(R14[7]), .Y(sigma0[21]) );
  XOR3X2 U205 ( .A(R14[19]), .B(R14[23]), .C(R14[2]), .Y(sigma0[16]) );
  XOR3X2 U206 ( .A(R14[23]), .B(R14[27]), .C(R14[6]), .Y(sigma0[20]) );
  XOR3X2 U207 ( .A(R1[30]), .B(R1[7]), .C(R1[5]), .Y(sigma1[20]) );
  XOR3X2 U208 ( .A(R1[31]), .B(R1[8]), .C(R1[6]), .Y(sigma1[21]) );
  XOR2X1 U209 ( .A(R1[7]), .B(R1[9]), .Y(sigma1[22]) );
  XOR3X2 U210 ( .A(R14[27]), .B(R14[31]), .C(R14[10]), .Y(sigma0[24]) );
  XOR3X2 U211 ( .A(R14[13]), .B(R14[30]), .C(R14[2]), .Y(sigma0[27]) );
  XOR3X2 U212 ( .A(R14[12]), .B(R14[29]), .C(R14[1]), .Y(sigma0[26]) );
  XOR3X2 U213 ( .A(R14[11]), .B(R14[28]), .C(R14[0]), .Y(sigma0[25]) );
  XOR2X1 U214 ( .A(R1[12]), .B(R1[14]), .Y(sigma1[27]) );
  XOR3X2 U215 ( .A(R14[14]), .B(R14[31]), .C(R14[3]), .Y(sigma0[28]) );
  XOR2X1 U216 ( .A(R14[4]), .B(R14[15]), .Y(sigma0[29]) );
  XOR2X1 U217 ( .A(R14[5]), .B(R14[16]), .Y(sigma0[30]) );
  XOR2X1 U218 ( .A(R1[14]), .B(R1[16]), .Y(sigma1[29]) );
  XOR2X1 U219 ( .A(R1[15]), .B(R1[17]), .Y(sigma1[30]) );
  OAI22X1 U220 ( .A0(n23), .A1(n561), .B0(n594), .B1(n560), .Y(n639) );
endmodule


module hash_core_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;
  wire   [31:2] carry;

  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_1 ( .A(A[1]), .B(B[1]), .CI(n29), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX4 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX4 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX4 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX4 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX4 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX4 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX4 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  NAND2X4 U1 ( .A(B[13]), .B(carry[13]), .Y(n9) );
  NAND2X2 U2 ( .A(B[21]), .B(n19), .Y(n22) );
  AND2X4 U3 ( .A(n23), .B(n21), .Y(n1) );
  NAND2BX4 U4 ( .AN(n5), .B(carry[21]), .Y(n21) );
  NAND2X4 U5 ( .A(n1), .B(n22), .Y(carry[22]) );
  NAND3X4 U6 ( .A(n26), .B(n28), .C(n27), .Y(carry[4]) );
  NAND2X4 U7 ( .A(A[3]), .B(carry[3]), .Y(n27) );
  NAND2X4 U8 ( .A(B[26]), .B(carry[26]), .Y(n13) );
  ADDFHX2 U9 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(n4) );
  INVX1 U10 ( .A(B[3]), .Y(n2) );
  INVX1 U11 ( .A(A[31]), .Y(n3) );
  ADDFHX2 U12 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(n6) );
  INVX1 U13 ( .A(A[21]), .Y(n5) );
  NAND2X1 U14 ( .A(B[21]), .B(A[21]), .Y(n23) );
  ADDFHX2 U15 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(n19) );
  NAND2BX4 U16 ( .AN(n2), .B(n24), .Y(n26) );
  XNOR3X4 U17 ( .A(n3), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  XOR2X1 U18 ( .A(A[13]), .B(B[13]), .Y(n7) );
  XOR2X1 U19 ( .A(carry[13]), .B(n7), .Y(SUM[13]) );
  NAND2X2 U20 ( .A(carry[13]), .B(A[13]), .Y(n8) );
  NAND2X4 U21 ( .A(B[13]), .B(A[13]), .Y(n10) );
  NAND3X4 U22 ( .A(n9), .B(n8), .C(n10), .Y(carry[14]) );
  XOR2X1 U23 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U24 ( .A(A[26]), .B(B[26]), .Y(n11) );
  XOR2X1 U25 ( .A(carry[26]), .B(n11), .Y(SUM[26]) );
  NAND2X4 U26 ( .A(A[26]), .B(n4), .Y(n12) );
  NAND2X4 U27 ( .A(B[26]), .B(A[26]), .Y(n14) );
  NAND3X4 U28 ( .A(n14), .B(n12), .C(n13), .Y(carry[27]) );
  XOR2X1 U29 ( .A(A[29]), .B(B[29]), .Y(n15) );
  XOR2X1 U30 ( .A(carry[29]), .B(n15), .Y(SUM[29]) );
  NAND2X4 U31 ( .A(A[29]), .B(n6), .Y(n16) );
  NAND2X4 U32 ( .A(B[29]), .B(carry[29]), .Y(n17) );
  NAND2X4 U33 ( .A(B[29]), .B(A[29]), .Y(n18) );
  NAND3X4 U34 ( .A(n18), .B(n16), .C(n17), .Y(carry[30]) );
  XOR2X1 U35 ( .A(A[21]), .B(B[21]), .Y(n20) );
  XOR2X1 U36 ( .A(n19), .B(n20), .Y(SUM[21]) );
  AND2X4 U37 ( .A(B[0]), .B(A[0]), .Y(n29) );
  XOR2X1 U38 ( .A(B[3]), .B(A[3]), .Y(n25) );
  ADDFHX4 U39 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(n24) );
  NAND2XL U40 ( .A(A[3]), .B(B[3]), .Y(n28) );
  XOR2X1 U41 ( .A(n24), .B(n25), .Y(SUM[3]) );
endmodule


module hash_core_DW01_add_1 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45;
  wire   [31:2] carry;

  ADDFHX4 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX4 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX4 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX4 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX4 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(n6), .CO(carry[29]), .S(SUM[28])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX4 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX4 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX4 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX4 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX4 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_1 ( .A(A[1]), .B(B[1]), .CI(n45), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX4 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  XNOR2X4 U1 ( .A(carry[31]), .B(n1), .Y(SUM[31]) );
  CLKINVX20 U2 ( .A(n38), .Y(n1) );
  AND2X4 U3 ( .A(B[0]), .B(A[0]), .Y(n45) );
  NAND2X4 U4 ( .A(carry[12]), .B(B[12]), .Y(n19) );
  XOR2XL U5 ( .A(B[5]), .B(A[5]), .Y(n30) );
  NAND2XL U6 ( .A(A[5]), .B(B[5]), .Y(n33) );
  ADDFHX2 U7 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(n8) );
  NAND2X4 U8 ( .A(B[5]), .B(n3), .Y(n31) );
  ADDFHX4 U9 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(n3) );
  NAND3X4 U10 ( .A(n19), .B(n20), .C(n21), .Y(carry[13]) );
  NAND2XL U11 ( .A(B[11]), .B(A[11]), .Y(n17) );
  INVX1 U12 ( .A(A[27]), .Y(n13) );
  INVX1 U13 ( .A(B[27]), .Y(n9) );
  INVX1 U14 ( .A(A[24]), .Y(n12) );
  NAND2X1 U15 ( .A(B[24]), .B(A[24]), .Y(n37) );
  AND2X4 U16 ( .A(n35), .B(n37), .Y(n2) );
  ADDFHX4 U17 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(n4) );
  ADDFHX4 U18 ( .A(A[28]), .B(B[28]), .CI(n6), .CO(n5) );
  NAND2X4 U19 ( .A(n40), .B(n43), .Y(n6) );
  ADDFHX2 U20 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(n10) );
  NAND2BX2 U21 ( .AN(n9), .B(carry[27]), .Y(n43) );
  NAND3X2 U22 ( .A(n15), .B(n17), .C(n16), .Y(carry[12]) );
  ADDFHX4 U23 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(n7) );
  NAND3X4 U24 ( .A(n17), .B(n15), .C(n16), .Y(n11) );
  NAND2BX4 U25 ( .AN(n12), .B(carry[24]), .Y(n35) );
  NAND2BX4 U26 ( .AN(n13), .B(n7), .Y(n42) );
  XOR2X1 U27 ( .A(A[11]), .B(B[11]), .Y(n14) );
  XOR2X1 U28 ( .A(n4), .B(n14), .Y(SUM[11]) );
  NAND2X4 U29 ( .A(A[11]), .B(n4), .Y(n15) );
  NAND2X4 U30 ( .A(B[11]), .B(carry[11]), .Y(n16) );
  XOR2XL U31 ( .A(B[12]), .B(A[12]), .Y(n18) );
  XOR2X1 U32 ( .A(n11), .B(n18), .Y(SUM[12]) );
  NAND2X4 U33 ( .A(n11), .B(A[12]), .Y(n20) );
  NAND2XL U34 ( .A(A[12]), .B(B[12]), .Y(n21) );
  XOR2X1 U35 ( .A(A[29]), .B(B[29]), .Y(n22) );
  XOR2X1 U36 ( .A(carry[29]), .B(n22), .Y(SUM[29]) );
  NAND2X4 U37 ( .A(A[29]), .B(n10), .Y(n23) );
  NAND2X4 U38 ( .A(B[29]), .B(n5), .Y(n24) );
  NAND2X4 U39 ( .A(B[29]), .B(A[29]), .Y(n25) );
  NAND3X4 U40 ( .A(n25), .B(n23), .C(n24), .Y(carry[30]) );
  XOR2X1 U41 ( .A(A[19]), .B(B[19]), .Y(n26) );
  XOR2X1 U42 ( .A(carry[19]), .B(n26), .Y(SUM[19]) );
  NAND2X4 U43 ( .A(A[19]), .B(n8), .Y(n27) );
  NAND2X4 U44 ( .A(B[19]), .B(carry[19]), .Y(n28) );
  NAND2X4 U45 ( .A(B[19]), .B(A[19]), .Y(n29) );
  NAND3X4 U46 ( .A(n29), .B(n27), .C(n28), .Y(carry[20]) );
  XOR2X1 U47 ( .A(n3), .B(n30), .Y(SUM[5]) );
  NAND2X4 U48 ( .A(A[5]), .B(carry[5]), .Y(n32) );
  NAND3X4 U49 ( .A(n33), .B(n31), .C(n32), .Y(carry[6]) );
  NAND2X4 U50 ( .A(n2), .B(n36), .Y(carry[25]) );
  NAND2X1 U51 ( .A(B[24]), .B(carry[24]), .Y(n36) );
  XOR2X1 U52 ( .A(A[24]), .B(B[24]), .Y(n34) );
  XOR2X1 U53 ( .A(carry[24]), .B(n34), .Y(SUM[24]) );
  XOR2X1 U54 ( .A(A[31]), .B(B[31]), .Y(n38) );
  NAND2X4 U55 ( .A(n44), .B(n42), .Y(n39) );
  NAND2X4 U56 ( .A(n40), .B(n43), .Y(carry[28]) );
  CLKINVX8 U57 ( .A(n39), .Y(n40) );
  NAND2X4 U58 ( .A(B[27]), .B(A[27]), .Y(n44) );
  XOR2X1 U59 ( .A(A[27]), .B(B[27]), .Y(n41) );
  XOR2X1 U60 ( .A(carry[27]), .B(n41), .Y(SUM[27]) );
  XOR2XL U61 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module hash_core_DW01_add_2 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20;
  wire   [31:2] carry;

  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX4 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX4 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n20), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX4 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX4 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX4 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX4 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX4 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX4 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX4 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX4 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  NAND2BX4 U1 ( .AN(n1), .B(carry[23]), .Y(n17) );
  CLKINVX20 U2 ( .A(A[23]), .Y(n1) );
  AND2X4 U3 ( .A(B[0]), .B(A[0]), .Y(n20) );
  NAND3X4 U4 ( .A(n10), .B(n8), .C(n9), .Y(carry[14]) );
  NAND3X4 U5 ( .A(n14), .B(n12), .C(n13), .Y(carry[28]) );
  NAND2X4 U6 ( .A(n2), .B(n18), .Y(carry[24]) );
  AND2X4 U7 ( .A(n19), .B(n17), .Y(n2) );
  NAND3X2 U8 ( .A(n6), .B(n4), .C(n5), .Y(carry[5]) );
  NAND2X2 U9 ( .A(A[13]), .B(carry[13]), .Y(n9) );
  NAND2X1 U10 ( .A(A[4]), .B(carry[4]), .Y(n5) );
  NAND2X1 U11 ( .A(B[23]), .B(A[23]), .Y(n19) );
  NAND2X1 U12 ( .A(B[27]), .B(A[27]), .Y(n14) );
  NAND2X1 U13 ( .A(A[13]), .B(B[13]), .Y(n10) );
  NAND2X2 U14 ( .A(B[13]), .B(carry[13]), .Y(n8) );
  NAND2X1 U15 ( .A(B[4]), .B(carry[4]), .Y(n4) );
  XOR2X1 U16 ( .A(n15), .B(n16), .Y(SUM[23]) );
  XOR2X1 U17 ( .A(A[23]), .B(B[23]), .Y(n16) );
  XOR2XL U18 ( .A(B[4]), .B(A[4]), .Y(n3) );
  XOR2X1 U19 ( .A(carry[4]), .B(n3), .Y(SUM[4]) );
  NAND2XL U20 ( .A(A[4]), .B(B[4]), .Y(n6) );
  XOR2XL U21 ( .A(B[13]), .B(A[13]), .Y(n7) );
  XOR2X1 U22 ( .A(carry[13]), .B(n7), .Y(SUM[13]) );
  XOR2X1 U23 ( .A(A[27]), .B(B[27]), .Y(n11) );
  XOR2X1 U24 ( .A(carry[27]), .B(n11), .Y(SUM[27]) );
  NAND2X2 U25 ( .A(A[27]), .B(carry[27]), .Y(n12) );
  NAND2X2 U26 ( .A(B[27]), .B(carry[27]), .Y(n13) );
  NAND2X1 U27 ( .A(B[23]), .B(carry[23]), .Y(n18) );
  ADDFHXL U28 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(n15) );
  XOR2XL U29 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module hash_core_DW01_add_4 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  wire   [31:2] carry;

  ADDFHX2 U1_1 ( .A(B[1]), .B(A[1]), .CI(n27), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX4 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX4 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX4 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX4 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX4 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX4 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX4 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX4 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  NAND2X2 U1 ( .A(B[28]), .B(carry[28]), .Y(n13) );
  INVX1 U2 ( .A(B[19]), .Y(n6) );
  NAND2X1 U3 ( .A(B[19]), .B(A[19]), .Y(n26) );
  INVX1 U4 ( .A(B[17]), .Y(n3) );
  INVX1 U5 ( .A(A[17]), .Y(n9) );
  NAND2X1 U6 ( .A(B[17]), .B(A[17]), .Y(n22) );
  INVX1 U7 ( .A(A[19]), .Y(n7) );
  INVX1 U8 ( .A(A[28]), .Y(n4) );
  XOR2X1 U9 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X4 U10 ( .A(n26), .B(n25), .Y(n1) );
  AND2X4 U11 ( .A(n22), .B(n20), .Y(n2) );
  NAND2BX1 U12 ( .AN(n3), .B(carry[17]), .Y(n21) );
  NAND2BX4 U13 ( .AN(n4), .B(n10), .Y(n12) );
  ADDFHX4 U14 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(n5) );
  NAND2BX4 U15 ( .AN(n6), .B(n5), .Y(n25) );
  NAND2BX1 U16 ( .AN(n7), .B(carry[19]), .Y(n24) );
  ADDFHX4 U17 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(n8) );
  NAND2BX4 U18 ( .AN(n9), .B(carry[17]), .Y(n20) );
  ADDFHX4 U19 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(n10) );
  XOR2XL U20 ( .A(A[28]), .B(B[28]), .Y(n11) );
  XOR2X1 U21 ( .A(n10), .B(n11), .Y(SUM[28]) );
  NAND2X4 U22 ( .A(B[28]), .B(A[28]), .Y(n14) );
  NAND3X4 U23 ( .A(n14), .B(n12), .C(n13), .Y(carry[29]) );
  XOR2XL U24 ( .A(A[21]), .B(B[21]), .Y(n15) );
  XOR2X1 U25 ( .A(n8), .B(n15), .Y(SUM[21]) );
  NAND2X4 U26 ( .A(n8), .B(A[21]), .Y(n16) );
  NAND2X4 U27 ( .A(B[21]), .B(carry[21]), .Y(n17) );
  NAND2X4 U28 ( .A(B[21]), .B(A[21]), .Y(n18) );
  NAND3X4 U29 ( .A(n18), .B(n16), .C(n17), .Y(carry[22]) );
  NAND2X4 U30 ( .A(n1), .B(n24), .Y(carry[20]) );
  NAND2X4 U31 ( .A(n2), .B(n21), .Y(carry[18]) );
  XOR2X1 U32 ( .A(A[17]), .B(B[17]), .Y(n19) );
  XOR2X1 U33 ( .A(carry[17]), .B(n19), .Y(SUM[17]) );
  AND2X4 U34 ( .A(B[0]), .B(A[0]), .Y(n27) );
  XOR2X1 U35 ( .A(A[19]), .B(B[19]), .Y(n23) );
  XOR2X1 U36 ( .A(carry[19]), .B(n23), .Y(SUM[19]) );
endmodule


module hash_core_DW01_add_5 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [31:2] carry;

  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n11), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX4 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX4 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX4 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX4 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  NAND3X2 U1 ( .A(n9), .B(n8), .C(n10), .Y(carry[7]) );
  NAND2BX2 U2 ( .AN(n1), .B(carry[6]), .Y(n9) );
  NAND2X2 U3 ( .A(A[6]), .B(carry[6]), .Y(n8) );
  INVX1 U4 ( .A(B[6]), .Y(n1) );
  INVX1 U5 ( .A(A[31]), .Y(n2) );
  XNOR3X4 U6 ( .A(n2), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  XOR2XL U7 ( .A(A[25]), .B(B[25]), .Y(n3) );
  XOR2X1 U8 ( .A(carry[25]), .B(n3), .Y(SUM[25]) );
  NAND2X4 U9 ( .A(A[25]), .B(carry[25]), .Y(n4) );
  NAND2X4 U10 ( .A(B[25]), .B(carry[25]), .Y(n5) );
  NAND2X4 U11 ( .A(B[25]), .B(A[25]), .Y(n6) );
  NAND3X4 U12 ( .A(n6), .B(n4), .C(n5), .Y(carry[26]) );
  AND2X4 U13 ( .A(A[0]), .B(B[0]), .Y(n11) );
  XOR2X1 U14 ( .A(A[6]), .B(B[6]), .Y(n7) );
  XOR2X1 U15 ( .A(carry[6]), .B(n7), .Y(SUM[6]) );
  NAND2XL U16 ( .A(B[6]), .B(A[6]), .Y(n10) );
  XOR2XL U17 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module hash_core_DW01_add_6 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22;
  wire   [31:2] carry;

  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX4 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX4 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .S(SUM[16]) );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX4 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX4 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX4 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  NAND3X4 U1 ( .A(n5), .B(n4), .C(n6), .Y(carry[27]) );
  NAND2X1 U2 ( .A(B[19]), .B(A[19]), .Y(n14) );
  NAND2X1 U3 ( .A(B[10]), .B(A[10]), .Y(n18) );
  NAND2X1 U4 ( .A(A[4]), .B(B[4]), .Y(n10) );
  AND2X2 U5 ( .A(B[0]), .B(A[0]), .Y(n1) );
  ADDFHX4 U6 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(n2) );
  XOR2X1 U7 ( .A(A[26]), .B(B[26]), .Y(n3) );
  XOR2X1 U8 ( .A(carry[26]), .B(n3), .Y(SUM[26]) );
  NAND2X2 U9 ( .A(A[26]), .B(carry[26]), .Y(n4) );
  NAND2X2 U10 ( .A(B[26]), .B(carry[26]), .Y(n5) );
  NAND2XL U11 ( .A(B[26]), .B(A[26]), .Y(n6) );
  XOR2XL U12 ( .A(B[4]), .B(A[4]), .Y(n7) );
  XOR2X1 U13 ( .A(carry[4]), .B(n7), .Y(SUM[4]) );
  NAND2X4 U14 ( .A(B[4]), .B(carry[4]), .Y(n8) );
  NAND2X4 U15 ( .A(A[4]), .B(carry[4]), .Y(n9) );
  NAND3X4 U16 ( .A(n10), .B(n8), .C(n9), .Y(carry[5]) );
  XOR2X1 U17 ( .A(A[19]), .B(B[19]), .Y(n11) );
  XOR2X1 U18 ( .A(carry[19]), .B(n11), .Y(SUM[19]) );
  NAND2X4 U19 ( .A(A[19]), .B(carry[19]), .Y(n12) );
  NAND2X4 U20 ( .A(B[19]), .B(carry[19]), .Y(n13) );
  NAND3X4 U21 ( .A(n14), .B(n12), .C(n13), .Y(carry[20]) );
  XOR2X1 U22 ( .A(A[10]), .B(B[10]), .Y(n15) );
  XOR2X1 U23 ( .A(carry[10]), .B(n15), .Y(SUM[10]) );
  NAND2X4 U24 ( .A(A[10]), .B(carry[10]), .Y(n16) );
  NAND2X4 U25 ( .A(B[10]), .B(carry[10]), .Y(n17) );
  NAND3X4 U26 ( .A(n18), .B(n16), .C(n17), .Y(carry[11]) );
  XOR2X1 U27 ( .A(A[17]), .B(B[17]), .Y(n19) );
  XOR2X1 U28 ( .A(n2), .B(n19), .Y(SUM[17]) );
  NAND2X4 U29 ( .A(A[17]), .B(n2), .Y(n20) );
  NAND2X4 U30 ( .A(B[17]), .B(n2), .Y(n21) );
  NAND2X4 U31 ( .A(B[17]), .B(A[17]), .Y(n22) );
  NAND3X4 U32 ( .A(n22), .B(n20), .C(n21), .Y(carry[18]) );
  XOR2XL U33 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module hash_core_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module hash_core_DW01_add_15 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229;

  OR2X4 U2 ( .A(A[9]), .B(B[9]), .Y(n206) );
  OAI21X4 U3 ( .A0(n68), .A1(n67), .B0(n69), .Y(n5) );
  NAND2X1 U4 ( .A(B[19]), .B(A[19]), .Y(n144) );
  OAI21X4 U5 ( .A0(n68), .A1(n67), .B0(n69), .Y(n56) );
  INVX8 U6 ( .A(n78), .Y(n68) );
  OAI21X2 U7 ( .A0(n95), .A1(n6), .B0(n2), .Y(n93) );
  NAND2X4 U8 ( .A(B[22]), .B(A[22]), .Y(n117) );
  INVX1 U9 ( .A(n192), .Y(n191) );
  OAI21X4 U10 ( .A0(n194), .A1(n16), .B0(n171), .Y(n192) );
  OR2X4 U11 ( .A(A[1]), .B(B[1]), .Y(n73) );
  XOR2X4 U12 ( .A(n93), .B(n94), .Y(SUM[27]) );
  NAND2X2 U13 ( .A(B[10]), .B(A[10]), .Y(n208) );
  NAND2X4 U14 ( .A(B[21]), .B(A[21]), .Y(n116) );
  OR2X4 U15 ( .A(A[21]), .B(B[21]), .Y(n126) );
  INVX4 U16 ( .A(n126), .Y(n114) );
  NOR2BX4 U17 ( .AN(n34), .B(n223), .Y(n219) );
  OAI21X2 U18 ( .A0(n58), .A1(n59), .B0(n60), .Y(n57) );
  NAND2X1 U19 ( .A(A[24]), .B(B[24]), .Y(n88) );
  NOR2X2 U20 ( .A(A[30]), .B(B[30]), .Y(n58) );
  NOR2X2 U21 ( .A(A[30]), .B(B[30]), .Y(n62) );
  INVX1 U22 ( .A(n185), .Y(n176) );
  CLKINVX3 U23 ( .A(n184), .Y(n183) );
  CLKINVX3 U24 ( .A(n160), .Y(n159) );
  NAND2X2 U25 ( .A(B[28]), .B(A[28]), .Y(n69) );
  NAND4BX2 U26 ( .AN(n16), .B(n186), .C(n187), .D(n188), .Y(n178) );
  OR2X2 U27 ( .A(A[20]), .B(B[20]), .Y(n130) );
  AOI21X2 U28 ( .A0(n141), .A1(n142), .B0(n143), .Y(n132) );
  INVX1 U29 ( .A(n144), .Y(n143) );
  CLKINVX3 U30 ( .A(n53), .Y(n7) );
  INVX1 U31 ( .A(n23), .Y(n201) );
  OAI2BB1X2 U32 ( .A0N(n126), .A1N(n127), .B0(n116), .Y(n124) );
  INVX1 U33 ( .A(n3), .Y(n4) );
  OAI21X1 U34 ( .A0(n191), .A1(n174), .B0(n172), .Y(n189) );
  NAND2X1 U35 ( .A(B[13]), .B(A[13]), .Y(n171) );
  XOR2X1 U36 ( .A(n77), .B(n76), .Y(SUM[29]) );
  AOI21X1 U37 ( .A0(n155), .A1(n156), .B0(n157), .Y(n154) );
  CLKINVX3 U38 ( .A(n206), .Y(n22) );
  CLKINVX4 U39 ( .A(n178), .Y(n177) );
  OR2X4 U40 ( .A(A[26]), .B(B[26]), .Y(n91) );
  NOR2BX1 U41 ( .AN(n116), .B(n114), .Y(n128) );
  NAND2X2 U42 ( .A(B[11]), .B(A[11]), .Y(n209) );
  BUFX1 U43 ( .A(n96), .Y(n2) );
  CLKBUFX2 U44 ( .A(n101), .Y(n1) );
  NAND2X1 U45 ( .A(n107), .B(n115), .Y(n127) );
  INVXL U46 ( .A(n104), .Y(n3) );
  XOR2X1 U47 ( .A(n14), .B(n68), .Y(SUM[28]) );
  AOI21X2 U48 ( .A0(n63), .A1(n5), .B0(n65), .Y(n64) );
  INVX4 U49 ( .A(n54), .Y(n8) );
  INVX4 U50 ( .A(n188), .Y(n173) );
  AOI21X2 U51 ( .A0(n176), .A1(n182), .B0(n183), .Y(n180) );
  OAI21X2 U52 ( .A0(n159), .A1(n145), .B0(n147), .Y(n156) );
  NOR2BX1 U53 ( .AN(n2), .B(n6), .Y(n98) );
  NOR2X4 U54 ( .A(B[26]), .B(A[26]), .Y(n6) );
  NAND2X4 U55 ( .A(A[26]), .B(B[26]), .Y(n96) );
  NAND4BBX4 U56 ( .AN(n26), .BN(n22), .C(n205), .D(n204), .Y(n175) );
  NAND2X4 U57 ( .A(n53), .B(n8), .Y(n9) );
  NAND2X2 U58 ( .A(n54), .B(n7), .Y(n10) );
  NAND2X4 U59 ( .A(n9), .B(n10), .Y(SUM[31]) );
  XNOR2X4 U60 ( .A(B[31]), .B(A[31]), .Y(n53) );
  NAND2X2 U61 ( .A(n11), .B(n12), .Y(n13) );
  NAND2X2 U62 ( .A(n13), .B(n181), .Y(n179) );
  INVX2 U63 ( .A(n180), .Y(n11) );
  CLKINVX2 U64 ( .A(n175), .Y(n12) );
  OAI2BB1X4 U65 ( .A0N(n202), .A1N(n203), .B0(n204), .Y(n181) );
  NAND2X4 U66 ( .A(n177), .B(n179), .Y(n164) );
  OAI21X2 U67 ( .A0(n224), .A1(n185), .B0(n184), .Y(n23) );
  OAI2BB1X4 U68 ( .A0N(n219), .A1N(n220), .B0(n31), .Y(n184) );
  XOR2X4 U69 ( .A(n121), .B(n122), .Y(SUM[23]) );
  OAI21X2 U70 ( .A0(n123), .A1(n118), .B0(n117), .Y(n121) );
  OAI21X1 U71 ( .A0(n201), .A1(n175), .B0(n181), .Y(n199) );
  AOI21X1 U72 ( .A0(n78), .A1(n70), .B0(n79), .Y(n77) );
  INVX2 U73 ( .A(n195), .Y(n194) );
  NAND2X4 U74 ( .A(B[9]), .B(A[9]), .Y(n21) );
  NAND4BBX2 U75 ( .AN(n39), .BN(n17), .C(n37), .D(n31), .Y(n185) );
  NAND2X4 U76 ( .A(B[7]), .B(A[7]), .Y(n29) );
  OR2X4 U77 ( .A(A[7]), .B(B[7]), .Y(n31) );
  NOR2X4 U78 ( .A(n138), .B(n137), .Y(n141) );
  NAND2X2 U79 ( .A(B[12]), .B(A[12]), .Y(n170) );
  OR2X4 U80 ( .A(A[11]), .B(B[11]), .Y(n204) );
  OR2X1 U81 ( .A(A[12]), .B(B[12]), .Y(n186) );
  OR2XL U82 ( .A(A[2]), .B(B[2]), .Y(n72) );
  NAND2X1 U83 ( .A(B[2]), .B(A[2]), .Y(n51) );
  AOI21XL U84 ( .A0(n205), .A1(n213), .B0(n214), .Y(n212) );
  NAND2X1 U85 ( .A(B[24]), .B(A[24]), .Y(n103) );
  NOR2X1 U86 ( .A(A[4]), .B(B[4]), .Y(n17) );
  NAND2XL U87 ( .A(n218), .B(n25), .Y(n19) );
  NAND2X1 U88 ( .A(B[17]), .B(A[17]), .Y(n147) );
  NAND2X2 U89 ( .A(B[14]), .B(A[14]), .Y(n172) );
  NAND2X2 U90 ( .A(B[27]), .B(A[27]), .Y(n86) );
  AOI21X4 U91 ( .A0(n83), .A1(n84), .B0(n85), .Y(n82) );
  NAND3X1 U92 ( .A(n205), .B(n206), .C(n207), .Y(n203) );
  INVX1 U93 ( .A(n210), .Y(n26) );
  NAND2XL U94 ( .A(n139), .B(n140), .Y(n134) );
  OAI21XL U95 ( .A0(n151), .A1(n152), .B0(n75), .Y(n229) );
  OAI21XL U96 ( .A0(n38), .A1(n39), .B0(n40), .Y(n35) );
  OAI211X2 U97 ( .A0(n16), .A1(n170), .B0(n171), .C0(n172), .Y(n167) );
  NAND2X2 U98 ( .A(n162), .B(n146), .Y(n160) );
  NAND2XL U99 ( .A(n69), .B(n70), .Y(n14) );
  NAND2X4 U100 ( .A(n99), .B(n89), .Y(n97) );
  NAND3XL U101 ( .A(n221), .B(n37), .C(n222), .Y(n220) );
  OAI21X2 U102 ( .A0(n197), .A1(n198), .B0(n170), .Y(n195) );
  INVX2 U103 ( .A(n199), .Y(n198) );
  AND2X2 U104 ( .A(n208), .B(n209), .Y(n202) );
  OAI21X2 U105 ( .A0(n226), .A1(n227), .B0(n47), .Y(n182) );
  NOR2BXL U106 ( .AN(n170), .B(n197), .Y(n200) );
  AND2X1 U107 ( .A(n103), .B(n105), .Y(n106) );
  NOR2BXL U108 ( .AN(n171), .B(n16), .Y(n196) );
  NOR2BXL U109 ( .AN(n21), .B(n22), .Y(n20) );
  AND2X1 U110 ( .A(n89), .B(n100), .Y(n102) );
  AND2X1 U111 ( .A(n113), .B(n120), .Y(n122) );
  INVXL U112 ( .A(n37), .Y(n33) );
  AND2X1 U113 ( .A(n146), .B(n139), .Y(n163) );
  AND2X1 U114 ( .A(n115), .B(n130), .Y(n131) );
  NOR2BXL U115 ( .AN(n40), .B(n39), .Y(n42) );
  INVXL U116 ( .A(n225), .Y(n48) );
  NOR2BXL U117 ( .AN(n75), .B(n151), .Y(n150) );
  INVXL U118 ( .A(n152), .Y(n74) );
  XOR2X1 U119 ( .A(B[30]), .B(A[30]), .Y(n18) );
  NAND2X2 U120 ( .A(B[18]), .B(A[18]), .Y(n148) );
  NAND2XL U121 ( .A(B[5]), .B(A[5]), .Y(n40) );
  NAND2XL U122 ( .A(B[1]), .B(A[1]), .Y(n75) );
  NAND2XL U123 ( .A(B[3]), .B(A[3]), .Y(n47) );
  NAND2X2 U124 ( .A(B[16]), .B(A[16]), .Y(n146) );
  NOR2BX1 U125 ( .AN(n152), .B(n15), .Y(SUM[0]) );
  NOR2XL U126 ( .A(A[0]), .B(B[0]), .Y(n15) );
  INVX1 U127 ( .A(n182), .Y(n224) );
  INVX1 U128 ( .A(n69), .Y(n79) );
  INVXL U129 ( .A(n119), .Y(n118) );
  INVX1 U130 ( .A(n221), .Y(n39) );
  INVX1 U131 ( .A(n186), .Y(n197) );
  NOR2BX1 U132 ( .AN(n117), .B(n118), .Y(n125) );
  INVX1 U133 ( .A(n124), .Y(n123) );
  NOR2BXL U134 ( .AN(n86), .B(n90), .Y(n94) );
  INVX1 U135 ( .A(n86), .Y(n85) );
  NAND2X1 U136 ( .A(n40), .B(n43), .Y(n222) );
  NAND2XL U137 ( .A(n63), .B(n66), .Y(n76) );
  XOR2X1 U138 ( .A(n156), .B(n158), .Y(SUM[18]) );
  NOR2BXL U139 ( .AN(n148), .B(n137), .Y(n158) );
  XOR2X1 U140 ( .A(n192), .B(n193), .Y(SUM[14]) );
  NOR2BXL U141 ( .AN(n172), .B(n174), .Y(n193) );
  XOR2X1 U142 ( .A(n153), .B(n154), .Y(SUM[19]) );
  NAND2XL U143 ( .A(n144), .B(n149), .Y(n153) );
  INVX1 U144 ( .A(n148), .Y(n157) );
  XOR2X1 U145 ( .A(n160), .B(n161), .Y(SUM[17]) );
  NOR2BXL U146 ( .AN(n147), .B(n145), .Y(n161) );
  NAND2X1 U147 ( .A(n21), .B(n25), .Y(n207) );
  INVX1 U148 ( .A(n29), .Y(n223) );
  XOR2X1 U149 ( .A(n1), .B(n102), .Y(SUM[25]) );
  XOR2X1 U150 ( .A(n97), .B(n98), .Y(SUM[26]) );
  XOR2X1 U151 ( .A(n127), .B(n128), .Y(SUM[21]) );
  XOR2X1 U152 ( .A(n129), .B(n131), .Y(SUM[20]) );
  XOR2X1 U153 ( .A(n124), .B(n125), .Y(SUM[22]) );
  OAI21XL U154 ( .A0(n217), .A1(n22), .B0(n21), .Y(n213) );
  INVX1 U155 ( .A(n19), .Y(n217) );
  NOR2X1 U156 ( .A(n228), .B(n229), .Y(n226) );
  NAND2X1 U157 ( .A(n72), .B(n225), .Y(n227) );
  INVX1 U158 ( .A(n51), .Y(n228) );
  INVX1 U159 ( .A(n208), .Y(n214) );
  INVX1 U160 ( .A(n73), .Y(n151) );
  NAND2X1 U161 ( .A(n23), .B(n210), .Y(n218) );
  XOR2X1 U162 ( .A(n199), .B(n200), .Y(SUM[12]) );
  XOR2X1 U163 ( .A(n213), .B(n215), .Y(SUM[10]) );
  NOR2BX1 U164 ( .AN(n208), .B(n216), .Y(n215) );
  INVX1 U165 ( .A(n205), .Y(n216) );
  XOR2X1 U166 ( .A(n19), .B(n20), .Y(SUM[9]) );
  OAI21XL U167 ( .A0(n17), .A1(n224), .B0(n43), .Y(n41) );
  INVX1 U168 ( .A(n41), .Y(n38) );
  XOR2X1 U169 ( .A(n23), .B(n24), .Y(SUM[8]) );
  NOR2BX1 U170 ( .AN(n25), .B(n26), .Y(n24) );
  XOR2X1 U171 ( .A(n41), .B(n42), .Y(SUM[5]) );
  XOR2X1 U172 ( .A(n35), .B(n36), .Y(SUM[6]) );
  NOR2BX1 U173 ( .AN(n34), .B(n33), .Y(n36) );
  INVX1 U174 ( .A(n31), .Y(n30) );
  XOR2X1 U175 ( .A(n27), .B(n28), .Y(SUM[7]) );
  OAI21XL U176 ( .A0(n32), .A1(n33), .B0(n34), .Y(n27) );
  NOR2BX1 U177 ( .AN(n29), .B(n30), .Y(n28) );
  INVX1 U178 ( .A(n35), .Y(n32) );
  NAND2X1 U179 ( .A(n204), .B(n209), .Y(n211) );
  INVX1 U180 ( .A(n72), .Y(n50) );
  XOR2X1 U181 ( .A(n52), .B(n71), .Y(SUM[2]) );
  NOR2BX1 U182 ( .AN(n51), .B(n50), .Y(n71) );
  OAI2BB1X1 U183 ( .A0N(n73), .A1N(n74), .B0(n75), .Y(n52) );
  XOR2X1 U184 ( .A(n182), .B(n44), .Y(SUM[4]) );
  NOR2BX1 U185 ( .AN(n43), .B(n17), .Y(n44) );
  XOR2X1 U186 ( .A(n45), .B(n46), .Y(SUM[3]) );
  OAI21XL U187 ( .A0(n49), .A1(n50), .B0(n51), .Y(n45) );
  NOR2BX1 U188 ( .AN(n47), .B(n48), .Y(n46) );
  INVX1 U189 ( .A(n52), .Y(n49) );
  XOR2X1 U190 ( .A(n74), .B(n150), .Y(SUM[1]) );
  NOR2X2 U191 ( .A(A[13]), .B(B[13]), .Y(n16) );
  NAND2X1 U192 ( .A(B[8]), .B(A[8]), .Y(n25) );
  XNOR2X4 U193 ( .A(n64), .B(n18), .Y(SUM[30]) );
  NAND2X1 U194 ( .A(B[6]), .B(A[6]), .Y(n34) );
  OR2X2 U195 ( .A(A[6]), .B(B[6]), .Y(n37) );
  OR2X2 U196 ( .A(A[16]), .B(B[16]), .Y(n139) );
  OR2X2 U197 ( .A(A[24]), .B(B[24]), .Y(n105) );
  OR2X2 U198 ( .A(A[8]), .B(B[8]), .Y(n210) );
  NAND2X2 U199 ( .A(B[30]), .B(A[30]), .Y(n60) );
  OR2X2 U200 ( .A(A[5]), .B(B[5]), .Y(n221) );
  NAND2X1 U201 ( .A(B[4]), .B(A[4]), .Y(n43) );
  OR2X2 U202 ( .A(A[3]), .B(B[3]), .Y(n225) );
  XOR2X1 U203 ( .A(n211), .B(n212), .Y(SUM[11]) );
  XOR2X1 U204 ( .A(n195), .B(n196), .Y(SUM[13]) );
  NAND2X1 U205 ( .A(B[0]), .B(A[0]), .Y(n152) );
  NAND2X4 U206 ( .A(n164), .B(n165), .Y(n135) );
  OR2XL U207 ( .A(A[25]), .B(B[25]), .Y(n100) );
  NAND2X1 U208 ( .A(B[23]), .B(A[23]), .Y(n113) );
  NAND2X2 U209 ( .A(B[29]), .B(A[29]), .Y(n66) );
  NAND2XL U210 ( .A(A[29]), .B(B[29]), .Y(n59) );
  NAND2XL U211 ( .A(n135), .B(n139), .Y(n162) );
  XOR2X1 U212 ( .A(n135), .B(n163), .Y(SUM[16]) );
  INVX4 U213 ( .A(n97), .Y(n95) );
  INVX8 U214 ( .A(n92), .Y(n90) );
  XOR2X1 U215 ( .A(n189), .B(n190), .Y(SUM[15]) );
  NOR2BXL U216 ( .AN(n169), .B(n173), .Y(n190) );
  INVX8 U217 ( .A(n155), .Y(n137) );
  INVX4 U218 ( .A(n149), .Y(n138) );
  NAND3BX2 U219 ( .AN(n87), .B(n91), .C(n92), .Y(n81) );
  AND2X4 U220 ( .A(n120), .B(n119), .Y(n110) );
  NAND3BX2 U221 ( .AN(n114), .B(n120), .C(n119), .Y(n108) );
  XOR2X1 U222 ( .A(n4), .B(n106), .Y(SUM[24]) );
  NAND2XL U223 ( .A(B[15]), .B(A[15]), .Y(n169) );
  AOI21X4 U224 ( .A0(n56), .A1(n55), .B0(n57), .Y(n54) );
  NOR2X4 U225 ( .A(n61), .B(n62), .Y(n55) );
  CLKINVX3 U226 ( .A(n63), .Y(n61) );
  CLKINVX3 U227 ( .A(n66), .Y(n65) );
  CLKINVX3 U228 ( .A(n70), .Y(n67) );
  OR2X4 U229 ( .A(A[29]), .B(B[29]), .Y(n63) );
  OAI21X4 U230 ( .A0(n80), .A1(n81), .B0(n82), .Y(n78) );
  OAI211X2 U231 ( .A0(n87), .A1(n88), .B0(n96), .C0(n89), .Y(n84) );
  NOR2X4 U232 ( .A(A[25]), .B(B[25]), .Y(n87) );
  NOR2X4 U233 ( .A(n90), .B(n6), .Y(n83) );
  OR2X4 U234 ( .A(A[28]), .B(B[28]), .Y(n70) );
  OR2X4 U235 ( .A(A[27]), .B(B[27]), .Y(n92) );
  NAND2X4 U236 ( .A(n100), .B(n101), .Y(n99) );
  NAND2X4 U237 ( .A(B[25]), .B(A[25]), .Y(n89) );
  NAND2X4 U238 ( .A(n80), .B(n103), .Y(n101) );
  NAND2X4 U239 ( .A(n104), .B(n105), .Y(n80) );
  OAI21X4 U240 ( .A0(n107), .A1(n108), .B0(n109), .Y(n104) );
  AOI21X4 U241 ( .A0(n110), .A1(n111), .B0(n112), .Y(n109) );
  CLKINVX3 U242 ( .A(n113), .Y(n112) );
  OAI211X2 U243 ( .A0(n114), .A1(n115), .B0(n116), .C0(n117), .Y(n111) );
  OR2X4 U244 ( .A(A[23]), .B(B[23]), .Y(n120) );
  OR2X4 U245 ( .A(A[22]), .B(B[22]), .Y(n119) );
  NAND2X4 U246 ( .A(n129), .B(n130), .Y(n107) );
  NAND2X4 U247 ( .A(B[20]), .B(A[20]), .Y(n115) );
  NAND2X4 U248 ( .A(n132), .B(n133), .Y(n129) );
  NAND3BX4 U249 ( .AN(n134), .B(n135), .C(n136), .Y(n133) );
  NOR2X4 U250 ( .A(n137), .B(n138), .Y(n136) );
  OAI211X2 U251 ( .A0(n145), .A1(n146), .B0(n147), .C0(n148), .Y(n142) );
  OR2X4 U252 ( .A(A[19]), .B(B[19]), .Y(n149) );
  OR2X4 U253 ( .A(A[18]), .B(B[18]), .Y(n155) );
  CLKINVX3 U254 ( .A(n140), .Y(n145) );
  OR2X4 U255 ( .A(A[17]), .B(B[17]), .Y(n140) );
  AOI21X4 U256 ( .A0(n166), .A1(n167), .B0(n168), .Y(n165) );
  CLKINVX3 U257 ( .A(n169), .Y(n168) );
  NOR2X4 U258 ( .A(n173), .B(n174), .Y(n166) );
  OR2X4 U259 ( .A(A[15]), .B(B[15]), .Y(n188) );
  CLKINVX3 U260 ( .A(n187), .Y(n174) );
  OR2X4 U261 ( .A(A[14]), .B(B[14]), .Y(n187) );
  OR2X4 U262 ( .A(A[10]), .B(B[10]), .Y(n205) );
endmodule


module hash_core_DW01_add_16 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228;

  XOR2X1 U2 ( .A(n126), .B(n127), .Y(SUM[22]) );
  CLKINVX4 U3 ( .A(n126), .Y(n125) );
  NOR2BX2 U4 ( .AN(n32), .B(n222), .Y(n218) );
  NOR2X4 U5 ( .A(n59), .B(n60), .Y(n53) );
  CLKINVX8 U6 ( .A(n61), .Y(n59) );
  NOR2X2 U7 ( .A(A[25]), .B(B[25]), .Y(n86) );
  NOR2BX1 U8 ( .AN(n118), .B(n120), .Y(n127) );
  INVX4 U9 ( .A(n121), .Y(n120) );
  XOR2X2 U10 ( .A(A[30]), .B(B[30]), .Y(n15) );
  NAND2X4 U11 ( .A(B[30]), .B(A[30]), .Y(n58) );
  NOR2X4 U12 ( .A(A[30]), .B(B[30]), .Y(n60) );
  INVXL U13 ( .A(n118), .Y(n4) );
  OR2X4 U14 ( .A(A[25]), .B(B[25]), .Y(n101) );
  INVX3 U15 ( .A(n52), .Y(n6) );
  NAND2X4 U16 ( .A(B[26]), .B(A[26]), .Y(n97) );
  NAND2X2 U17 ( .A(B[21]), .B(A[21]), .Y(n117) );
  INVX8 U18 ( .A(n128), .Y(n115) );
  OR2X4 U19 ( .A(A[21]), .B(B[21]), .Y(n128) );
  OAI21X1 U20 ( .A0(n200), .A1(n177), .B0(n182), .Y(n198) );
  CLKINVX3 U21 ( .A(n21), .Y(n200) );
  NAND2X4 U22 ( .A(B[11]), .B(A[11]), .Y(n208) );
  OAI2BB1X4 U23 ( .A0N(n128), .A1N(n129), .B0(n117), .Y(n126) );
  NOR2X2 U24 ( .A(n66), .B(n65), .Y(n9) );
  INVX4 U25 ( .A(n183), .Y(n223) );
  OAI21X4 U26 ( .A0(n225), .A1(n226), .B0(n45), .Y(n183) );
  OAI211X2 U27 ( .A0(n115), .A1(n116), .B0(n117), .C0(n118), .Y(n112) );
  AOI21X2 U28 ( .A0(n178), .A1(n183), .B0(n184), .Y(n181) );
  INVXL U29 ( .A(n173), .Y(n12) );
  INVXL U30 ( .A(n13), .Y(n11) );
  NOR2X2 U31 ( .A(n9), .B(n77), .Y(n75) );
  OAI2BB1X2 U32 ( .A0N(n201), .A1N(n202), .B0(n203), .Y(n182) );
  NAND4BBX2 U33 ( .AN(n24), .BN(n20), .C(n204), .D(n203), .Y(n177) );
  OAI21X2 U34 ( .A0(n56), .A1(n57), .B0(n58), .Y(n55) );
  NAND2X1 U35 ( .A(A[24]), .B(B[24]), .Y(n87) );
  OR2X2 U36 ( .A(A[22]), .B(B[22]), .Y(n121) );
  NOR2X2 U37 ( .A(A[13]), .B(B[13]), .Y(n13) );
  NAND2X1 U38 ( .A(B[13]), .B(A[13]), .Y(n173) );
  NAND2X1 U39 ( .A(B[8]), .B(A[8]), .Y(n23) );
  CLKINVX3 U40 ( .A(n93), .Y(n89) );
  INVX2 U41 ( .A(n101), .Y(n91) );
  NAND2X2 U42 ( .A(B[25]), .B(A[25]), .Y(n88) );
  NAND2X1 U43 ( .A(B[22]), .B(A[22]), .Y(n118) );
  INVX1 U44 ( .A(n10), .Y(n192) );
  CLKINVX3 U45 ( .A(n162), .Y(n161) );
  NAND2X2 U46 ( .A(B[20]), .B(A[20]), .Y(n116) );
  AOI21X2 U47 ( .A0(n143), .A1(n144), .B0(n145), .Y(n134) );
  NAND2X1 U48 ( .A(n108), .B(n116), .Y(n129) );
  XNOR2X2 U49 ( .A(n62), .B(n15), .Y(SUM[30]) );
  INVX1 U50 ( .A(n64), .Y(n63) );
  OR2X2 U51 ( .A(A[28]), .B(B[28]), .Y(n68) );
  OAI21X4 U52 ( .A0(n181), .A1(n177), .B0(n182), .Y(n180) );
  NAND2X1 U53 ( .A(B[17]), .B(A[17]), .Y(n149) );
  AOI21X1 U54 ( .A0(n194), .A1(n11), .B0(n12), .Y(n10) );
  OAI21X2 U55 ( .A0(n196), .A1(n197), .B0(n172), .Y(n194) );
  NAND2X2 U56 ( .A(B[9]), .B(A[9]), .Y(n19) );
  NAND2X1 U57 ( .A(B[29]), .B(A[29]), .Y(n57) );
  NOR2X4 U58 ( .A(B[30]), .B(A[30]), .Y(n56) );
  OAI21X2 U59 ( .A0(n161), .A1(n147), .B0(n149), .Y(n158) );
  INVXL U60 ( .A(n105), .Y(n1) );
  INVX2 U61 ( .A(n1), .Y(n2) );
  INVX4 U62 ( .A(n142), .Y(n147) );
  INVX2 U63 ( .A(n114), .Y(n113) );
  XOR2X1 U64 ( .A(n78), .B(n66), .Y(SUM[28]) );
  NAND2X1 U65 ( .A(n67), .B(n68), .Y(n78) );
  CLKINVX8 U66 ( .A(n92), .Y(n90) );
  NAND2XL U67 ( .A(n137), .B(n141), .Y(n164) );
  NAND2X1 U68 ( .A(n141), .B(n142), .Y(n136) );
  CLKINVX2 U69 ( .A(n185), .Y(n184) );
  INVX3 U70 ( .A(n189), .Y(n175) );
  NOR2X4 U71 ( .A(n125), .B(n120), .Y(n3) );
  OR2X4 U72 ( .A(n3), .B(n4), .Y(n123) );
  XOR2X4 U73 ( .A(n123), .B(n124), .Y(SUM[23]) );
  NAND2X4 U74 ( .A(n51), .B(n6), .Y(n7) );
  NAND2X4 U75 ( .A(n5), .B(n52), .Y(n8) );
  NAND2X4 U76 ( .A(n7), .B(n8), .Y(SUM[31]) );
  INVX4 U77 ( .A(n51), .Y(n5) );
  INVX2 U78 ( .A(n67), .Y(n77) );
  XOR2X4 U79 ( .A(n74), .B(n75), .Y(SUM[29]) );
  AOI21X2 U80 ( .A0(n61), .A1(n54), .B0(n63), .Y(n62) );
  NAND2X2 U81 ( .A(n100), .B(n88), .Y(n98) );
  NOR2BX2 U82 ( .AN(n88), .B(n91), .Y(n103) );
  XNOR2X4 U83 ( .A(B[31]), .B(A[31]), .Y(n51) );
  NAND2X2 U84 ( .A(n79), .B(n104), .Y(n102) );
  NAND2X2 U85 ( .A(B[19]), .B(A[19]), .Y(n146) );
  OR2XL U86 ( .A(A[8]), .B(B[8]), .Y(n209) );
  OR2XL U87 ( .A(A[2]), .B(B[2]), .Y(n70) );
  NAND2X1 U88 ( .A(B[2]), .B(A[2]), .Y(n49) );
  AOI21X1 U89 ( .A0(n157), .A1(n158), .B0(n159), .Y(n156) );
  NAND3X1 U90 ( .A(n204), .B(n205), .C(n206), .Y(n202) );
  NAND2X1 U91 ( .A(B[7]), .B(A[7]), .Y(n27) );
  OR2X2 U92 ( .A(A[7]), .B(B[7]), .Y(n29) );
  NOR2XL U93 ( .A(A[4]), .B(B[4]), .Y(n14) );
  XOR2X1 U94 ( .A(n98), .B(n99), .Y(SUM[26]) );
  NAND4BBX2 U95 ( .AN(n37), .BN(n14), .C(n35), .D(n29), .Y(n186) );
  OAI21X2 U96 ( .A0(n10), .A1(n176), .B0(n174), .Y(n190) );
  NOR2BX1 U97 ( .AN(n172), .B(n196), .Y(n199) );
  OAI21XL U98 ( .A0(n153), .A1(n154), .B0(n73), .Y(n228) );
  OAI21XL U99 ( .A0(n36), .A1(n37), .B0(n38), .Y(n33) );
  NAND2X1 U100 ( .A(B[29]), .B(A[29]), .Y(n64) );
  NAND2XL U101 ( .A(B[24]), .B(A[24]), .Y(n104) );
  NAND2X2 U102 ( .A(B[14]), .B(A[14]), .Y(n174) );
  NAND2X2 U103 ( .A(B[10]), .B(A[10]), .Y(n207) );
  OR2X2 U104 ( .A(A[24]), .B(B[24]), .Y(n106) );
  OR2X2 U105 ( .A(A[5]), .B(B[5]), .Y(n220) );
  INVX2 U106 ( .A(n198), .Y(n197) );
  NAND2X2 U107 ( .A(n164), .B(n148), .Y(n162) );
  INVXL U108 ( .A(n150), .Y(n159) );
  AND2X2 U109 ( .A(n207), .B(n208), .Y(n201) );
  OAI21X4 U110 ( .A0(n96), .A1(n90), .B0(n97), .Y(n94) );
  INVX4 U111 ( .A(n98), .Y(n96) );
  NAND4BX2 U112 ( .AN(n13), .B(n187), .C(n188), .D(n189), .Y(n179) );
  NOR2BXL U113 ( .AN(n19), .B(n20), .Y(n18) );
  AND2X1 U114 ( .A(n148), .B(n141), .Y(n165) );
  NOR2BXL U115 ( .AN(n23), .B(n24), .Y(n22) );
  INVXL U116 ( .A(n35), .Y(n31) );
  AND2X1 U117 ( .A(n116), .B(n132), .Y(n133) );
  INVXL U118 ( .A(n224), .Y(n46) );
  NOR2BXL U119 ( .AN(n73), .B(n153), .Y(n152) );
  INVXL U120 ( .A(n154), .Y(n72) );
  NAND2X2 U121 ( .A(B[5]), .B(A[5]), .Y(n38) );
  OR2X4 U122 ( .A(A[9]), .B(B[9]), .Y(n205) );
  NAND2X2 U123 ( .A(B[12]), .B(A[12]), .Y(n172) );
  NAND2XL U124 ( .A(B[1]), .B(A[1]), .Y(n73) );
  NAND2XL U125 ( .A(B[3]), .B(A[3]), .Y(n45) );
  NAND2X2 U126 ( .A(B[27]), .B(A[27]), .Y(n85) );
  OR2XL U127 ( .A(A[12]), .B(B[12]), .Y(n187) );
  OR2X4 U128 ( .A(A[16]), .B(B[16]), .Y(n141) );
  NOR2XL U129 ( .A(A[0]), .B(B[0]), .Y(n16) );
  OAI21X4 U130 ( .A0(n223), .A1(n186), .B0(n185), .Y(n21) );
  OAI2BB1X4 U131 ( .A0N(n218), .A1N(n219), .B0(n29), .Y(n185) );
  INVX1 U132 ( .A(n186), .Y(n178) );
  OAI211X1 U133 ( .A0(n13), .A1(n172), .B0(n173), .C0(n174), .Y(n169) );
  NOR2BXL U134 ( .AN(n97), .B(n90), .Y(n99) );
  INVX1 U135 ( .A(n85), .Y(n84) );
  INVX1 U136 ( .A(n205), .Y(n20) );
  INVX1 U137 ( .A(n220), .Y(n37) );
  NOR2BXL U138 ( .AN(n114), .B(n119), .Y(n124) );
  NOR2BXL U139 ( .AN(n117), .B(n115), .Y(n130) );
  INVX1 U140 ( .A(n146), .Y(n145) );
  INVX1 U141 ( .A(n209), .Y(n24) );
  NAND3X1 U142 ( .A(n220), .B(n35), .C(n221), .Y(n219) );
  NAND2X1 U143 ( .A(n38), .B(n41), .Y(n221) );
  XOR2X1 U144 ( .A(n102), .B(n103), .Y(SUM[25]) );
  XOR2X1 U145 ( .A(n190), .B(n191), .Y(SUM[15]) );
  XOR2X1 U146 ( .A(n192), .B(n193), .Y(SUM[14]) );
  NOR2BXL U147 ( .AN(n174), .B(n176), .Y(n193) );
  NAND2XL U148 ( .A(n61), .B(n64), .Y(n74) );
  XOR2X1 U149 ( .A(n155), .B(n156), .Y(SUM[19]) );
  NAND2XL U150 ( .A(n146), .B(n151), .Y(n155) );
  NAND2X1 U151 ( .A(n19), .B(n23), .Y(n206) );
  NAND2X2 U152 ( .A(n101), .B(n102), .Y(n100) );
  INVX1 U153 ( .A(n27), .Y(n222) );
  AND2X2 U154 ( .A(n104), .B(n106), .Y(n107) );
  XOR2X1 U155 ( .A(n158), .B(n160), .Y(SUM[18]) );
  XOR2X1 U156 ( .A(n129), .B(n130), .Y(SUM[21]) );
  XOR2X1 U157 ( .A(n131), .B(n133), .Y(SUM[20]) );
  XOR2X1 U158 ( .A(n162), .B(n163), .Y(SUM[17]) );
  OAI21XL U159 ( .A0(n216), .A1(n20), .B0(n19), .Y(n212) );
  INVX1 U160 ( .A(n17), .Y(n216) );
  NOR2X1 U161 ( .A(n227), .B(n228), .Y(n225) );
  NAND2X1 U162 ( .A(n70), .B(n224), .Y(n226) );
  INVX1 U163 ( .A(n49), .Y(n227) );
  AOI21XL U164 ( .A0(n204), .A1(n212), .B0(n213), .Y(n211) );
  INVX1 U165 ( .A(n207), .Y(n213) );
  INVX1 U166 ( .A(n187), .Y(n196) );
  INVX1 U167 ( .A(n71), .Y(n153) );
  NOR2BXL U168 ( .AN(n149), .B(n147), .Y(n163) );
  NOR2BXL U169 ( .AN(n150), .B(n139), .Y(n160) );
  NAND2X1 U170 ( .A(n217), .B(n23), .Y(n17) );
  NAND2X1 U171 ( .A(n21), .B(n209), .Y(n217) );
  XOR2X1 U172 ( .A(n212), .B(n214), .Y(SUM[10]) );
  NOR2BX1 U173 ( .AN(n207), .B(n215), .Y(n214) );
  INVXL U174 ( .A(n204), .Y(n215) );
  XOR2X1 U175 ( .A(n198), .B(n199), .Y(SUM[12]) );
  XOR2X1 U176 ( .A(n194), .B(n195), .Y(SUM[13]) );
  NOR2BX1 U177 ( .AN(n173), .B(n13), .Y(n195) );
  XOR2X1 U178 ( .A(n17), .B(n18), .Y(SUM[9]) );
  NAND2XL U179 ( .A(n203), .B(n208), .Y(n210) );
  XOR2X1 U180 ( .A(n210), .B(n211), .Y(SUM[11]) );
  NOR2BX1 U181 ( .AN(n154), .B(n16), .Y(SUM[0]) );
  OAI21XL U182 ( .A0(n14), .A1(n223), .B0(n41), .Y(n39) );
  INVX1 U183 ( .A(n39), .Y(n36) );
  XOR2X1 U184 ( .A(n39), .B(n40), .Y(SUM[5]) );
  NOR2BX1 U185 ( .AN(n38), .B(n37), .Y(n40) );
  XOR2X1 U186 ( .A(n33), .B(n34), .Y(SUM[6]) );
  NOR2BX1 U187 ( .AN(n32), .B(n31), .Y(n34) );
  INVX1 U188 ( .A(n29), .Y(n28) );
  XOR2X1 U189 ( .A(n21), .B(n22), .Y(SUM[8]) );
  XOR2X1 U190 ( .A(n25), .B(n26), .Y(SUM[7]) );
  OAI21XL U191 ( .A0(n30), .A1(n31), .B0(n32), .Y(n25) );
  NOR2BX1 U192 ( .AN(n27), .B(n28), .Y(n26) );
  INVX1 U193 ( .A(n33), .Y(n30) );
  INVX1 U194 ( .A(n70), .Y(n48) );
  XOR2X1 U195 ( .A(n50), .B(n69), .Y(SUM[2]) );
  NOR2BX1 U196 ( .AN(n49), .B(n48), .Y(n69) );
  OAI2BB1X1 U197 ( .A0N(n71), .A1N(n72), .B0(n73), .Y(n50) );
  XOR2X1 U198 ( .A(n183), .B(n42), .Y(SUM[4]) );
  NOR2BX1 U199 ( .AN(n41), .B(n14), .Y(n42) );
  XOR2X1 U200 ( .A(n43), .B(n44), .Y(SUM[3]) );
  OAI21XL U201 ( .A0(n47), .A1(n48), .B0(n49), .Y(n43) );
  NOR2BX1 U202 ( .AN(n45), .B(n46), .Y(n44) );
  INVX1 U203 ( .A(n50), .Y(n47) );
  XOR2X1 U204 ( .A(n72), .B(n152), .Y(SUM[1]) );
  NAND2X2 U205 ( .A(B[28]), .B(A[28]), .Y(n67) );
  NAND2X1 U206 ( .A(B[6]), .B(A[6]), .Y(n32) );
  OR2X2 U207 ( .A(A[6]), .B(B[6]), .Y(n35) );
  NAND2X2 U208 ( .A(B[18]), .B(A[18]), .Y(n150) );
  OR2X2 U209 ( .A(A[20]), .B(B[20]), .Y(n132) );
  NAND2X1 U210 ( .A(B[4]), .B(A[4]), .Y(n41) );
  OR2X2 U211 ( .A(A[3]), .B(B[3]), .Y(n224) );
  OR2X2 U212 ( .A(A[1]), .B(B[1]), .Y(n71) );
  NAND2X1 U213 ( .A(B[0]), .B(A[0]), .Y(n154) );
  NAND2X4 U214 ( .A(n166), .B(n167), .Y(n137) );
  NAND2X1 U215 ( .A(B[23]), .B(A[23]), .Y(n114) );
  NAND3BX2 U216 ( .AN(n91), .B(n92), .C(n93), .Y(n80) );
  XOR2X1 U217 ( .A(n137), .B(n165), .Y(SUM[16]) );
  INVX8 U218 ( .A(n76), .Y(n66) );
  NAND2XL U219 ( .A(B[15]), .B(A[15]), .Y(n171) );
  NOR2BXL U220 ( .AN(n171), .B(n175), .Y(n191) );
  INVX8 U221 ( .A(n157), .Y(n139) );
  NAND3BX2 U222 ( .AN(n115), .B(n121), .C(n122), .Y(n109) );
  NOR2BXL U223 ( .AN(n85), .B(n89), .Y(n95) );
  INVX8 U224 ( .A(n122), .Y(n119) );
  INVX8 U225 ( .A(n151), .Y(n140) );
  XOR2X1 U226 ( .A(n2), .B(n107), .Y(SUM[24]) );
  AOI21X4 U227 ( .A0(n54), .A1(n53), .B0(n55), .Y(n52) );
  OAI21X4 U228 ( .A0(n65), .A1(n66), .B0(n67), .Y(n54) );
  CLKINVX3 U229 ( .A(n68), .Y(n65) );
  OR2X4 U230 ( .A(A[29]), .B(B[29]), .Y(n61) );
  OAI21X4 U231 ( .A0(n79), .A1(n80), .B0(n81), .Y(n76) );
  AOI21X4 U232 ( .A0(n82), .A1(n83), .B0(n84), .Y(n81) );
  OAI211X2 U233 ( .A0(n86), .A1(n87), .B0(n88), .C0(n97), .Y(n83) );
  NOR2X4 U234 ( .A(n89), .B(n90), .Y(n82) );
  XOR2X4 U235 ( .A(n94), .B(n95), .Y(SUM[27]) );
  OR2X4 U236 ( .A(A[27]), .B(B[27]), .Y(n93) );
  OR2X4 U237 ( .A(A[26]), .B(B[26]), .Y(n92) );
  NAND2X4 U238 ( .A(n105), .B(n106), .Y(n79) );
  OAI21X4 U239 ( .A0(n108), .A1(n109), .B0(n110), .Y(n105) );
  AOI21X4 U240 ( .A0(n111), .A1(n112), .B0(n113), .Y(n110) );
  NOR2X4 U241 ( .A(n119), .B(n120), .Y(n111) );
  OR2X4 U242 ( .A(A[23]), .B(B[23]), .Y(n122) );
  NAND2X4 U243 ( .A(n131), .B(n132), .Y(n108) );
  NAND2X4 U244 ( .A(n134), .B(n135), .Y(n131) );
  NAND3BX4 U245 ( .AN(n136), .B(n137), .C(n138), .Y(n135) );
  NOR2X4 U246 ( .A(n139), .B(n140), .Y(n138) );
  OAI211X2 U247 ( .A0(n147), .A1(n148), .B0(n149), .C0(n150), .Y(n144) );
  NOR2X4 U248 ( .A(n140), .B(n139), .Y(n143) );
  OR2X4 U249 ( .A(A[19]), .B(B[19]), .Y(n151) );
  OR2X4 U250 ( .A(A[18]), .B(B[18]), .Y(n157) );
  OR2X4 U251 ( .A(A[17]), .B(B[17]), .Y(n142) );
  NAND2X4 U252 ( .A(B[16]), .B(A[16]), .Y(n148) );
  AOI21X4 U253 ( .A0(n168), .A1(n169), .B0(n170), .Y(n167) );
  CLKINVX3 U254 ( .A(n171), .Y(n170) );
  NOR2X4 U255 ( .A(n175), .B(n176), .Y(n168) );
  NAND2BX4 U256 ( .AN(n179), .B(n180), .Y(n166) );
  OR2X4 U257 ( .A(A[15]), .B(B[15]), .Y(n189) );
  CLKINVX3 U258 ( .A(n188), .Y(n176) );
  OR2X4 U259 ( .A(A[14]), .B(B[14]), .Y(n188) );
  OR2X4 U260 ( .A(A[11]), .B(B[11]), .Y(n203) );
  OR2X4 U261 ( .A(A[10]), .B(B[10]), .Y(n204) );
endmodule


module hash_core_DW01_add_20 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209;

  OAI21X1 U2 ( .A0(n59), .A1(n60), .B0(n61), .Y(n57) );
  AOI21X1 U3 ( .A0(n69), .A1(n70), .B0(n71), .Y(n60) );
  XOR2X2 U4 ( .A(n138), .B(n139), .Y(SUM[19]) );
  OAI21X2 U5 ( .A0(n177), .A1(n10), .B0(n161), .Y(n175) );
  NAND3XL U6 ( .A(A[0]), .B(B[0]), .C(n65), .Y(n64) );
  OAI2BB1X2 U7 ( .A0N(B[0]), .A1N(A[0]), .B0(n66), .Y(n207) );
  NAND2X4 U8 ( .A(n119), .B(n120), .Y(n99) );
  OAI21X2 U9 ( .A0(n123), .A1(n124), .B0(n125), .Y(n119) );
  OR2X2 U10 ( .A(A[18]), .B(B[18]), .Y(n135) );
  NAND2X1 U11 ( .A(n21), .B(n192), .Y(n191) );
  OAI21XL U12 ( .A0(n154), .A1(n12), .B0(n155), .Y(n153) );
  INVX1 U13 ( .A(n159), .Y(n158) );
  OAI21XL U14 ( .A0(n10), .A1(n160), .B0(n161), .Y(n157) );
  NAND2X1 U15 ( .A(n95), .B(n96), .Y(n75) );
  INVX2 U16 ( .A(n19), .Y(n200) );
  OAI21X2 U17 ( .A0(n183), .A1(n162), .B0(n184), .Y(n181) );
  NAND2X1 U18 ( .A(B[4]), .B(A[4]), .Y(n40) );
  INVX1 U19 ( .A(n204), .Y(n31) );
  XOR2X2 U20 ( .A(n173), .B(n174), .Y(SUM[15]) );
  XOR2X1 U21 ( .A(n175), .B(n176), .Y(SUM[14]) );
  OAI21XL U22 ( .A0(n51), .A1(n52), .B0(n53), .Y(n47) );
  NAND2X1 U23 ( .A(n92), .B(n87), .Y(n90) );
  NAND2X1 U24 ( .A(n76), .B(n93), .Y(n92) );
  NAND2X2 U25 ( .A(n40), .B(n35), .Y(n205) );
  OAI2BB1X4 U26 ( .A0N(n8), .A1N(n39), .B0(n169), .Y(n23) );
  NAND2X4 U27 ( .A(n146), .B(n147), .Y(n123) );
  INVX4 U28 ( .A(n23), .Y(n183) );
  OAI21X4 U29 ( .A0(n200), .A1(n22), .B0(n21), .Y(n196) );
  NOR2X4 U30 ( .A(A[13]), .B(B[13]), .Y(n10) );
  NAND2XL U31 ( .A(B[13]), .B(A[13]), .Y(n161) );
  NAND3BX2 U32 ( .AN(n172), .B(n49), .C(n171), .Y(n39) );
  OAI21X4 U33 ( .A0(n185), .A1(n186), .B0(n187), .Y(n167) );
  XNOR2X1 U34 ( .A(n114), .B(n7), .Y(SUM[22]) );
  XNOR2X1 U35 ( .A(n57), .B(n4), .Y(SUM[30]) );
  NOR2X2 U36 ( .A(n166), .B(n167), .Y(n150) );
  XOR2X1 U37 ( .A(n63), .B(n51), .Y(SUM[2]) );
  NAND3BXL U38 ( .AN(n14), .B(n135), .C(n136), .Y(n124) );
  NOR2BX1 U39 ( .AN(n40), .B(n46), .Y(n45) );
  NOR2BXL U40 ( .AN(n28), .B(n29), .Y(n27) );
  XOR2X1 U41 ( .A(n26), .B(n27), .Y(SUM[7]) );
  AND2X2 U42 ( .A(n83), .B(n78), .Y(n9) );
  NAND3XL U43 ( .A(n37), .B(n204), .C(n205), .Y(n202) );
  NOR2BX1 U44 ( .AN(n49), .B(n172), .Y(n170) );
  INVX1 U45 ( .A(n83), .Y(n91) );
  AOI21XL U46 ( .A0(n78), .A1(n90), .B0(n91), .Y(n89) );
  NAND4BXL U47 ( .AN(n11), .B(n193), .C(n188), .D(n189), .Y(n162) );
  NAND2X1 U48 ( .A(B[2]), .B(A[2]), .Y(n53) );
  OR2X2 U49 ( .A(A[1]), .B(B[1]), .Y(n65) );
  NAND2X1 U50 ( .A(B[6]), .B(A[6]), .Y(n32) );
  OR2X2 U51 ( .A(A[5]), .B(B[5]), .Y(n37) );
  OR2X2 U52 ( .A(A[17]), .B(B[17]), .Y(n136) );
  AND2X2 U53 ( .A(n1), .B(n2), .Y(n8) );
  NOR2X1 U54 ( .A(n41), .B(n46), .Y(n1) );
  NOR2X1 U55 ( .A(n29), .B(n31), .Y(n2) );
  OAI21X4 U56 ( .A0(n150), .A1(n151), .B0(n152), .Y(n146) );
  NAND2XL U57 ( .A(n53), .B(n67), .Y(n63) );
  NAND3X1 U58 ( .A(n3), .B(n35), .C(n36), .Y(n33) );
  OR2XL U59 ( .A(n40), .B(n41), .Y(n3) );
  XOR2X2 U60 ( .A(n88), .B(n89), .Y(SUM[27]) );
  XOR2X2 U61 ( .A(n90), .B(n9), .Y(SUM[26]) );
  NOR2BX1 U62 ( .AN(n134), .B(n126), .Y(n125) );
  OAI21X1 U63 ( .A0(n13), .A1(n180), .B0(n160), .Y(n178) );
  NAND2X1 U64 ( .A(n55), .B(n58), .Y(n4) );
  NOR2BXL U65 ( .AN(n159), .B(n165), .Y(n176) );
  INVX2 U66 ( .A(n193), .Y(n22) );
  AND2X2 U67 ( .A(n32), .B(n28), .Y(n201) );
  NAND2BXL U68 ( .AN(n53), .B(n208), .Y(n209) );
  XNOR2X1 U69 ( .A(n95), .B(n5), .Y(SUM[24]) );
  NAND2X1 U70 ( .A(n86), .B(n96), .Y(n5) );
  XNOR2X1 U71 ( .A(n69), .B(n6), .Y(SUM[28]) );
  NAND2X1 U72 ( .A(n72), .B(n70), .Y(n6) );
  NAND2X1 U73 ( .A(n107), .B(n102), .Y(n7) );
  INVXL U74 ( .A(n189), .Y(n199) );
  AOI21XL U75 ( .A0(n102), .A1(n114), .B0(n115), .Y(n113) );
  NOR2BXL U76 ( .AN(n128), .B(n129), .Y(n142) );
  XOR2XL U77 ( .A(n68), .B(n60), .Y(SUM[29]) );
  NOR2BXL U78 ( .AN(n134), .B(n14), .Y(n139) );
  NOR2BXL U79 ( .AN(n21), .B(n22), .Y(n20) );
  NAND2XL U80 ( .A(n99), .B(n110), .Y(n117) );
  NAND2XL U81 ( .A(n123), .B(n132), .Y(n144) );
  NAND2XL U82 ( .A(n57), .B(n58), .Y(n56) );
  NOR2XL U83 ( .A(A[0]), .B(B[0]), .Y(n16) );
  AND2X1 U84 ( .A(B[0]), .B(A[0]), .Y(n17) );
  NAND2X2 U85 ( .A(B[1]), .B(A[1]), .Y(n66) );
  NAND2XL U86 ( .A(B[0]), .B(A[0]), .Y(n18) );
  NAND2XL U87 ( .A(B[9]), .B(A[9]), .Y(n21) );
  NAND2XL U88 ( .A(B[7]), .B(A[7]), .Y(n28) );
  NOR2XL U89 ( .A(A[12]), .B(B[12]), .Y(n13) );
  NOR2XL U90 ( .A(A[8]), .B(B[8]), .Y(n11) );
  NAND2XL U91 ( .A(B[11]), .B(A[11]), .Y(n187) );
  NAND2XL U92 ( .A(B[15]), .B(A[15]), .Y(n155) );
  NAND2XL U93 ( .A(B[19]), .B(A[19]), .Y(n134) );
  OR2XL U94 ( .A(A[16]), .B(B[16]), .Y(n147) );
  INVX1 U95 ( .A(n167), .Y(n184) );
  NAND2X1 U96 ( .A(n163), .B(n164), .Y(n151) );
  INVX1 U97 ( .A(n153), .Y(n152) );
  OAI21XL U98 ( .A0(n11), .A1(n183), .B0(n25), .Y(n19) );
  NOR2BX1 U99 ( .AN(n155), .B(n12), .Y(n174) );
  OAI2BB1X1 U100 ( .A0N(n156), .A1N(n175), .B0(n159), .Y(n173) );
  INVX1 U101 ( .A(n67), .Y(n52) );
  INVX1 U102 ( .A(n208), .Y(n50) );
  XOR2X1 U103 ( .A(n194), .B(n195), .Y(SUM[11]) );
  NAND2X1 U104 ( .A(n187), .B(n188), .Y(n194) );
  AOI21X1 U105 ( .A0(n189), .A1(n196), .B0(n197), .Y(n195) );
  INVX1 U106 ( .A(n192), .Y(n197) );
  INVX1 U107 ( .A(n178), .Y(n177) );
  INVX1 U108 ( .A(n181), .Y(n180) );
  NAND2X1 U109 ( .A(n188), .B(n189), .Y(n186) );
  NOR2X1 U110 ( .A(n190), .B(n191), .Y(n185) );
  NAND3X1 U111 ( .A(n37), .B(n38), .C(n39), .Y(n36) );
  INVX1 U112 ( .A(n37), .Y(n41) );
  INVX1 U113 ( .A(n38), .Y(n46) );
  INVX1 U114 ( .A(n203), .Y(n29) );
  XOR2X1 U115 ( .A(n39), .B(n45), .Y(SUM[4]) );
  XOR2X1 U116 ( .A(n196), .B(n198), .Y(SUM[10]) );
  NOR2BX1 U117 ( .AN(n192), .B(n199), .Y(n198) );
  XOR2X1 U118 ( .A(n181), .B(n182), .Y(SUM[12]) );
  NOR2BX1 U119 ( .AN(n160), .B(n13), .Y(n182) );
  XOR2X1 U120 ( .A(n33), .B(n34), .Y(SUM[6]) );
  NOR2BX1 U121 ( .AN(n32), .B(n31), .Y(n34) );
  XOR2X1 U122 ( .A(n47), .B(n48), .Y(SUM[3]) );
  NOR2BX1 U123 ( .AN(n49), .B(n50), .Y(n48) );
  XOR2X1 U124 ( .A(n42), .B(n43), .Y(SUM[5]) );
  NAND2X1 U125 ( .A(n37), .B(n35), .Y(n42) );
  AOI21X1 U126 ( .A0(n39), .A1(n38), .B0(n44), .Y(n43) );
  INVX1 U127 ( .A(n40), .Y(n44) );
  XOR2X1 U128 ( .A(n23), .B(n24), .Y(SUM[8]) );
  NOR2BX1 U129 ( .AN(n25), .B(n11), .Y(n24) );
  AOI21X1 U130 ( .A0(n168), .A1(n169), .B0(n162), .Y(n166) );
  OAI2BB1X1 U131 ( .A0N(n170), .A1N(n171), .B0(n8), .Y(n168) );
  AOI21X1 U132 ( .A0(n156), .A1(n157), .B0(n158), .Y(n154) );
  NAND2X1 U133 ( .A(n116), .B(n111), .Y(n114) );
  NAND2X1 U134 ( .A(n100), .B(n117), .Y(n116) );
  OAI2BB1X1 U135 ( .A0N(n201), .A1N(n202), .B0(n203), .Y(n169) );
  NOR2X1 U136 ( .A(n22), .B(n25), .Y(n190) );
  NAND2X1 U137 ( .A(n143), .B(n133), .Y(n141) );
  NAND2X1 U138 ( .A(n136), .B(n144), .Y(n143) );
  XOR2X1 U139 ( .A(n178), .B(n179), .Y(SUM[13]) );
  NOR2BX1 U140 ( .AN(n161), .B(n10), .Y(n179) );
  XOR2X1 U141 ( .A(n141), .B(n142), .Y(SUM[18]) );
  OAI21XL U142 ( .A0(n140), .A1(n129), .B0(n128), .Y(n138) );
  INVX1 U143 ( .A(n141), .Y(n140) );
  XOR2X1 U144 ( .A(n19), .B(n20), .Y(SUM[9]) );
  OAI21XL U145 ( .A0(n30), .A1(n31), .B0(n32), .Y(n26) );
  INVX1 U146 ( .A(n33), .Y(n30) );
  NAND2X1 U147 ( .A(n66), .B(n65), .Y(n137) );
  INVX1 U148 ( .A(n209), .Y(n172) );
  INVX1 U149 ( .A(n72), .Y(n71) );
  NAND2X1 U150 ( .A(n81), .B(n77), .Y(n88) );
  INVX1 U151 ( .A(n62), .Y(n59) );
  INVX1 U152 ( .A(n135), .Y(n129) );
  XOR2X1 U153 ( .A(n119), .B(n121), .Y(SUM[20]) );
  NOR2BX1 U154 ( .AN(n110), .B(n122), .Y(n121) );
  INVX1 U155 ( .A(n120), .Y(n122) );
  INVX1 U156 ( .A(n136), .Y(n131) );
  XOR2X1 U157 ( .A(n117), .B(n118), .Y(SUM[21]) );
  NOR2BX1 U158 ( .AN(n111), .B(n109), .Y(n118) );
  INVX1 U159 ( .A(n156), .Y(n165) );
  AOI21X1 U160 ( .A0(n127), .A1(n128), .B0(n14), .Y(n126) );
  NAND2BX1 U161 ( .AN(n129), .B(n130), .Y(n127) );
  OAI21XL U162 ( .A0(n131), .A1(n132), .B0(n133), .Y(n130) );
  XOR2X1 U163 ( .A(n146), .B(n148), .Y(SUM[16]) );
  NOR2BX1 U164 ( .AN(n132), .B(n149), .Y(n148) );
  INVX1 U165 ( .A(n147), .Y(n149) );
  NAND2X1 U166 ( .A(n97), .B(n98), .Y(n95) );
  AOI21X1 U167 ( .A0(n103), .A1(n101), .B0(n104), .Y(n97) );
  NAND4BXL U168 ( .AN(n99), .B(n100), .C(n101), .D(n102), .Y(n98) );
  INVX1 U169 ( .A(n105), .Y(n104) );
  XOR2X1 U170 ( .A(n144), .B(n145), .Y(SUM[17]) );
  NOR2BX1 U171 ( .AN(n133), .B(n131), .Y(n145) );
  NAND2X1 U172 ( .A(n61), .B(n62), .Y(n68) );
  XOR2X1 U173 ( .A(n112), .B(n113), .Y(SUM[23]) );
  NAND2X1 U174 ( .A(n105), .B(n101), .Y(n112) );
  INVX1 U175 ( .A(n107), .Y(n115) );
  NAND2X1 U176 ( .A(n75), .B(n86), .Y(n93) );
  NAND2X1 U177 ( .A(n73), .B(n74), .Y(n69) );
  AOI21X1 U178 ( .A0(n79), .A1(n77), .B0(n80), .Y(n73) );
  NAND4BXL U179 ( .AN(n75), .B(n76), .C(n77), .D(n78), .Y(n74) );
  INVX1 U180 ( .A(n81), .Y(n80) );
  NOR2X1 U181 ( .A(n10), .B(n13), .Y(n163) );
  XOR2X1 U182 ( .A(n93), .B(n94), .Y(SUM[25]) );
  NOR2BX1 U183 ( .AN(n87), .B(n85), .Y(n94) );
  NOR2X1 U184 ( .A(n12), .B(n165), .Y(n164) );
  INVX1 U185 ( .A(n100), .Y(n109) );
  NAND2X1 U186 ( .A(n106), .B(n107), .Y(n103) );
  NAND2X1 U187 ( .A(n102), .B(n108), .Y(n106) );
  OAI21XL U188 ( .A0(n109), .A1(n110), .B0(n111), .Y(n108) );
  NAND2X1 U189 ( .A(n55), .B(n56), .Y(n54) );
  INVX1 U190 ( .A(n76), .Y(n85) );
  NAND2X1 U191 ( .A(n82), .B(n83), .Y(n79) );
  NAND2X1 U192 ( .A(n78), .B(n84), .Y(n82) );
  OAI21XL U193 ( .A0(n85), .A1(n86), .B0(n87), .Y(n84) );
  NAND3X1 U194 ( .A(n206), .B(n65), .C(n207), .Y(n171) );
  NOR2X1 U195 ( .A(n50), .B(n52), .Y(n206) );
  OR2X2 U196 ( .A(A[3]), .B(B[3]), .Y(n208) );
  OR2X2 U197 ( .A(A[2]), .B(B[2]), .Y(n67) );
  XOR3X2 U198 ( .A(B[31]), .B(A[31]), .C(n54), .Y(SUM[31]) );
  AND2X2 U199 ( .A(n66), .B(n64), .Y(n51) );
  OR2X2 U200 ( .A(A[10]), .B(B[10]), .Y(n189) );
  NAND2X1 U201 ( .A(B[5]), .B(A[5]), .Y(n35) );
  NAND2X1 U202 ( .A(B[8]), .B(A[8]), .Y(n25) );
  OR2X2 U203 ( .A(A[11]), .B(B[11]), .Y(n188) );
  NAND2X1 U204 ( .A(B[10]), .B(A[10]), .Y(n192) );
  NAND2X1 U205 ( .A(B[3]), .B(A[3]), .Y(n49) );
  OR2X2 U206 ( .A(A[4]), .B(B[4]), .Y(n38) );
  XOR2X1 U207 ( .A(n18), .B(n137), .Y(SUM[1]) );
  OR2X2 U208 ( .A(A[9]), .B(B[9]), .Y(n193) );
  OR2X2 U209 ( .A(A[6]), .B(B[6]), .Y(n204) );
  OR2X2 U210 ( .A(A[7]), .B(B[7]), .Y(n203) );
  NOR2X1 U211 ( .A(A[15]), .B(B[15]), .Y(n12) );
  NOR2X1 U212 ( .A(A[19]), .B(B[19]), .Y(n14) );
  NAND2X1 U213 ( .A(B[12]), .B(A[12]), .Y(n160) );
  NAND2X1 U214 ( .A(B[17]), .B(A[17]), .Y(n133) );
  NAND2X1 U215 ( .A(B[14]), .B(A[14]), .Y(n159) );
  NOR2X1 U216 ( .A(n16), .B(n17), .Y(SUM[0]) );
  OR2X2 U217 ( .A(A[14]), .B(B[14]), .Y(n156) );
  OR2X2 U218 ( .A(A[22]), .B(B[22]), .Y(n102) );
  NAND2X1 U219 ( .A(B[22]), .B(A[22]), .Y(n107) );
  NAND2X1 U220 ( .A(B[16]), .B(A[16]), .Y(n132) );
  NAND2X1 U221 ( .A(B[20]), .B(A[20]), .Y(n110) );
  NAND2X1 U222 ( .A(B[18]), .B(A[18]), .Y(n128) );
  OR2X2 U223 ( .A(A[23]), .B(B[23]), .Y(n101) );
  NAND2X1 U224 ( .A(B[21]), .B(A[21]), .Y(n111) );
  OR2X2 U225 ( .A(A[21]), .B(B[21]), .Y(n100) );
  OR2X2 U226 ( .A(A[20]), .B(B[20]), .Y(n120) );
  OR2X2 U227 ( .A(A[26]), .B(B[26]), .Y(n78) );
  NAND2X1 U228 ( .A(B[24]), .B(A[24]), .Y(n86) );
  NAND2X1 U229 ( .A(B[26]), .B(A[26]), .Y(n83) );
  OR2X2 U230 ( .A(A[27]), .B(B[27]), .Y(n77) );
  NAND2X1 U231 ( .A(B[25]), .B(A[25]), .Y(n87) );
  OR2X2 U232 ( .A(A[25]), .B(B[25]), .Y(n76) );
  NAND2X1 U233 ( .A(B[23]), .B(A[23]), .Y(n105) );
  NAND2X1 U234 ( .A(B[27]), .B(A[27]), .Y(n81) );
  OR2X2 U235 ( .A(A[28]), .B(B[28]), .Y(n70) );
  OR2X2 U236 ( .A(A[24]), .B(B[24]), .Y(n96) );
  NAND2X1 U237 ( .A(B[30]), .B(A[30]), .Y(n55) );
  NAND2X1 U238 ( .A(B[29]), .B(A[29]), .Y(n61) );
  NAND2X1 U239 ( .A(B[28]), .B(A[28]), .Y(n72) );
  OR2X2 U240 ( .A(A[30]), .B(B[30]), .Y(n58) );
  OR2X2 U241 ( .A(A[29]), .B(B[29]), .Y(n62) );
endmodule


module hash_core_DW01_add_19 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n333, n334, n335, n336, n337, n1, n2, n4, n6, n7, n8, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332;

  NAND2X4 U2 ( .A(B[1]), .B(A[1]), .Y(n133) );
  CLKBUFX8 U3 ( .A(n139), .Y(n4) );
  NAND2BX4 U4 ( .AN(n1), .B(n311), .Y(n280) );
  NAND2X2 U5 ( .A(n309), .B(n310), .Y(n1) );
  NAND2X2 U6 ( .A(n94), .B(n95), .Y(n93) );
  INVXL U7 ( .A(n291), .Y(n321) );
  AND2X4 U8 ( .A(n281), .B(n282), .Y(n2) );
  NOR2X4 U9 ( .A(n2), .B(n283), .Y(n278) );
  CLKINVX2 U10 ( .A(n284), .Y(n283) );
  XOR2X2 U11 ( .A(n224), .B(n267), .Y(n336) );
  NOR2BX4 U12 ( .AN(n21), .B(n6), .Y(n323) );
  CLKBUFX8 U13 ( .A(n321), .Y(n6) );
  XOR2X2 U14 ( .A(n151), .B(n152), .Y(n333) );
  NAND2X4 U15 ( .A(n12), .B(n245), .Y(n272) );
  NAND2X2 U16 ( .A(B[26]), .B(A[26]), .Y(n155) );
  NAND4BX2 U17 ( .AN(n46), .B(n290), .C(n75), .D(n67), .Y(n325) );
  NOR2X2 U18 ( .A(n144), .B(n145), .Y(n161) );
  BUFX12 U19 ( .A(n45), .Y(SUM[14]) );
  AOI21X2 U20 ( .A0(n118), .A1(n119), .B0(n120), .Y(n117) );
  NAND3X4 U21 ( .A(n50), .B(n122), .C(n123), .Y(n118) );
  NAND3BX2 U22 ( .AN(n249), .B(n250), .C(n242), .Y(n248) );
  OAI21X1 U23 ( .A0(n144), .A1(n149), .B0(n150), .Y(n146) );
  NAND2X4 U24 ( .A(B[22]), .B(A[22]), .Y(n170) );
  NAND2BX4 U25 ( .AN(n102), .B(n90), .Y(n94) );
  NAND2X2 U26 ( .A(n90), .B(n95), .Y(n103) );
  INVX4 U27 ( .A(n90), .Y(n73) );
  NAND2X2 U28 ( .A(n91), .B(n90), .Y(n329) );
  NAND3BX1 U29 ( .AN(n262), .B(n242), .C(n263), .Y(n260) );
  NAND2X2 U30 ( .A(n138), .B(n4), .Y(n43) );
  OAI21X4 U31 ( .A0(n11), .A1(n146), .B0(n147), .Y(n138) );
  INVX8 U32 ( .A(n156), .Y(n144) );
  BUFX20 U33 ( .A(n335), .Y(SUM[21]) );
  NAND3BX2 U34 ( .AN(n96), .B(n98), .C(n97), .Y(n105) );
  INVX8 U35 ( .A(n285), .Y(n96) );
  BUFX12 U36 ( .A(n333), .Y(SUM[27]) );
  NOR2X2 U37 ( .A(n56), .B(n143), .Y(n147) );
  AOI21X4 U38 ( .A0(n238), .A1(n239), .B0(n240), .Y(n235) );
  OAI21X1 U39 ( .A0(n251), .A1(n252), .B0(n253), .Y(n250) );
  NAND2X1 U40 ( .A(B[14]), .B(A[14]), .Y(n293) );
  NOR2XL U41 ( .A(A[14]), .B(B[14]), .Y(n22) );
  OAI2BB1X2 U42 ( .A0N(n247), .A1N(n248), .B0(n210), .Y(n246) );
  NOR2X2 U43 ( .A(n225), .B(n226), .Y(n222) );
  INVX8 U44 ( .A(n238), .Y(n226) );
  NAND2X2 U45 ( .A(n15), .B(n242), .Y(n239) );
  NOR2X1 U46 ( .A(n196), .B(n195), .Y(n198) );
  INVX4 U47 ( .A(n185), .Y(n196) );
  INVX4 U48 ( .A(B[24]), .Y(n7) );
  CLKINVX8 U49 ( .A(n7), .Y(n8) );
  XOR2X4 U50 ( .A(n71), .B(n107), .Y(SUM[4]) );
  NOR2BX2 U51 ( .AN(n229), .B(n226), .Y(n267) );
  NAND2BX2 U52 ( .AN(n229), .B(n230), .Y(n209) );
  OR2X4 U53 ( .A(A[17]), .B(B[17]), .Y(n230) );
  BUFX8 U54 ( .A(n336), .Y(SUM[16]) );
  NAND2X4 U55 ( .A(B[8]), .B(A[8]), .Y(n64) );
  INVX8 U56 ( .A(n184), .Y(n195) );
  AOI21X4 U57 ( .A0(n91), .A1(n92), .B0(n93), .Y(n88) );
  NAND2X2 U58 ( .A(B[2]), .B(A[2]), .Y(n114) );
  INVX1 U59 ( .A(n53), .Y(n30) );
  NAND2BX2 U60 ( .AN(n187), .B(n185), .Y(n168) );
  NAND2X2 U61 ( .A(n184), .B(n214), .Y(n35) );
  NAND2BX2 U62 ( .AN(n215), .B(n202), .Y(n214) );
  INVX4 U63 ( .A(n302), .Y(n275) );
  INVX2 U64 ( .A(n323), .Y(n24) );
  NAND2X1 U65 ( .A(n256), .B(n302), .Y(n312) );
  INVX2 U66 ( .A(n111), .Y(n110) );
  NAND2X2 U67 ( .A(n115), .B(n27), .Y(n28) );
  INVX2 U68 ( .A(n129), .Y(n27) );
  XOR2X2 U69 ( .A(n116), .B(n117), .Y(SUM[31]) );
  NAND2X2 U70 ( .A(n156), .B(n148), .Y(n154) );
  CLKINVX3 U71 ( .A(n286), .Y(n281) );
  INVX4 U72 ( .A(n148), .Y(n143) );
  NAND2BX2 U73 ( .AN(n256), .B(n287), .Y(n264) );
  OAI21XL U74 ( .A0(A[9]), .A1(B[9]), .B0(n290), .Y(n327) );
  BUFX3 U75 ( .A(n310), .Y(n21) );
  NOR2X1 U76 ( .A(n292), .B(n275), .Y(n308) );
  NOR2X2 U77 ( .A(n68), .B(n69), .Y(n66) );
  NAND3BX2 U78 ( .AN(n70), .B(n71), .C(n72), .Y(n63) );
  NOR3X2 U79 ( .A(n69), .B(n73), .C(n74), .Y(n72) );
  NAND2X1 U80 ( .A(B[9]), .B(A[9]), .Y(n61) );
  AND2X2 U81 ( .A(n263), .B(n241), .Y(n15) );
  NAND2X1 U82 ( .A(B[18]), .B(A[18]), .Y(n237) );
  NAND2X2 U83 ( .A(B[17]), .B(A[17]), .Y(n210) );
  CLKINVX3 U84 ( .A(n230), .Y(n225) );
  NAND2X1 U85 ( .A(n229), .B(n263), .Y(n249) );
  OAI21XL U86 ( .A0(n255), .A1(n256), .B0(n257), .Y(n251) );
  INVX4 U87 ( .A(n173), .Y(n179) );
  NAND2X2 U88 ( .A(n10), .B(n165), .Y(n176) );
  NAND2X1 U89 ( .A(n178), .B(n172), .Y(n177) );
  INVX4 U90 ( .A(n157), .Y(n145) );
  INVX1 U91 ( .A(n150), .Y(n163) );
  OAI21X1 U92 ( .A0(n256), .A1(n255), .B0(n257), .Y(n299) );
  OR2X2 U93 ( .A(A[3]), .B(B[3]), .Y(n111) );
  NOR2BX2 U94 ( .AN(n114), .B(n113), .Y(n129) );
  OR2X2 U95 ( .A(A[1]), .B(B[1]), .Y(n131) );
  NAND3X2 U96 ( .A(n124), .B(n125), .C(n126), .Y(n123) );
  INVX1 U97 ( .A(n125), .Y(n128) );
  NAND2X1 U98 ( .A(B[27]), .B(A[27]), .Y(n139) );
  NAND2X1 U99 ( .A(n150), .B(n149), .Y(n158) );
  BUFX3 U100 ( .A(n337), .Y(SUM[0]) );
  NOR2BX2 U101 ( .AN(n263), .B(n276), .Y(n295) );
  INVX1 U102 ( .A(n263), .Y(n270) );
  OAI21XL U103 ( .A0(A[13]), .A1(B[13]), .B0(n302), .Y(n301) );
  AND2X2 U104 ( .A(n177), .B(n167), .Y(n10) );
  AND2X2 U105 ( .A(B[26]), .B(A[26]), .Y(n11) );
  INVX1 U106 ( .A(n187), .Y(n193) );
  AND2X2 U107 ( .A(n288), .B(n287), .Y(n12) );
  AND2X2 U108 ( .A(n207), .B(n237), .Y(n13) );
  AND2X2 U109 ( .A(n206), .B(n208), .Y(n14) );
  NOR2X4 U110 ( .A(n62), .B(n69), .Y(n316) );
  NAND2X1 U111 ( .A(n207), .B(n208), .Y(n204) );
  BUFX8 U112 ( .A(n183), .Y(n16) );
  NAND2XL U113 ( .A(n230), .B(n210), .Y(n258) );
  NAND3BX4 U114 ( .AN(n329), .B(n71), .C(n330), .Y(n17) );
  NAND3BX2 U115 ( .AN(n329), .B(n71), .C(n330), .Y(n80) );
  BUFX3 U116 ( .A(A[15]), .Y(n18) );
  NAND2X1 U117 ( .A(n210), .B(n229), .Y(n240) );
  AND3X4 U118 ( .A(n309), .B(n313), .C(n300), .Y(n48) );
  CLKINVX2 U119 ( .A(n300), .Y(n305) );
  INVX3 U120 ( .A(n296), .Y(n31) );
  NAND2X1 U121 ( .A(n308), .B(n280), .Y(n307) );
  INVX2 U122 ( .A(n280), .Y(n279) );
  XOR2X2 U123 ( .A(n86), .B(n87), .Y(SUM[7]) );
  NOR3X4 U124 ( .A(n188), .B(n195), .C(n196), .Y(n194) );
  NAND2X2 U125 ( .A(B[14]), .B(A[14]), .Y(n254) );
  NOR2BX2 U126 ( .AN(n98), .B(n110), .Y(n109) );
  OAI2BB1X2 U127 ( .A0N(n227), .A1N(n217), .B0(n206), .Y(n221) );
  BUFX3 U128 ( .A(A[23]), .Y(n19) );
  NAND2X4 U129 ( .A(B[12]), .B(A[12]), .Y(n256) );
  OAI21X4 U130 ( .A0(n320), .A1(n6), .B0(n21), .Y(n318) );
  AND2X2 U131 ( .A(n172), .B(n185), .Y(n57) );
  NOR4BBX4 U132 ( .AN(n280), .BN(n20), .C(n275), .D(n292), .Y(n298) );
  OR2XL U133 ( .A(A[13]), .B(B[13]), .Y(n20) );
  NAND2X2 U134 ( .A(B[13]), .B(A[13]), .Y(n257) );
  CLKINVX3 U135 ( .A(n287), .Y(n255) );
  NAND3BX4 U136 ( .AN(n243), .B(n244), .C(n245), .Y(n241) );
  OAI21X4 U137 ( .A0(n193), .A1(n183), .B0(n194), .Y(n192) );
  NAND2X2 U138 ( .A(n320), .B(n323), .Y(n26) );
  NAND3BX2 U139 ( .AN(n164), .B(n165), .C(n166), .Y(n162) );
  NAND2X2 U140 ( .A(B[15]), .B(n18), .Y(n263) );
  NAND2X2 U141 ( .A(n322), .B(n24), .Y(n25) );
  NOR2BX4 U142 ( .AN(n76), .B(n68), .Y(n330) );
  AOI2BB1X4 U143 ( .A0N(n17), .A1N(n327), .B0(n328), .Y(n324) );
  OAI21X4 U144 ( .A0(n62), .A1(n64), .B0(n61), .Y(n328) );
  INVX4 U145 ( .A(n322), .Y(n320) );
  AND2X2 U146 ( .A(n254), .B(n245), .Y(n53) );
  INVX8 U147 ( .A(n289), .Y(n62) );
  AND3X2 U148 ( .A(n264), .B(n257), .C(n265), .Y(n34) );
  OAI2BB1X2 U149 ( .A0N(B[9]), .A1N(A[9]), .B0(n64), .Y(n317) );
  NOR2X4 U150 ( .A(n143), .B(n56), .Y(n142) );
  NOR2BX2 U151 ( .AN(n61), .B(n62), .Y(n60) );
  NAND2X2 U152 ( .A(B[3]), .B(A[3]), .Y(n98) );
  OAI21X2 U153 ( .A0(A[11]), .A1(B[11]), .B0(n291), .Y(n314) );
  NOR2X2 U154 ( .A(n34), .B(n266), .Y(n262) );
  NAND2X2 U155 ( .A(n245), .B(n244), .Y(n266) );
  AND3X1 U156 ( .A(n168), .B(n169), .C(n170), .Y(n23) );
  NOR2X1 U157 ( .A(n23), .B(n171), .Y(n164) );
  NAND2X1 U158 ( .A(n172), .B(n173), .Y(n171) );
  NAND2X4 U159 ( .A(n25), .B(n26), .Y(SUM[10]) );
  NAND2X4 U160 ( .A(B[23]), .B(n19), .Y(n167) );
  NOR2X4 U161 ( .A(B[15]), .B(A[15]), .Y(n276) );
  NAND2X2 U162 ( .A(B[11]), .B(A[11]), .Y(n309) );
  NAND2X2 U163 ( .A(n112), .B(n129), .Y(n29) );
  NAND2X4 U164 ( .A(n28), .B(n29), .Y(SUM[2]) );
  OAI2BB1X2 U165 ( .A0N(n131), .A1N(n132), .B0(n133), .Y(n115) );
  NAND2X2 U166 ( .A(n53), .B(n296), .Y(n32) );
  NAND2X4 U167 ( .A(n30), .B(n31), .Y(n33) );
  NAND2X4 U168 ( .A(n32), .B(n33), .Y(n45) );
  AND2X4 U169 ( .A(n35), .B(n187), .Y(n213) );
  NAND2BX2 U170 ( .AN(n201), .B(n202), .Y(n199) );
  NAND2X1 U171 ( .A(n79), .B(n17), .Y(n77) );
  OR2X4 U172 ( .A(A[21]), .B(B[21]), .Y(n185) );
  BUFX12 U173 ( .A(n334), .Y(SUM[26]) );
  NOR2BX4 U174 ( .AN(n133), .B(n232), .Y(n231) );
  NOR2X2 U175 ( .A(n276), .B(n58), .Y(n253) );
  NOR2X4 U176 ( .A(n179), .B(n188), .Y(n186) );
  OAI21X2 U177 ( .A0(n188), .A1(n169), .B0(n170), .Y(n191) );
  INVX4 U178 ( .A(n172), .Y(n188) );
  NAND3BX1 U179 ( .AN(n96), .B(n98), .C(n97), .Y(n92) );
  AND2X2 U180 ( .A(n156), .B(n150), .Y(n42) );
  NAND2X2 U181 ( .A(B[25]), .B(A[25]), .Y(n150) );
  INVX4 U182 ( .A(n91), .Y(n74) );
  NAND2X4 U183 ( .A(B[21]), .B(A[21]), .Y(n169) );
  NAND2BX2 U184 ( .AN(n52), .B(n288), .Y(n313) );
  OR2X4 U185 ( .A(A[8]), .B(B[8]), .Y(n290) );
  INVX8 U186 ( .A(n290), .Y(n69) );
  AOI21X4 U187 ( .A0(n305), .A1(n302), .B0(n306), .Y(n304) );
  OR2X4 U188 ( .A(A[12]), .B(B[12]), .Y(n302) );
  INVX2 U189 ( .A(n169), .Y(n200) );
  NAND2X1 U190 ( .A(n185), .B(n169), .Y(n212) );
  NAND3X2 U191 ( .A(n138), .B(n4), .C(n137), .Y(n126) );
  NOR2BX2 U192 ( .AN(n4), .B(n56), .Y(n152) );
  BUFX4 U193 ( .A(n22), .Y(n58) );
  NAND2X2 U194 ( .A(n307), .B(n256), .Y(n306) );
  INVX8 U195 ( .A(n39), .Y(SUM[30]) );
  NAND2X4 U196 ( .A(B[4]), .B(A[4]), .Y(n102) );
  OAI21X2 U197 ( .A0(n112), .A1(n113), .B0(n114), .Y(n108) );
  INVX2 U198 ( .A(n115), .Y(n112) );
  NAND2X4 U199 ( .A(B[5]), .B(A[5]), .Y(n95) );
  AOI21X4 U200 ( .A0(n135), .A1(n124), .B0(n136), .Y(n134) );
  NAND2BX1 U201 ( .AN(n43), .B(n137), .Y(n135) );
  OR2X4 U202 ( .A(A[20]), .B(B[20]), .Y(n184) );
  XOR2X4 U203 ( .A(n132), .B(n231), .Y(SUM[1]) );
  OR2X4 U204 ( .A(A[10]), .B(B[10]), .Y(n291) );
  XOR2X4 U205 ( .A(n108), .B(n109), .Y(SUM[3]) );
  AOI21X2 U206 ( .A0(B[11]), .A1(A[11]), .B0(n292), .Y(n319) );
  NAND4BX4 U207 ( .AN(n331), .B(n332), .C(n131), .D(n130), .Y(n97) );
  NOR2XL U208 ( .A(A[3]), .B(B[3]), .Y(n331) );
  NAND2XL U209 ( .A(n133), .B(n233), .Y(n332) );
  OAI21X4 U210 ( .A0(n235), .A1(n236), .B0(n237), .Y(n234) );
  NAND2X4 U211 ( .A(n75), .B(n67), .Y(n284) );
  OR2X4 U212 ( .A(A[24]), .B(n8), .Y(n157) );
  XNOR2X4 U213 ( .A(n118), .B(n49), .Y(n39) );
  AND2X2 U214 ( .A(n121), .B(n119), .Y(n49) );
  XNOR2X4 U215 ( .A(n41), .B(n134), .Y(SUM[29]) );
  NAND2X4 U216 ( .A(n8), .B(A[24]), .Y(n149) );
  NAND2X2 U217 ( .A(B[20]), .B(A[20]), .Y(n187) );
  AOI21X4 U218 ( .A0(n105), .A1(n91), .B0(n106), .Y(n104) );
  NAND2X2 U219 ( .A(n66), .B(n67), .Y(n65) );
  NOR2BX2 U220 ( .AN(n167), .B(n179), .Y(n190) );
  OAI2BB1X4 U221 ( .A0N(n175), .A1N(n176), .B0(n149), .Y(n174) );
  XOR2X4 U222 ( .A(n103), .B(n104), .Y(SUM[5]) );
  NOR2BX4 U223 ( .AN(n102), .B(n74), .Y(n107) );
  NAND3X4 U224 ( .A(n83), .B(n85), .C(n84), .Y(n67) );
  NAND2XL U225 ( .A(n172), .B(n170), .Y(n44) );
  XNOR2X4 U226 ( .A(n141), .B(n180), .Y(n55) );
  INVX8 U227 ( .A(n55), .Y(SUM[24]) );
  INVXL U228 ( .A(n83), .Y(n82) );
  XOR2X4 U229 ( .A(n99), .B(n40), .Y(SUM[6]) );
  AND2X1 U230 ( .A(n85), .B(n76), .Y(n40) );
  AND2X1 U231 ( .A(n122), .B(n125), .Y(n41) );
  AND2X1 U232 ( .A(n127), .B(n124), .Y(n140) );
  NAND3X4 U233 ( .A(n161), .B(n141), .C(n142), .Y(n137) );
  NOR2X4 U234 ( .A(n218), .B(n219), .Y(n227) );
  XOR2X4 U235 ( .A(n44), .B(n197), .Y(SUM[22]) );
  INVXL U236 ( .A(n121), .Y(n120) );
  OAI21X4 U237 ( .A0(n277), .A1(n278), .B0(n279), .Y(n273) );
  AND3X4 U238 ( .A(n211), .B(n210), .C(n209), .Y(n203) );
  INVXL U239 ( .A(n254), .Y(n252) );
  CLKINVX3 U240 ( .A(n233), .Y(n132) );
  OR2X4 U241 ( .A(A[2]), .B(B[2]), .Y(n130) );
  OR2X4 U242 ( .A(B[5]), .B(A[5]), .Y(n90) );
  OR2X4 U243 ( .A(A[4]), .B(B[4]), .Y(n91) );
  OR2X4 U244 ( .A(A[22]), .B(B[22]), .Y(n172) );
  OR2X4 U245 ( .A(A[25]), .B(B[25]), .Y(n156) );
  OR2X4 U246 ( .A(A[26]), .B(B[26]), .Y(n148) );
  NOR2XL U247 ( .A(A[9]), .B(B[9]), .Y(n46) );
  NAND2X2 U248 ( .A(B[10]), .B(A[10]), .Y(n310) );
  NOR2BX1 U249 ( .AN(n233), .B(n47), .Y(n337) );
  NOR2XL U250 ( .A(A[0]), .B(B[0]), .Y(n47) );
  NOR2XL U251 ( .A(n179), .B(n145), .Y(n175) );
  NAND2X1 U252 ( .A(n148), .B(n155), .Y(n159) );
  NOR2BX1 U253 ( .AN(n187), .B(n195), .Y(n220) );
  NOR2BX1 U254 ( .AN(n64), .B(n69), .Y(n78) );
  INVX1 U255 ( .A(n102), .Y(n106) );
  NAND4BXL U256 ( .AN(n73), .B(n91), .C(n76), .D(n75), .Y(n286) );
  XOR2X4 U257 ( .A(n48), .B(n312), .Y(SUM[12]) );
  INVX1 U258 ( .A(n127), .Y(n136) );
  INVX1 U259 ( .A(n131), .Y(n232) );
  NAND2XL U260 ( .A(n287), .B(n257), .Y(n303) );
  OR2X2 U261 ( .A(n127), .B(n128), .Y(n50) );
  INVX1 U262 ( .A(n130), .Y(n113) );
  NAND2X1 U263 ( .A(n95), .B(n102), .Y(n326) );
  XNOR2X4 U264 ( .A(n294), .B(n295), .Y(n51) );
  INVX8 U265 ( .A(n51), .Y(SUM[15]) );
  INVXL U266 ( .A(n229), .Y(n261) );
  AND2X1 U267 ( .A(n311), .B(n310), .Y(n52) );
  OAI21X2 U268 ( .A0(n203), .A1(n204), .B0(n205), .Y(n201) );
  XNOR2X4 U269 ( .A(n258), .B(n259), .Y(n54) );
  INVX8 U270 ( .A(n54), .Y(SUM[17]) );
  NOR2X4 U271 ( .A(A[27]), .B(B[27]), .Y(n56) );
  NAND4BX4 U272 ( .AN(n182), .B(n183), .C(n57), .D(n184), .Y(n165) );
  NAND2X2 U273 ( .A(B[19]), .B(A[19]), .Y(n206) );
  NAND3X2 U274 ( .A(n168), .B(n169), .C(n170), .Y(n178) );
  NAND2X1 U275 ( .A(B[28]), .B(A[28]), .Y(n127) );
  OR2X2 U276 ( .A(A[28]), .B(B[28]), .Y(n124) );
  OR2X2 U277 ( .A(A[29]), .B(B[29]), .Y(n125) );
  NAND3X2 U278 ( .A(n209), .B(n210), .C(n228), .Y(n217) );
  NAND2XL U279 ( .A(B[18]), .B(A[18]), .Y(n228) );
  NAND2XL U280 ( .A(B[18]), .B(A[18]), .Y(n211) );
  OR2X2 U281 ( .A(A[30]), .B(B[30]), .Y(n119) );
  NAND2X1 U282 ( .A(B[29]), .B(A[29]), .Y(n122) );
  NAND2X1 U283 ( .A(B[30]), .B(A[30]), .Y(n121) );
  NAND2X1 U284 ( .A(B[0]), .B(A[0]), .Y(n233) );
  XNOR2X1 U285 ( .A(B[31]), .B(A[31]), .Y(n116) );
  NAND3BX4 U286 ( .AN(n96), .B(n98), .C(n97), .Y(n71) );
  NAND2X1 U287 ( .A(n75), .B(n76), .Y(n70) );
  OAI21X2 U288 ( .A0(n296), .A1(n58), .B0(n254), .Y(n294) );
  NOR2X1 U289 ( .A(n19), .B(B[23]), .Y(n182) );
  NAND3X1 U290 ( .A(n289), .B(n290), .C(n291), .Y(n277) );
  INVX4 U291 ( .A(n242), .Y(n271) );
  INVX8 U292 ( .A(n207), .Y(n219) );
  INVX8 U293 ( .A(n208), .Y(n218) );
  NOR2X2 U294 ( .A(n218), .B(n219), .Y(n216) );
  NAND2X1 U295 ( .A(n230), .B(n207), .Y(n236) );
  NAND2XL U296 ( .A(B[14]), .B(A[14]), .Y(n265) );
  NAND2XL U297 ( .A(n245), .B(n244), .Y(n268) );
  NAND2X1 U298 ( .A(B[7]), .B(A[7]), .Y(n83) );
  AOI21X1 U299 ( .A0(B[7]), .A1(A[7]), .B0(n68), .Y(n87) );
  INVX8 U300 ( .A(n288), .Y(n292) );
  NOR2X2 U301 ( .A(n225), .B(n226), .Y(n247) );
  INVX8 U302 ( .A(n75), .Y(n68) );
  NOR2X2 U303 ( .A(n81), .B(n82), .Y(n79) );
  NAND2X1 U304 ( .A(n95), .B(n94), .Y(n100) );
  NAND2XL U305 ( .A(n90), .B(n76), .Y(n89) );
  NAND3X2 U306 ( .A(n90), .B(n91), .C(n71), .Y(n101) );
  AOI21X1 U307 ( .A0(n84), .A1(n85), .B0(n68), .Y(n81) );
  NAND3XL U308 ( .A(n98), .B(n285), .C(n97), .Y(n282) );
  NAND2X2 U309 ( .A(B[6]), .B(A[6]), .Y(n85) );
  NAND2X4 U310 ( .A(n284), .B(n80), .Y(n315) );
  XOR2X4 U311 ( .A(n59), .B(n60), .Y(SUM[9]) );
  NAND3X4 U312 ( .A(n63), .B(n64), .C(n65), .Y(n59) );
  XOR2X4 U313 ( .A(n77), .B(n78), .Y(SUM[8]) );
  OAI21X4 U314 ( .A0(n88), .A1(n89), .B0(n85), .Y(n86) );
  NAND2BX4 U315 ( .AN(n100), .B(n101), .Y(n99) );
  XOR2X4 U316 ( .A(n126), .B(n140), .Y(SUM[28]) );
  OAI21X4 U317 ( .A0(n153), .A1(n154), .B0(n155), .Y(n151) );
  AOI21X4 U318 ( .A0(n157), .A1(n141), .B0(n158), .Y(n153) );
  XOR2X4 U319 ( .A(n159), .B(n160), .Y(n334) );
  AOI21X4 U320 ( .A0(n161), .A1(n162), .B0(n163), .Y(n160) );
  AND2X2 U321 ( .A(n149), .B(n167), .Y(n166) );
  XOR2X4 U322 ( .A(n174), .B(n42), .Y(SUM[25]) );
  NOR2BX4 U323 ( .AN(n149), .B(n145), .Y(n180) );
  NAND2BX4 U324 ( .AN(n181), .B(n165), .Y(n141) );
  OAI2BB1X4 U325 ( .A0N(n186), .A1N(n178), .B0(n167), .Y(n181) );
  XOR2X4 U326 ( .A(n189), .B(n190), .Y(SUM[23]) );
  OR2X4 U327 ( .A(A[23]), .B(B[23]), .Y(n173) );
  NAND2BX4 U328 ( .AN(n191), .B(n192), .Y(n189) );
  AOI21X4 U329 ( .A0(n198), .A1(n199), .B0(n200), .Y(n197) );
  AND2X2 U330 ( .A(n187), .B(n206), .Y(n205) );
  XOR2X4 U331 ( .A(n213), .B(n212), .Y(n335) );
  OAI2BB1X4 U332 ( .A0N(n216), .A1N(n217), .B0(n206), .Y(n215) );
  XOR2X4 U333 ( .A(n16), .B(n220), .Y(SUM[20]) );
  NAND2BX4 U334 ( .AN(n221), .B(n202), .Y(n183) );
  NAND3X4 U335 ( .A(n222), .B(n223), .C(n224), .Y(n202) );
  NOR2X4 U336 ( .A(n218), .B(n219), .Y(n223) );
  XOR2X4 U337 ( .A(n234), .B(n14), .Y(SUM[19]) );
  OR2X4 U338 ( .A(A[19]), .B(B[19]), .Y(n208) );
  XOR2X4 U339 ( .A(n246), .B(n13), .Y(SUM[18]) );
  OR2X4 U340 ( .A(A[18]), .B(B[18]), .Y(n207) );
  AOI21X4 U341 ( .A0(n238), .A1(n260), .B0(n261), .Y(n259) );
  OR2X4 U342 ( .A(A[16]), .B(B[16]), .Y(n238) );
  NAND2X4 U343 ( .A(B[16]), .B(A[16]), .Y(n229) );
  OAI21X4 U344 ( .A0(n243), .A1(n268), .B0(n269), .Y(n224) );
  NOR2X4 U345 ( .A(n270), .B(n271), .Y(n269) );
  NAND3BX4 U346 ( .AN(n272), .B(n273), .C(n274), .Y(n242) );
  NOR2X4 U347 ( .A(n275), .B(n276), .Y(n274) );
  AND3X4 U348 ( .A(n257), .B(n293), .C(n264), .Y(n243) );
  OR2X4 U349 ( .A(B[15]), .B(A[15]), .Y(n244) );
  NOR3X4 U350 ( .A(n298), .B(n297), .C(n299), .Y(n296) );
  NOR2X4 U351 ( .A(n300), .B(n301), .Y(n297) );
  OR2X4 U352 ( .A(A[14]), .B(B[14]), .Y(n245) );
  XOR2X4 U353 ( .A(n303), .B(n304), .Y(SUM[13]) );
  OR2X4 U354 ( .A(B[13]), .B(A[13]), .Y(n287) );
  NAND3BX4 U355 ( .AN(n314), .B(n315), .C(n316), .Y(n300) );
  NAND3X4 U356 ( .A(n291), .B(n289), .C(n317), .Y(n311) );
  XOR2X4 U357 ( .A(n318), .B(n319), .Y(SUM[11]) );
  OR2X4 U358 ( .A(A[11]), .B(B[11]), .Y(n288) );
  NAND2X4 U359 ( .A(n324), .B(n325), .Y(n322) );
  NAND3X4 U360 ( .A(n90), .B(n76), .C(n326), .Y(n84) );
  OR2X4 U361 ( .A(A[9]), .B(B[9]), .Y(n289) );
  OR2X4 U362 ( .A(A[7]), .B(B[7]), .Y(n75) );
  OR2X4 U363 ( .A(A[6]), .B(B[6]), .Y(n76) );
  NAND2BX4 U364 ( .AN(n114), .B(n111), .Y(n285) );
endmodule


module hash_core_DW01_add_26 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n267, n268, n269, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266;

  AOI21X4 U2 ( .A0(n130), .A1(n129), .B0(n131), .Y(n127) );
  NAND2X1 U3 ( .A(B[30]), .B(A[30]), .Y(n78) );
  AOI21X1 U4 ( .A0(n84), .A1(n85), .B0(n86), .Y(n79) );
  AOI2BB1X2 U5 ( .A0N(n87), .A1N(n88), .B0(n89), .Y(n84) );
  INVX2 U6 ( .A(n48), .Y(n241) );
  INVX4 U7 ( .A(n11), .Y(SUM[24]) );
  AOI21X4 U8 ( .A0(n193), .A1(n188), .B0(n194), .Y(n176) );
  NOR2BX2 U9 ( .AN(n58), .B(n57), .Y(n60) );
  NAND2X2 U10 ( .A(B[6]), .B(A[6]), .Y(n58) );
  NOR2BXL U11 ( .AN(n217), .B(n43), .Y(n235) );
  BUFX8 U12 ( .A(n269), .Y(SUM[18]) );
  INVX4 U13 ( .A(n106), .Y(n198) );
  CLKINVX4 U14 ( .A(n8), .Y(n2) );
  INVX8 U15 ( .A(n2), .Y(n3) );
  NAND2XL U16 ( .A(B[9]), .B(A[9]), .Y(n8) );
  NOR2X4 U17 ( .A(n185), .B(n186), .Y(n179) );
  BUFX8 U18 ( .A(n268), .Y(SUM[21]) );
  NAND2X1 U19 ( .A(B[24]), .B(A[24]), .Y(n148) );
  XOR2X2 U20 ( .A(n107), .B(n197), .Y(SUM[1]) );
  CLKINVX4 U21 ( .A(n74), .Y(n265) );
  OAI21X2 U22 ( .A0(n72), .A1(n73), .B0(n74), .Y(n68) );
  NOR2BX2 U23 ( .AN(n74), .B(n73), .Y(n104) );
  NAND2X2 U24 ( .A(B[2]), .B(A[2]), .Y(n74) );
  INVX4 U25 ( .A(n191), .Y(n208) );
  NAND2X2 U26 ( .A(n191), .B(n192), .Y(n187) );
  OR2X4 U27 ( .A(A[16]), .B(B[16]), .Y(n191) );
  OAI21X2 U28 ( .A0(n79), .A1(n80), .B0(n81), .Y(n77) );
  NAND2X1 U29 ( .A(B[1]), .B(A[1]), .Y(n108) );
  OAI21X4 U30 ( .A0(n222), .A1(n218), .B0(n223), .Y(n221) );
  NAND2X2 U31 ( .A(n105), .B(n262), .Y(n264) );
  OR2X4 U32 ( .A(A[3]), .B(B[3]), .Y(n262) );
  NAND2X4 U33 ( .A(B[12]), .B(A[12]), .Y(n215) );
  BUFX8 U34 ( .A(n136), .Y(n5) );
  NAND2XL U35 ( .A(B[23]), .B(A[23]), .Y(n136) );
  NOR2X4 U36 ( .A(A[4]), .B(B[4]), .Y(n38) );
  NOR2X2 U37 ( .A(n265), .B(n266), .Y(n263) );
  OAI21X1 U38 ( .A0(n198), .A1(n199), .B0(n108), .Y(n266) );
  BUFX8 U39 ( .A(n148), .Y(n6) );
  INVX1 U40 ( .A(n214), .Y(n213) );
  NAND3X2 U41 ( .A(A[24]), .B(B[24]), .C(n118), .Y(n133) );
  CLKINVX2 U42 ( .A(n37), .Y(n31) );
  NOR2X2 U43 ( .A(n183), .B(n195), .Y(n194) );
  CLKINVX3 U44 ( .A(n182), .Y(n181) );
  INVX1 U45 ( .A(A[20]), .Y(n14) );
  NAND2X1 U46 ( .A(B[20]), .B(A[20]), .Y(n171) );
  INVX1 U47 ( .A(n173), .Y(n175) );
  OR2X2 U48 ( .A(A[1]), .B(B[1]), .Y(n106) );
  INVX4 U49 ( .A(n188), .Y(n184) );
  NOR2X1 U50 ( .A(n82), .B(n41), .Y(n81) );
  INVX1 U51 ( .A(n102), .Y(n101) );
  NAND2X1 U52 ( .A(B[18]), .B(A[18]), .Y(n195) );
  INVX1 U53 ( .A(n100), .Y(n86) );
  BUFX3 U54 ( .A(n149), .Y(n17) );
  NAND2X1 U55 ( .A(B[26]), .B(A[26]), .Y(n128) );
  INVX1 U56 ( .A(n28), .Y(n66) );
  INVX1 U57 ( .A(n199), .Y(n107) );
  NOR2BX1 U58 ( .AN(n50), .B(n51), .Y(n49) );
  INVX1 U59 ( .A(n251), .Y(n51) );
  CLKINVX3 U60 ( .A(n9), .Y(SUM[6]) );
  NAND2X2 U61 ( .A(n22), .B(n23), .Y(SUM[9]) );
  INVX1 U62 ( .A(n46), .Y(n21) );
  CLKBUFX8 U63 ( .A(n267), .Y(SUM[22]) );
  NOR2BX1 U64 ( .AN(n161), .B(n165), .Y(n167) );
  INVX2 U65 ( .A(n234), .Y(n233) );
  NOR2BX1 U66 ( .AN(n196), .B(n185), .Y(n205) );
  NAND2X2 U67 ( .A(n24), .B(n53), .Y(n27) );
  XOR2X2 U68 ( .A(n63), .B(n64), .Y(SUM[5]) );
  OAI21X4 U69 ( .A0(n263), .A1(n264), .B0(n70), .Y(n224) );
  BUFX3 U70 ( .A(n83), .Y(n7) );
  OR2X2 U71 ( .A(A[26]), .B(B[26]), .Y(n90) );
  NOR2X2 U72 ( .A(A[26]), .B(B[26]), .Y(n116) );
  INVX1 U73 ( .A(n229), .Y(n238) );
  OR2X2 U74 ( .A(A[12]), .B(B[12]), .Y(n229) );
  NAND2X1 U75 ( .A(B[29]), .B(A[29]), .Y(n83) );
  XNOR2X1 U76 ( .A(n59), .B(n60), .Y(n9) );
  AND2X2 U77 ( .A(B[26]), .B(A[26]), .Y(n10) );
  XNOR2X1 U78 ( .A(n155), .B(n120), .Y(n11) );
  AND2X4 U79 ( .A(n206), .B(n186), .Y(n12) );
  NAND2X1 U80 ( .A(n45), .B(n21), .Y(n22) );
  INVX3 U81 ( .A(n120), .Y(n154) );
  NOR2BX1 U82 ( .AN(n215), .B(n238), .Y(n240) );
  OAI21X1 U83 ( .A0(n241), .A1(n218), .B0(n223), .Y(n13) );
  NOR2BX4 U84 ( .AN(n248), .B(n249), .Y(n242) );
  AOI21X4 U85 ( .A0(n245), .A1(n254), .B0(n255), .Y(n253) );
  NOR2X2 U86 ( .A(B[27]), .B(A[27]), .Y(n117) );
  NOR2X1 U87 ( .A(B[27]), .B(A[27]), .Y(n126) );
  NAND3BX4 U88 ( .AN(n14), .B(B[20]), .C(n159), .Y(n158) );
  NAND3X4 U89 ( .A(n245), .B(n246), .C(n247), .Y(n243) );
  NAND4X4 U90 ( .A(n251), .B(n246), .C(n245), .D(n244), .Y(n218) );
  NAND2X2 U91 ( .A(B[8]), .B(A[8]), .Y(n50) );
  INVXL U92 ( .A(n172), .Y(n15) );
  INVX2 U93 ( .A(n15), .Y(n16) );
  NOR2BX4 U94 ( .AN(n5), .B(n141), .Y(n163) );
  INVX1 U95 ( .A(n156), .Y(n141) );
  INVXL U96 ( .A(n42), .Y(n35) );
  NOR2BXL U97 ( .AN(n216), .B(n42), .Y(n237) );
  AOI21X4 U98 ( .A0(B[21]), .A1(A[21]), .B0(n160), .Y(n157) );
  INVX4 U99 ( .A(n161), .Y(n160) );
  NOR2BX1 U100 ( .AN(n62), .B(n37), .Y(n64) );
  NAND2X2 U101 ( .A(B[5]), .B(A[5]), .Y(n62) );
  AOI21X1 U102 ( .A0(n219), .A1(n224), .B0(n225), .Y(n222) );
  INVX2 U103 ( .A(n226), .Y(n225) );
  NAND2X1 U104 ( .A(B[28]), .B(A[28]), .Y(n113) );
  NAND2X2 U105 ( .A(B[13]), .B(A[13]), .Y(n216) );
  OR2X2 U106 ( .A(B[27]), .B(A[27]), .Y(n39) );
  NAND2X1 U107 ( .A(n97), .B(n7), .Y(n109) );
  OAI2BB1X4 U108 ( .A0N(n236), .A1N(n35), .B0(n216), .Y(n234) );
  NOR2X4 U109 ( .A(n33), .B(n43), .Y(n211) );
  NOR2X4 U110 ( .A(B[15]), .B(A[15]), .Y(n33) );
  NOR2BXL U111 ( .AN(n214), .B(n33), .Y(n232) );
  NOR2X4 U112 ( .A(A[14]), .B(B[14]), .Y(n43) );
  AOI21X2 U113 ( .A0(n98), .A1(n85), .B0(n99), .Y(n94) );
  NOR2X2 U114 ( .A(n89), .B(n101), .Y(n98) );
  NAND2X2 U115 ( .A(n190), .B(n191), .Y(n206) );
  XOR2X2 U116 ( .A(n168), .B(n170), .Y(n268) );
  NAND4BX2 U117 ( .AN(n187), .B(n190), .C(n189), .D(n188), .Y(n177) );
  INVX2 U118 ( .A(n97), .Y(n82) );
  OAI21X2 U119 ( .A0(n82), .A1(n96), .B0(n7), .Y(n95) );
  NOR2BX2 U120 ( .AN(n6), .B(n146), .Y(n155) );
  NAND2XL U121 ( .A(B[19]), .B(A[19]), .Y(n182) );
  XOR2X4 U122 ( .A(n234), .B(n235), .Y(SUM[14]) );
  CLKINVX4 U123 ( .A(n250), .Y(n249) );
  NAND3BX4 U124 ( .AN(n149), .B(n5), .C(n151), .Y(n120) );
  NAND2X2 U125 ( .A(B[21]), .B(A[21]), .Y(n169) );
  AND2X4 U126 ( .A(n77), .B(n78), .Y(n32) );
  NAND2X4 U127 ( .A(B[15]), .B(A[15]), .Y(n214) );
  AND2X4 U128 ( .A(B[4]), .B(A[4]), .Y(n28) );
  AND2X4 U129 ( .A(n211), .B(n212), .Y(n18) );
  NOR2X4 U130 ( .A(n18), .B(n213), .Y(n210) );
  NAND2X4 U131 ( .A(B[14]), .B(A[14]), .Y(n217) );
  OAI21X4 U132 ( .A0(n56), .A1(n57), .B0(n58), .Y(n52) );
  INVX4 U133 ( .A(n138), .Y(n165) );
  NAND3BX2 U134 ( .AN(n37), .B(n260), .C(n61), .Y(n259) );
  NAND4BBX4 U135 ( .AN(n37), .BN(n38), .C(n61), .D(n261), .Y(n227) );
  NOR2X4 U136 ( .A(A[5]), .B(B[5]), .Y(n37) );
  NOR2BX4 U137 ( .AN(n54), .B(n55), .Y(n53) );
  NAND2X2 U138 ( .A(B[7]), .B(A[7]), .Y(n54) );
  XOR2X4 U139 ( .A(B[31]), .B(A[31]), .Y(n76) );
  XOR2X2 U140 ( .A(n236), .B(n237), .Y(SUM[13]) );
  XOR2X1 U141 ( .A(n48), .B(n49), .Y(SUM[8]) );
  INVXL U142 ( .A(n195), .Y(n203) );
  NOR2BXL U143 ( .AN(n195), .B(n184), .Y(n204) );
  NAND2X2 U144 ( .A(B[17]), .B(A[17]), .Y(n196) );
  NOR2X2 U145 ( .A(A[30]), .B(B[30]), .Y(n41) );
  NOR2X4 U146 ( .A(B[13]), .B(A[13]), .Y(n42) );
  NAND3BX2 U147 ( .AN(n134), .B(n135), .C(n5), .Y(n130) );
  OR2X4 U148 ( .A(A[2]), .B(B[2]), .Y(n105) );
  NAND2X2 U149 ( .A(n257), .B(n46), .Y(n23) );
  NAND2X2 U150 ( .A(n52), .B(n25), .Y(n26) );
  NAND2X4 U151 ( .A(n26), .B(n27), .Y(SUM[7]) );
  CLKINVX4 U152 ( .A(n52), .Y(n24) );
  INVXL U153 ( .A(n53), .Y(n25) );
  XOR2X4 U154 ( .A(n253), .B(n252), .Y(SUM[11]) );
  OR2X4 U155 ( .A(n65), .B(n227), .Y(n29) );
  NAND2X4 U156 ( .A(n29), .B(n226), .Y(n48) );
  AND2X2 U157 ( .A(n48), .B(n251), .Y(n36) );
  NOR2X2 U158 ( .A(n38), .B(n65), .Y(n30) );
  OR2X4 U159 ( .A(n30), .B(n28), .Y(n63) );
  INVX4 U160 ( .A(n224), .Y(n65) );
  OAI2BB1X4 U161 ( .A0N(n63), .A1N(n31), .B0(n62), .Y(n59) );
  NAND2X2 U162 ( .A(n62), .B(n66), .Y(n260) );
  INVX1 U163 ( .A(n91), .Y(n87) );
  OAI2BB1X4 U164 ( .A0N(n121), .A1N(n118), .B0(n122), .Y(n91) );
  NAND2BXL U165 ( .AN(n41), .B(n78), .Y(n92) );
  INVX4 U166 ( .A(n45), .Y(n257) );
  NOR3BX4 U167 ( .AN(n156), .B(n140), .C(n139), .Y(n149) );
  NAND3X4 U168 ( .A(n102), .B(n103), .C(n85), .Y(n111) );
  CLKINVX2 U169 ( .A(n123), .Y(n132) );
  XOR2X2 U170 ( .A(n166), .B(n167), .Y(n267) );
  OAI2BB1X1 U171 ( .A0N(n106), .A1N(n107), .B0(n108), .Y(n75) );
  OAI2BB1X4 U172 ( .A0N(n229), .A1N(n239), .B0(n215), .Y(n236) );
  INVXL U173 ( .A(n248), .Y(n255) );
  AND2X1 U174 ( .A(n248), .B(n245), .Y(n256) );
  OAI21X4 U175 ( .A0(n257), .A1(n47), .B0(n3), .Y(n254) );
  NOR2BXL U176 ( .AN(n108), .B(n198), .Y(n197) );
  NAND2XL U177 ( .A(n97), .B(n100), .Y(n99) );
  OAI2BB1X4 U178 ( .A0N(n159), .A1N(n168), .B0(n169), .Y(n166) );
  AND2X1 U179 ( .A(n123), .B(n118), .Y(n153) );
  NAND2X4 U180 ( .A(n159), .B(n138), .Y(n139) );
  INVXL U181 ( .A(n262), .Y(n71) );
  AND2X1 U182 ( .A(n169), .B(n159), .Y(n170) );
  NAND2XL U183 ( .A(B[3]), .B(A[3]), .Y(n70) );
  NAND2XL U184 ( .A(B[0]), .B(A[0]), .Y(n199) );
  XNOR2X4 U185 ( .A(n32), .B(n76), .Y(SUM[31]) );
  AND3X4 U186 ( .A(n120), .B(n119), .C(n118), .Y(n40) );
  NOR2BX1 U187 ( .AN(n199), .B(n34), .Y(SUM[0]) );
  NOR2XL U188 ( .A(A[0]), .B(B[0]), .Y(n34) );
  INVXL U189 ( .A(n227), .Y(n219) );
  NOR2XL U190 ( .A(n139), .B(n140), .Y(n134) );
  XOR2X1 U191 ( .A(n190), .B(n207), .Y(SUM[16]) );
  NOR2BX1 U192 ( .AN(n186), .B(n208), .Y(n207) );
  XOR2X2 U193 ( .A(n202), .B(n204), .Y(n269) );
  INVX1 U194 ( .A(n59), .Y(n56) );
  NOR2BX1 U195 ( .AN(n3), .B(n47), .Y(n46) );
  NAND2XL U196 ( .A(n182), .B(n189), .Y(n200) );
  NAND2XL U197 ( .A(n244), .B(n250), .Y(n252) );
  XOR2X1 U198 ( .A(n224), .B(n67), .Y(SUM[4]) );
  NOR2BX1 U199 ( .AN(n66), .B(n38), .Y(n67) );
  INVX1 U200 ( .A(n113), .Y(n112) );
  NAND2X1 U201 ( .A(n128), .B(n90), .Y(n143) );
  INVXL U202 ( .A(n61), .Y(n57) );
  INVX1 U203 ( .A(n103), .Y(n89) );
  NAND2BX4 U204 ( .AN(n36), .B(n50), .Y(n45) );
  NAND2XL U205 ( .A(n137), .B(n138), .Y(n135) );
  XOR2X1 U206 ( .A(n68), .B(n69), .Y(SUM[3]) );
  NOR2BX1 U207 ( .AN(n70), .B(n71), .Y(n69) );
  INVX1 U208 ( .A(n75), .Y(n72) );
  XOR2X1 U209 ( .A(n75), .B(n104), .Y(SUM[2]) );
  INVX1 U210 ( .A(n105), .Y(n73) );
  NAND2X2 U211 ( .A(B[16]), .B(A[16]), .Y(n186) );
  NAND3X4 U212 ( .A(n39), .B(n90), .C(n91), .Y(n102) );
  NAND2X2 U213 ( .A(B[10]), .B(A[10]), .Y(n248) );
  NAND2X4 U214 ( .A(n40), .B(n115), .Y(n85) );
  NAND2XL U215 ( .A(A[28]), .B(B[28]), .Y(n96) );
  OAI2BB1X1 U216 ( .A0N(B[28]), .A1N(A[28]), .B0(n7), .Y(n80) );
  NAND2X4 U217 ( .A(n209), .B(n210), .Y(n190) );
  XOR2X1 U218 ( .A(n16), .B(n174), .Y(SUM[20]) );
  OAI21X4 U219 ( .A0(n147), .A1(n146), .B0(n6), .Y(n145) );
  NAND2X2 U220 ( .A(B[25]), .B(A[25]), .Y(n123) );
  NOR2X4 U221 ( .A(n17), .B(n150), .Y(n147) );
  NAND2X2 U222 ( .A(n119), .B(n118), .Y(n142) );
  NAND2X2 U223 ( .A(B[11]), .B(A[11]), .Y(n250) );
  OAI21XL U224 ( .A0(B[27]), .A1(A[27]), .B0(n90), .Y(n88) );
  XNOR2X4 U225 ( .A(n12), .B(n205), .Y(SUM[17]) );
  INVX4 U226 ( .A(n166), .Y(n164) );
  INVX8 U227 ( .A(n192), .Y(n185) );
  AND2X1 U228 ( .A(A[24]), .B(B[24]), .Y(n121) );
  XOR2X1 U229 ( .A(n13), .B(n240), .Y(SUM[12]) );
  INVX8 U230 ( .A(n189), .Y(n183) );
  XOR2X4 U231 ( .A(n92), .B(n93), .Y(SUM[30]) );
  NOR2X4 U232 ( .A(n94), .B(n95), .Y(n93) );
  XOR2X4 U233 ( .A(n109), .B(n110), .Y(SUM[29]) );
  AOI21X4 U234 ( .A0(n111), .A1(n100), .B0(n112), .Y(n110) );
  OR2X4 U235 ( .A(A[29]), .B(B[29]), .Y(n97) );
  XOR2X4 U236 ( .A(n111), .B(n114), .Y(SUM[28]) );
  NOR2BX4 U237 ( .AN(n113), .B(n86), .Y(n114) );
  OR2X4 U238 ( .A(A[28]), .B(B[28]), .Y(n100) );
  NOR2X4 U239 ( .A(n116), .B(n117), .Y(n115) );
  NOR2BX4 U240 ( .AN(n123), .B(n10), .Y(n122) );
  XOR2X4 U241 ( .A(n124), .B(n125), .Y(SUM[27]) );
  NOR2BX4 U242 ( .AN(n103), .B(n126), .Y(n125) );
  NAND2X4 U243 ( .A(B[27]), .B(A[27]), .Y(n103) );
  OAI21X4 U244 ( .A0(n127), .A1(n116), .B0(n128), .Y(n124) );
  NAND2BX4 U245 ( .AN(n132), .B(n133), .Y(n131) );
  NOR2X4 U246 ( .A(n141), .B(n142), .Y(n129) );
  XOR2X4 U247 ( .A(n143), .B(n144), .Y(SUM[26]) );
  AOI21X4 U248 ( .A0(n118), .A1(n145), .B0(n132), .Y(n144) );
  NAND2X4 U249 ( .A(n151), .B(n5), .Y(n150) );
  XOR2X4 U250 ( .A(n152), .B(n153), .Y(SUM[25]) );
  OR2X4 U251 ( .A(A[25]), .B(B[25]), .Y(n118) );
  OAI21X4 U252 ( .A0(n146), .A1(n154), .B0(n6), .Y(n152) );
  CLKINVX3 U253 ( .A(n119), .Y(n146) );
  OR2X4 U254 ( .A(A[24]), .B(B[24]), .Y(n119) );
  NAND3X4 U255 ( .A(n138), .B(n156), .C(n137), .Y(n151) );
  NAND2X4 U256 ( .A(n157), .B(n158), .Y(n137) );
  XOR2X4 U257 ( .A(n162), .B(n163), .Y(SUM[23]) );
  OR2X4 U258 ( .A(A[23]), .B(B[23]), .Y(n156) );
  OAI21X4 U259 ( .A0(n164), .A1(n165), .B0(n161), .Y(n162) );
  OR2X4 U260 ( .A(B[22]), .B(A[22]), .Y(n138) );
  NAND2X4 U261 ( .A(B[22]), .B(A[22]), .Y(n161) );
  OR2X4 U262 ( .A(A[21]), .B(B[21]), .Y(n159) );
  NAND2X4 U263 ( .A(n140), .B(n171), .Y(n168) );
  NAND2X4 U264 ( .A(n173), .B(n172), .Y(n140) );
  NOR2BX4 U265 ( .AN(n171), .B(n175), .Y(n174) );
  OR2X4 U266 ( .A(A[20]), .B(B[20]), .Y(n173) );
  NAND3X4 U267 ( .A(n176), .B(n177), .C(n178), .Y(n172) );
  AOI21X4 U268 ( .A0(n179), .A1(n180), .B0(n181), .Y(n178) );
  NOR2X4 U269 ( .A(n183), .B(n184), .Y(n180) );
  NOR2X4 U270 ( .A(n183), .B(n196), .Y(n193) );
  XOR2X4 U271 ( .A(n201), .B(n200), .Y(SUM[19]) );
  AOI21X4 U272 ( .A0(n202), .A1(n188), .B0(n203), .Y(n201) );
  OR2X4 U273 ( .A(B[19]), .B(A[19]), .Y(n189) );
  OR2X4 U274 ( .A(A[18]), .B(B[18]), .Y(n188) );
  OAI21X4 U275 ( .A0(n12), .A1(n185), .B0(n196), .Y(n202) );
  OR2X4 U276 ( .A(A[17]), .B(B[17]), .Y(n192) );
  OAI211X2 U277 ( .A0(n42), .A1(n215), .B0(n216), .C0(n217), .Y(n212) );
  NAND2BX4 U278 ( .AN(n220), .B(n221), .Y(n209) );
  NAND3BX4 U279 ( .AN(n228), .B(n229), .C(n230), .Y(n220) );
  NOR2X4 U280 ( .A(n43), .B(n42), .Y(n230) );
  NOR2X4 U281 ( .A(A[15]), .B(B[15]), .Y(n228) );
  XOR2X4 U282 ( .A(n231), .B(n232), .Y(SUM[15]) );
  OAI21X4 U283 ( .A0(n233), .A1(n43), .B0(n217), .Y(n231) );
  OAI21X4 U284 ( .A0(n241), .A1(n218), .B0(n223), .Y(n239) );
  OAI2BB1X4 U285 ( .A0N(n242), .A1N(n243), .B0(n244), .Y(n223) );
  NAND2X4 U286 ( .A(n3), .B(n50), .Y(n247) );
  OR2X4 U287 ( .A(B[11]), .B(A[11]), .Y(n244) );
  XOR2X4 U288 ( .A(n254), .B(n256), .Y(SUM[10]) );
  OR2X4 U289 ( .A(A[10]), .B(B[10]), .Y(n245) );
  CLKINVX3 U290 ( .A(n246), .Y(n47) );
  OR2X4 U291 ( .A(A[9]), .B(B[9]), .Y(n246) );
  OR2X4 U292 ( .A(A[8]), .B(B[8]), .Y(n251) );
  NAND2BX4 U293 ( .AN(n55), .B(n258), .Y(n226) );
  NAND3X4 U294 ( .A(n259), .B(n58), .C(n54), .Y(n258) );
  CLKINVX3 U295 ( .A(n261), .Y(n55) );
  OR2X4 U296 ( .A(B[7]), .B(A[7]), .Y(n261) );
  OR2X4 U297 ( .A(A[6]), .B(B[6]), .Y(n61) );
endmodule


module hash_core_DW01_add_27 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n271, n272, n273, n274, n275, n2, n4, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n21, n22, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270;

  OAI21X4 U2 ( .A0(n224), .A1(n220), .B0(n225), .Y(n223) );
  OAI21X4 U3 ( .A0(n25), .A1(n265), .B0(n63), .Y(n61) );
  OR2X2 U4 ( .A(B[27]), .B(A[27]), .Y(n37) );
  NAND3BX2 U5 ( .AN(n10), .B(B[20]), .C(n159), .Y(n158) );
  OR2X4 U6 ( .A(A[21]), .B(B[21]), .Y(n159) );
  NAND2X4 U7 ( .A(n150), .B(n135), .Y(n149) );
  OR2X4 U8 ( .A(A[16]), .B(B[16]), .Y(n191) );
  BUFX3 U9 ( .A(n273), .Y(SUM[8]) );
  NOR2BXL U10 ( .AN(n215), .B(n38), .Y(n233) );
  OR2X4 U11 ( .A(A[15]), .B(B[15]), .Y(n41) );
  OAI21X4 U12 ( .A0(n145), .A1(n146), .B0(n147), .Y(n144) );
  NOR2X2 U13 ( .A(A[15]), .B(B[15]), .Y(n38) );
  NOR2X1 U14 ( .A(n269), .B(n270), .Y(n267) );
  OAI21X1 U15 ( .A0(n198), .A1(n199), .B0(n107), .Y(n270) );
  CLKINVX8 U16 ( .A(n206), .Y(n205) );
  CLKBUFX8 U17 ( .A(n56), .Y(n2) );
  NAND2XL U18 ( .A(B[6]), .B(A[6]), .Y(n56) );
  XOR2X4 U19 ( .A(n202), .B(n204), .Y(SUM[18]) );
  NAND2X2 U20 ( .A(n210), .B(n211), .Y(n190) );
  NOR2BX4 U21 ( .AN(n122), .B(n153), .Y(n152) );
  NAND2X1 U22 ( .A(B[13]), .B(A[13]), .Y(n218) );
  INVX8 U23 ( .A(n239), .Y(n216) );
  CLKBUFX8 U24 ( .A(n218), .Y(n21) );
  XOR2X2 U25 ( .A(n64), .B(n65), .Y(SUM[4]) );
  NAND2X2 U26 ( .A(B[17]), .B(A[17]), .Y(n196) );
  NAND2XL U27 ( .A(B[19]), .B(A[19]), .Y(n182) );
  BUFX3 U28 ( .A(n275), .Y(SUM[5]) );
  OAI21X4 U29 ( .A0(n54), .A1(n55), .B0(n2), .Y(n50) );
  XOR2X4 U30 ( .A(n255), .B(n256), .Y(SUM[11]) );
  OR2X4 U31 ( .A(A[21]), .B(B[21]), .Y(n8) );
  BUFX8 U32 ( .A(n82), .Y(n4) );
  OR2X4 U33 ( .A(A[13]), .B(B[13]), .Y(n239) );
  NOR2X1 U34 ( .A(A[4]), .B(B[4]), .Y(n35) );
  NAND2X4 U35 ( .A(B[4]), .B(A[4]), .Y(n63) );
  BUFX4 U36 ( .A(n274), .Y(SUM[6]) );
  NAND2X2 U37 ( .A(B[24]), .B(A[24]), .Y(n147) );
  NAND2X4 U38 ( .A(n28), .B(n60), .Y(n57) );
  XOR2X2 U39 ( .A(n172), .B(n174), .Y(SUM[20]) );
  NOR2BX2 U40 ( .AN(n171), .B(n175), .Y(n174) );
  NAND3X2 U41 ( .A(n248), .B(n249), .C(n250), .Y(n246) );
  CLKINVX3 U42 ( .A(n188), .Y(n184) );
  AND2X2 U43 ( .A(n117), .B(n118), .Y(n18) );
  INVX2 U44 ( .A(n46), .Y(n244) );
  NAND2BX2 U45 ( .AN(n131), .B(n132), .Y(n130) );
  NAND2X2 U46 ( .A(n61), .B(n27), .Y(n28) );
  INVX2 U47 ( .A(n34), .Y(n27) );
  AOI21X2 U48 ( .A0(n97), .A1(n84), .B0(n98), .Y(n93) );
  INVX1 U49 ( .A(A[20]), .Y(n10) );
  CLKINVX3 U50 ( .A(n253), .Y(n252) );
  INVX1 U51 ( .A(n90), .Y(n86) );
  OR2X2 U52 ( .A(B[18]), .B(A[18]), .Y(n188) );
  NAND2BX2 U53 ( .AN(n53), .B(n261), .Y(n228) );
  NAND3BX1 U54 ( .AN(n34), .B(n263), .C(n59), .Y(n262) );
  NAND2X1 U55 ( .A(n118), .B(n117), .Y(n141) );
  NAND3X1 U56 ( .A(A[24]), .B(B[24]), .C(n117), .Y(n132) );
  CLKINVX3 U57 ( .A(n96), .Y(n81) );
  INVX1 U58 ( .A(n105), .Y(n198) );
  BUFX3 U59 ( .A(n195), .Y(n11) );
  OR2X2 U60 ( .A(A[8]), .B(B[8]), .Y(n254) );
  OR2X2 U61 ( .A(A[3]), .B(B[3]), .Y(n266) );
  OR2X2 U62 ( .A(B[25]), .B(A[25]), .Y(n13) );
  CLKINVX3 U63 ( .A(n118), .Y(n145) );
  INVX4 U64 ( .A(n119), .Y(n154) );
  NOR2X1 U65 ( .A(A[30]), .B(B[30]), .Y(n39) );
  NOR2X2 U66 ( .A(n115), .B(n116), .Y(n114) );
  NAND2X1 U67 ( .A(n96), .B(n99), .Y(n98) );
  XOR2X1 U68 ( .A(B[31]), .B(A[31]), .Y(n75) );
  CLKINVX3 U69 ( .A(n113), .Y(n32) );
  NOR2BX2 U70 ( .AN(n112), .B(n85), .Y(n113) );
  XOR2X1 U71 ( .A(n46), .B(n47), .Y(n273) );
  NOR2BX1 U72 ( .AN(n48), .B(n49), .Y(n47) );
  INVX1 U73 ( .A(n254), .Y(n49) );
  BUFX3 U74 ( .A(n272), .Y(SUM[9]) );
  XOR2X2 U75 ( .A(n257), .B(n259), .Y(SUM[10]) );
  BUFX3 U76 ( .A(n271), .Y(SUM[12]) );
  NOR2BX1 U77 ( .AN(n60), .B(n34), .Y(n62) );
  NOR2BX1 U78 ( .AN(n72), .B(n71), .Y(n103) );
  NOR2BX2 U79 ( .AN(n102), .B(n125), .Y(n124) );
  XOR2X1 U80 ( .A(n57), .B(n58), .Y(n274) );
  OAI2BB1XL U81 ( .A0N(B[28]), .A1N(A[28]), .B0(n4), .Y(n79) );
  NAND2X2 U82 ( .A(n96), .B(n4), .Y(n108) );
  OR2X2 U83 ( .A(A[26]), .B(B[26]), .Y(n89) );
  NOR2X2 U84 ( .A(A[26]), .B(B[26]), .Y(n115) );
  NAND2X1 U85 ( .A(B[9]), .B(A[9]), .Y(n6) );
  NAND2X1 U86 ( .A(B[29]), .B(A[29]), .Y(n82) );
  AND2X2 U87 ( .A(B[26]), .B(A[26]), .Y(n7) );
  NAND2X2 U88 ( .A(A[12]), .B(B[12]), .Y(n217) );
  INVX1 U89 ( .A(n265), .Y(n64) );
  INVX1 U90 ( .A(n8), .Y(n170) );
  INVX1 U91 ( .A(n249), .Y(n45) );
  NAND2BX4 U92 ( .AN(n19), .B(n136), .Y(n150) );
  INVX1 U93 ( .A(n173), .Y(n175) );
  NOR2X2 U94 ( .A(n38), .B(n40), .Y(n212) );
  NOR2BXL U95 ( .AN(n219), .B(n40), .Y(n236) );
  NAND2XL U96 ( .A(n136), .B(n137), .Y(n134) );
  CLKINVX2 U97 ( .A(n137), .Y(n164) );
  INVX1 U98 ( .A(n215), .Y(n214) );
  NAND2X2 U99 ( .A(B[15]), .B(A[15]), .Y(n215) );
  NAND4X4 U100 ( .A(n254), .B(n249), .C(n248), .D(n247), .Y(n220) );
  AOI21X4 U101 ( .A0(n248), .A1(n257), .B0(n258), .Y(n256) );
  NAND3X4 U102 ( .A(n41), .B(n230), .C(n231), .Y(n222) );
  NOR2X2 U103 ( .A(n140), .B(n141), .Y(n128) );
  BUFX8 U104 ( .A(n188), .Y(n9) );
  INVX2 U105 ( .A(n101), .Y(n100) );
  NOR2BXL U106 ( .AN(n52), .B(n53), .Y(n51) );
  NAND2X1 U107 ( .A(B[7]), .B(A[7]), .Y(n52) );
  AOI21X4 U108 ( .A0(B[21]), .A1(A[21]), .B0(n160), .Y(n157) );
  AND2X4 U109 ( .A(n119), .B(n18), .Y(n36) );
  NOR2BX1 U110 ( .AN(n11), .B(n184), .Y(n204) );
  NAND2X2 U111 ( .A(B[20]), .B(A[20]), .Y(n171) );
  NAND2X2 U112 ( .A(B[14]), .B(A[14]), .Y(n219) );
  NOR2BX4 U113 ( .AN(n147), .B(n145), .Y(n155) );
  OAI2BB1X4 U114 ( .A0N(n237), .A1N(n239), .B0(n21), .Y(n235) );
  INVX4 U115 ( .A(n161), .Y(n160) );
  NOR2X2 U116 ( .A(B[27]), .B(A[27]), .Y(n116) );
  AOI21X1 U117 ( .A0(n179), .A1(n180), .B0(n181), .Y(n12) );
  NOR2X4 U118 ( .A(n185), .B(n186), .Y(n179) );
  CLKINVX3 U119 ( .A(n122), .Y(n131) );
  INVX4 U120 ( .A(n182), .Y(n181) );
  OAI2BB1X2 U121 ( .A0N(n120), .A1N(n13), .B0(n121), .Y(n90) );
  NOR2X4 U122 ( .A(n183), .B(n11), .Y(n194) );
  NAND3X4 U123 ( .A(n178), .B(n177), .C(n176), .Y(n14) );
  NAND3XL U124 ( .A(n12), .B(n176), .C(n177), .Y(n172) );
  NAND2X4 U125 ( .A(n208), .B(n186), .Y(n206) );
  NAND2X2 U126 ( .A(B[16]), .B(A[16]), .Y(n186) );
  NAND2X4 U127 ( .A(n210), .B(n211), .Y(n15) );
  OAI2BB1X4 U128 ( .A0N(n165), .A1N(n16), .B0(n161), .Y(n162) );
  CLKINVX20 U129 ( .A(n164), .Y(n16) );
  OR2X4 U130 ( .A(A[17]), .B(B[17]), .Y(n192) );
  NAND2X2 U131 ( .A(B[23]), .B(A[23]), .Y(n135) );
  OR2X2 U132 ( .A(n265), .B(n229), .Y(n29) );
  NOR2X2 U133 ( .A(n149), .B(n148), .Y(n146) );
  NAND3X4 U134 ( .A(n37), .B(n89), .C(n90), .Y(n101) );
  NOR2X4 U135 ( .A(n93), .B(n94), .Y(n92) );
  OAI21X2 U136 ( .A0(n81), .A1(n95), .B0(n4), .Y(n94) );
  CLKINVX4 U137 ( .A(n183), .Y(n17) );
  NAND3X2 U138 ( .A(n101), .B(n102), .C(n84), .Y(n110) );
  XOR2X2 U139 ( .A(n206), .B(n207), .Y(SUM[17]) );
  NAND2X1 U140 ( .A(n60), .B(n63), .Y(n263) );
  NAND2X2 U141 ( .A(B[5]), .B(A[5]), .Y(n60) );
  NOR2BX1 U142 ( .AN(n24), .B(n185), .Y(n207) );
  INVX8 U143 ( .A(n192), .Y(n185) );
  NAND2BX4 U144 ( .AN(n222), .B(n223), .Y(n210) );
  AND2X1 U145 ( .A(n139), .B(n171), .Y(n42) );
  NAND2X2 U146 ( .A(n76), .B(n77), .Y(n74) );
  OAI21X1 U147 ( .A0(n78), .A1(n79), .B0(n80), .Y(n76) );
  INVX4 U148 ( .A(n99), .Y(n85) );
  XOR2X4 U149 ( .A(n50), .B(n51), .Y(SUM[7]) );
  NAND4BX4 U150 ( .AN(n187), .B(n9), .C(n17), .D(n15), .Y(n177) );
  OR2X4 U151 ( .A(A[24]), .B(B[24]), .Y(n118) );
  NAND2X2 U152 ( .A(B[10]), .B(A[10]), .Y(n251) );
  NAND2X2 U153 ( .A(n137), .B(n156), .Y(n19) );
  NAND2X4 U154 ( .A(B[2]), .B(A[2]), .Y(n72) );
  NAND2X4 U155 ( .A(n8), .B(n137), .Y(n138) );
  OAI21X4 U156 ( .A0(n260), .A1(n45), .B0(n6), .Y(n257) );
  INVX2 U157 ( .A(n43), .Y(n260) );
  NOR2BX2 U158 ( .AN(n135), .B(n140), .Y(n163) );
  INVX8 U159 ( .A(n26), .Y(n40) );
  NAND2X1 U160 ( .A(B[26]), .B(A[26]), .Y(n127) );
  NOR2BX4 U161 ( .AN(n161), .B(n164), .Y(n166) );
  BUFX8 U162 ( .A(n110), .Y(n22) );
  NAND2X1 U163 ( .A(n139), .B(n171), .Y(n167) );
  OR2X4 U164 ( .A(A[14]), .B(B[14]), .Y(n26) );
  XOR2X4 U165 ( .A(n91), .B(n92), .Y(SUM[30]) );
  OAI21X4 U166 ( .A0(n145), .A1(n154), .B0(n147), .Y(n151) );
  XOR2X4 U167 ( .A(n74), .B(n75), .Y(SUM[31]) );
  BUFX8 U168 ( .A(n196), .Y(n24) );
  NAND2X2 U169 ( .A(n6), .B(n48), .Y(n250) );
  NAND2X4 U170 ( .A(n30), .B(n48), .Y(n43) );
  NAND2X2 U171 ( .A(B[8]), .B(A[8]), .Y(n48) );
  BUFX4 U172 ( .A(n35), .Y(n25) );
  NAND2X1 U173 ( .A(B[1]), .B(A[1]), .Y(n107) );
  OR2X4 U174 ( .A(A[2]), .B(B[2]), .Y(n104) );
  NOR2X4 U175 ( .A(A[5]), .B(B[5]), .Y(n34) );
  INVX4 U176 ( .A(n57), .Y(n54) );
  XOR2X2 U177 ( .A(n237), .B(n238), .Y(SUM[13]) );
  NAND2X4 U178 ( .A(n29), .B(n228), .Y(n46) );
  NAND4BBX2 U179 ( .AN(n34), .BN(n25), .C(n59), .D(n264), .Y(n229) );
  NAND3BX2 U180 ( .AN(n133), .B(n134), .C(n135), .Y(n129) );
  NOR2BX1 U181 ( .AN(n217), .B(n240), .Y(n243) );
  NAND2X2 U182 ( .A(n46), .B(n254), .Y(n30) );
  OR2X4 U183 ( .A(A[6]), .B(B[6]), .Y(n59) );
  OR2X4 U184 ( .A(A[7]), .B(B[7]), .Y(n264) );
  OR2X2 U185 ( .A(B[12]), .B(A[12]), .Y(n230) );
  OAI2BB1XL U186 ( .A0N(n105), .A1N(n106), .B0(n107), .Y(n73) );
  NAND2XL U187 ( .A(B[0]), .B(A[0]), .Y(n199) );
  NAND2X4 U188 ( .A(n104), .B(n266), .Y(n268) );
  NOR2BX1 U189 ( .AN(n6), .B(n45), .Y(n44) );
  INVX1 U190 ( .A(n112), .Y(n111) );
  XOR2X1 U191 ( .A(n154), .B(n155), .Y(n33) );
  INVX4 U192 ( .A(n33), .Y(SUM[24]) );
  AOI21X4 U193 ( .A0(n9), .A1(n202), .B0(n203), .Y(n201) );
  NOR2BX1 U194 ( .AN(n68), .B(n69), .Y(n67) );
  AOI2BB1X2 U195 ( .A0N(n86), .A1N(n87), .B0(n88), .Y(n83) );
  NAND2XL U196 ( .A(B[30]), .B(A[30]), .Y(n77) );
  INVXL U197 ( .A(n229), .Y(n221) );
  NOR2BXL U198 ( .AN(n2), .B(n55), .Y(n58) );
  AND2X1 U199 ( .A(n251), .B(n248), .Y(n259) );
  NAND3X2 U200 ( .A(n262), .B(n2), .C(n52), .Y(n261) );
  NAND2X2 U201 ( .A(n127), .B(n89), .Y(n142) );
  AND2X1 U202 ( .A(n186), .B(n191), .Y(n209) );
  INVXL U203 ( .A(n11), .Y(n203) );
  NAND2XL U204 ( .A(B[3]), .B(A[3]), .Y(n68) );
  NOR2BXL U205 ( .AN(n107), .B(n198), .Y(n197) );
  OR2X4 U206 ( .A(A[28]), .B(B[28]), .Y(n99) );
  NAND2X4 U207 ( .A(B[27]), .B(A[27]), .Y(n102) );
  OR2X4 U208 ( .A(A[1]), .B(B[1]), .Y(n105) );
  NOR2BX1 U209 ( .AN(n199), .B(n31), .Y(SUM[0]) );
  NOR2XL U210 ( .A(A[0]), .B(B[0]), .Y(n31) );
  OAI21X2 U211 ( .A0(n267), .A1(n268), .B0(n68), .Y(n226) );
  AOI21X2 U212 ( .A0(n221), .A1(n64), .B0(n227), .Y(n224) );
  INVXL U213 ( .A(n228), .Y(n227) );
  INVX1 U214 ( .A(n226), .Y(n265) );
  NAND2BX1 U215 ( .AN(n39), .B(n77), .Y(n91) );
  NOR2BX1 U216 ( .AN(n21), .B(n216), .Y(n238) );
  INVX1 U217 ( .A(n72), .Y(n269) );
  XOR2X1 U218 ( .A(n242), .B(n243), .Y(n271) );
  XOR2X1 U219 ( .A(n61), .B(n62), .Y(n275) );
  XOR2X1 U220 ( .A(n43), .B(n44), .Y(n272) );
  NAND2XL U221 ( .A(n247), .B(n253), .Y(n255) );
  INVX1 U222 ( .A(n251), .Y(n258) );
  XNOR2X4 U223 ( .A(n42), .B(n169), .Y(SUM[21]) );
  NOR2BX1 U224 ( .AN(n63), .B(n25), .Y(n65) );
  INVXL U225 ( .A(n13), .Y(n153) );
  XNOR2X4 U226 ( .A(n22), .B(n32), .Y(SUM[28]) );
  INVX1 U227 ( .A(n59), .Y(n55) );
  INVX1 U228 ( .A(n102), .Y(n88) );
  INVXL U229 ( .A(n156), .Y(n140) );
  INVX1 U230 ( .A(n230), .Y(n240) );
  NOR2X2 U231 ( .A(n88), .B(n100), .Y(n97) );
  NOR2BX2 U232 ( .AN(n251), .B(n252), .Y(n245) );
  INVX1 U233 ( .A(n264), .Y(n53) );
  XOR2X1 U234 ( .A(n66), .B(n67), .Y(SUM[3]) );
  OAI21XL U235 ( .A0(n70), .A1(n71), .B0(n72), .Y(n66) );
  INVX1 U236 ( .A(n73), .Y(n70) );
  XOR2X1 U237 ( .A(n73), .B(n103), .Y(SUM[2]) );
  INVX1 U238 ( .A(n104), .Y(n71) );
  INVX1 U239 ( .A(n266), .Y(n69) );
  NAND2X4 U240 ( .A(n36), .B(n114), .Y(n84) );
  AOI21XL U241 ( .A0(n83), .A1(n84), .B0(n85), .Y(n78) );
  NOR2X1 U242 ( .A(n81), .B(n39), .Y(n80) );
  NAND2XL U243 ( .A(B[28]), .B(A[28]), .Y(n112) );
  NAND2XL U244 ( .A(A[28]), .B(B[28]), .Y(n95) );
  XOR2X1 U245 ( .A(n106), .B(n197), .Y(SUM[1]) );
  INVX1 U246 ( .A(n199), .Y(n106) );
  NAND2X4 U247 ( .A(n190), .B(n191), .Y(n208) );
  NOR2XL U248 ( .A(n138), .B(n139), .Y(n133) );
  NAND2X2 U249 ( .A(B[25]), .B(A[25]), .Y(n122) );
  OR2X2 U250 ( .A(A[9]), .B(B[9]), .Y(n249) );
  NAND2X1 U251 ( .A(B[18]), .B(A[18]), .Y(n195) );
  NAND2X2 U252 ( .A(B[11]), .B(A[11]), .Y(n253) );
  OAI21XL U253 ( .A0(B[27]), .A1(A[27]), .B0(n89), .Y(n87) );
  NOR2X1 U254 ( .A(B[27]), .B(A[27]), .Y(n125) );
  NAND2XL U255 ( .A(B[21]), .B(A[21]), .Y(n168) );
  XOR2X1 U256 ( .A(n190), .B(n209), .Y(SUM[16]) );
  NAND2XL U257 ( .A(n182), .B(n189), .Y(n200) );
  INVX4 U258 ( .A(n242), .Y(n241) );
  AND2X1 U259 ( .A(A[24]), .B(B[24]), .Y(n120) );
  INVX4 U260 ( .A(n235), .Y(n234) );
  INVX8 U261 ( .A(n189), .Y(n183) );
  XOR2X4 U262 ( .A(n108), .B(n109), .Y(SUM[29]) );
  AOI21X4 U263 ( .A0(n22), .A1(n99), .B0(n111), .Y(n109) );
  OR2X4 U264 ( .A(A[29]), .B(B[29]), .Y(n96) );
  NOR2BX4 U265 ( .AN(n122), .B(n7), .Y(n121) );
  XOR2X4 U266 ( .A(n123), .B(n124), .Y(SUM[27]) );
  OAI21X4 U267 ( .A0(n126), .A1(n115), .B0(n127), .Y(n123) );
  AOI21X4 U268 ( .A0(n128), .A1(n129), .B0(n130), .Y(n126) );
  XOR2X4 U269 ( .A(n143), .B(n142), .Y(SUM[26]) );
  AOI21X4 U270 ( .A0(n144), .A1(n13), .B0(n131), .Y(n143) );
  XOR2X4 U271 ( .A(n151), .B(n152), .Y(SUM[25]) );
  OR2X4 U272 ( .A(B[25]), .B(A[25]), .Y(n117) );
  NAND3BX4 U273 ( .AN(n148), .B(n150), .C(n135), .Y(n119) );
  NAND2X4 U274 ( .A(n158), .B(n157), .Y(n136) );
  NOR3BX4 U275 ( .AN(n156), .B(n139), .C(n138), .Y(n148) );
  XOR2X4 U276 ( .A(n162), .B(n163), .Y(SUM[23]) );
  OR2X4 U277 ( .A(A[23]), .B(B[23]), .Y(n156) );
  XOR2X4 U278 ( .A(n165), .B(n166), .Y(SUM[22]) );
  OR2X4 U279 ( .A(B[22]), .B(A[22]), .Y(n137) );
  NAND2X4 U280 ( .A(B[22]), .B(A[22]), .Y(n161) );
  OAI2BB1X4 U281 ( .A0N(n8), .A1N(n167), .B0(n168), .Y(n165) );
  NOR2BX4 U282 ( .AN(n168), .B(n170), .Y(n169) );
  NAND2X4 U283 ( .A(n14), .B(n173), .Y(n139) );
  OR2X4 U284 ( .A(A[20]), .B(B[20]), .Y(n173) );
  AOI21X4 U285 ( .A0(n179), .A1(n180), .B0(n181), .Y(n178) );
  NOR2X4 U286 ( .A(n183), .B(n184), .Y(n180) );
  NAND2X4 U287 ( .A(n191), .B(n192), .Y(n187) );
  AOI21X4 U288 ( .A0(n193), .A1(n9), .B0(n194), .Y(n176) );
  NOR2X4 U289 ( .A(n183), .B(n24), .Y(n193) );
  XOR2X4 U290 ( .A(n200), .B(n201), .Y(SUM[19]) );
  OR2X4 U291 ( .A(B[19]), .B(A[19]), .Y(n189) );
  OAI21X4 U292 ( .A0(n205), .A1(n185), .B0(n24), .Y(n202) );
  AOI21X4 U293 ( .A0(n212), .A1(n213), .B0(n214), .Y(n211) );
  OAI211X2 U294 ( .A0(n216), .A1(n217), .B0(n21), .C0(n219), .Y(n213) );
  NOR2X4 U295 ( .A(n40), .B(n216), .Y(n231) );
  XOR2X4 U296 ( .A(n232), .B(n233), .Y(SUM[15]) );
  OAI21X4 U297 ( .A0(n234), .A1(n40), .B0(n219), .Y(n232) );
  XOR2X4 U298 ( .A(n235), .B(n236), .Y(SUM[14]) );
  OAI21X4 U299 ( .A0(n241), .A1(n240), .B0(n217), .Y(n237) );
  OAI21X4 U300 ( .A0(n244), .A1(n220), .B0(n225), .Y(n242) );
  OAI2BB1X4 U301 ( .A0N(n245), .A1N(n246), .B0(n247), .Y(n225) );
  OR2X4 U302 ( .A(A[11]), .B(B[11]), .Y(n247) );
  OR2X4 U303 ( .A(A[10]), .B(B[10]), .Y(n248) );
endmodule


module hash_core_DW01_add_30 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n236, n237, n1, n2, n3, n4, n5, n6, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235;

  AND2X2 U2 ( .A(n15), .B(n234), .Y(n14) );
  AOI21X2 U3 ( .A0(n26), .A1(n216), .B0(n221), .Y(n223) );
  OR2X4 U4 ( .A(A[1]), .B(B[1]), .Y(n78) );
  NAND2X2 U5 ( .A(B[1]), .B(A[1]), .Y(n80) );
  AOI21X2 U6 ( .A0(n126), .A1(n132), .B0(n133), .Y(n131) );
  NAND2X1 U7 ( .A(B[9]), .B(A[9]), .Y(n28) );
  BUFX8 U8 ( .A(n46), .Y(n1) );
  NAND2XL U9 ( .A(B[5]), .B(A[5]), .Y(n46) );
  XOR2X2 U10 ( .A(n67), .B(n77), .Y(SUM[2]) );
  OAI2BB1X2 U11 ( .A0N(n78), .A1N(n79), .B0(n80), .Y(n67) );
  AOI2BB1XL U12 ( .A0N(n45), .A1N(n1), .B0(n47), .Y(n44) );
  NOR2X2 U13 ( .A(n17), .B(n45), .Y(n235) );
  NOR2BX1 U14 ( .AN(n48), .B(n45), .Y(n52) );
  NOR2X1 U15 ( .A(n17), .B(n45), .Y(n229) );
  CLKINVX3 U16 ( .A(n50), .Y(n45) );
  OR2X4 U17 ( .A(n53), .B(n60), .Y(n10) );
  AOI21X2 U18 ( .A0(n1), .A1(n56), .B0(n53), .Y(n228) );
  INVX2 U19 ( .A(n49), .Y(n53) );
  XOR2X2 U20 ( .A(n30), .B(n31), .Y(SUM[8]) );
  NOR2X2 U21 ( .A(n180), .B(n38), .Y(n204) );
  CLKINVX3 U22 ( .A(n180), .Y(n206) );
  NOR2X2 U23 ( .A(n180), .B(n38), .Y(n183) );
  NAND2X4 U24 ( .A(n214), .B(n215), .Y(n180) );
  OR2X4 U25 ( .A(A[5]), .B(B[5]), .Y(n49) );
  AOI21X1 U26 ( .A0(n183), .A1(n184), .B0(n185), .Y(n181) );
  INVX1 U27 ( .A(n170), .Y(n169) );
  INVX1 U28 ( .A(n153), .Y(n145) );
  NOR2BXL U29 ( .AN(n56), .B(n60), .Y(n59) );
  OAI21XL U30 ( .A0(n16), .A1(n177), .B0(n178), .Y(n175) );
  NOR2X1 U31 ( .A(n33), .B(n29), .Y(n215) );
  OR2X2 U32 ( .A(A[23]), .B(B[23]), .Y(n120) );
  OR2X2 U33 ( .A(A[10]), .B(B[10]), .Y(n220) );
  NAND2X2 U34 ( .A(n232), .B(n233), .Y(n187) );
  AOI21X1 U35 ( .A0(n80), .A1(n159), .B0(n158), .Y(n232) );
  NOR2X1 U36 ( .A(n64), .B(n19), .Y(n233) );
  OR2X2 U37 ( .A(A[3]), .B(B[3]), .Y(n234) );
  INVX1 U38 ( .A(n196), .Y(n176) );
  INVX4 U39 ( .A(n199), .Y(n198) );
  NAND2X1 U40 ( .A(B[8]), .B(A[8]), .Y(n32) );
  INVX1 U41 ( .A(n226), .Y(n33) );
  OAI2BB1X2 U42 ( .A0N(n228), .A1N(n229), .B0(n230), .Y(n37) );
  NAND2X1 U43 ( .A(B[12]), .B(A[12]), .Y(n177) );
  INVX1 U44 ( .A(n22), .Y(n9) );
  NOR2X1 U45 ( .A(A[11]), .B(B[11]), .Y(n18) );
  NAND2X1 U46 ( .A(B[10]), .B(A[10]), .Y(n212) );
  AOI21X2 U47 ( .A0(n26), .A1(n216), .B0(n221), .Y(n219) );
  NOR2X2 U48 ( .A(A[2]), .B(B[2]), .Y(n19) );
  NAND2X1 U49 ( .A(B[3]), .B(A[3]), .Y(n63) );
  INVX1 U50 ( .A(n78), .Y(n158) );
  BUFX3 U51 ( .A(n237), .Y(SUM[9]) );
  BUFX3 U52 ( .A(n236), .Y(SUM[18]) );
  NAND2X1 U53 ( .A(B[7]), .B(A[7]), .Y(n41) );
  OR2X2 U54 ( .A(A[6]), .B(B[6]), .Y(n50) );
  NOR2X2 U55 ( .A(A[7]), .B(B[7]), .Y(n17) );
  XOR2X1 U56 ( .A(n79), .B(n157), .Y(SUM[1]) );
  NOR2BX1 U57 ( .AN(n80), .B(n158), .Y(n157) );
  XOR2X2 U58 ( .A(n102), .B(n103), .Y(SUM[27]) );
  NAND2X4 U59 ( .A(n109), .B(n110), .Y(n88) );
  XOR2X2 U60 ( .A(n35), .B(n59), .Y(SUM[4]) );
  XOR2X4 U61 ( .A(n199), .B(n200), .Y(SUM[13]) );
  OAI2BB1X2 U62 ( .A0N(n9), .A1N(n144), .B0(n155), .Y(n166) );
  OAI2BB1X4 U63 ( .A0N(n224), .A1N(n35), .B0(n225), .Y(n26) );
  NAND2X1 U64 ( .A(B[4]), .B(A[4]), .Y(n56) );
  XOR2X4 U65 ( .A(n193), .B(n194), .Y(SUM[15]) );
  AOI21X1 U66 ( .A0(n37), .A1(n226), .B0(n227), .Y(n225) );
  XOR2X2 U67 ( .A(n130), .B(n131), .Y(SUM[23]) );
  AOI21X2 U68 ( .A0(n174), .A1(n195), .B0(n176), .Y(n194) );
  XOR2X4 U69 ( .A(n160), .B(n161), .Y(SUM[19]) );
  OAI21X2 U70 ( .A0(n162), .A1(n145), .B0(n152), .Y(n160) );
  INVX8 U71 ( .A(n216), .Y(n29) );
  XOR2X2 U72 ( .A(n222), .B(n223), .Y(SUM[10]) );
  NAND2X4 U73 ( .A(n113), .B(n114), .Y(n109) );
  NAND3X4 U74 ( .A(n115), .B(n116), .C(n117), .Y(n114) );
  OAI21X1 U75 ( .A0(n104), .A1(n94), .B0(n93), .Y(n102) );
  INVXL U76 ( .A(n105), .Y(n104) );
  NAND2XL U77 ( .A(n132), .B(n3), .Y(n4) );
  NAND2X2 U78 ( .A(n2), .B(n134), .Y(n5) );
  NAND2X2 U79 ( .A(n4), .B(n5), .Y(SUM[22]) );
  INVXL U80 ( .A(n132), .Y(n2) );
  INVX1 U81 ( .A(n134), .Y(n3) );
  OAI21X4 U82 ( .A0(n135), .A1(n23), .B0(n129), .Y(n132) );
  OR2X4 U83 ( .A(n219), .B(n213), .Y(n6) );
  NAND2X4 U84 ( .A(n6), .B(n212), .Y(n217) );
  OAI2BB1X4 U85 ( .A0N(n204), .A1N(n35), .B0(n205), .Y(n202) );
  AOI21X2 U86 ( .A0(n206), .A1(n37), .B0(n185), .Y(n205) );
  OAI21X4 U87 ( .A0(n165), .A1(n20), .B0(n156), .Y(n163) );
  INVX4 U88 ( .A(n136), .Y(n135) );
  OAI21X4 U89 ( .A0(n24), .A1(n138), .B0(n128), .Y(n136) );
  XOR2X4 U90 ( .A(n217), .B(n218), .Y(SUM[11]) );
  NAND2X4 U91 ( .A(B[2]), .B(A[2]), .Y(n66) );
  NOR2X2 U92 ( .A(A[13]), .B(B[13]), .Y(n16) );
  NAND2XL U93 ( .A(B[13]), .B(A[13]), .Y(n178) );
  NOR2X2 U94 ( .A(n213), .B(n18), .Y(n214) );
  NOR2BX2 U95 ( .AN(n63), .B(n64), .Y(n62) );
  XNOR2X1 U96 ( .A(n71), .B(n11), .Y(SUM[30]) );
  OR2X4 U97 ( .A(A[4]), .B(B[4]), .Y(n54) );
  NAND2XL U98 ( .A(B[17]), .B(A[17]), .Y(n156) );
  NOR2XL U99 ( .A(n188), .B(n14), .Y(n186) );
  XOR2X2 U100 ( .A(n61), .B(n62), .Y(SUM[3]) );
  OAI21X4 U101 ( .A0(n42), .A1(n53), .B0(n1), .Y(n51) );
  AOI21X1 U102 ( .A0(n174), .A1(n175), .B0(n176), .Y(n171) );
  XOR2X1 U103 ( .A(n26), .B(n27), .Y(n237) );
  NAND2XL U104 ( .A(n49), .B(n1), .Y(n57) );
  INVX4 U105 ( .A(n202), .Y(n201) );
  INVX2 U106 ( .A(n220), .Y(n213) );
  NOR2X1 U107 ( .A(A[17]), .B(B[17]), .Y(n20) );
  NAND2XL U108 ( .A(B[6]), .B(A[6]), .Y(n48) );
  NAND2X1 U109 ( .A(B[24]), .B(A[24]), .Y(n97) );
  OR2X2 U110 ( .A(A[22]), .B(B[22]), .Y(n126) );
  OAI21X4 U111 ( .A0(n179), .A1(n13), .B0(n169), .Y(n144) );
  NAND2BXL U112 ( .AN(n180), .B(n37), .Y(n182) );
  INVXL U113 ( .A(n37), .Y(n36) );
  OAI21X2 U114 ( .A0(n65), .A1(n19), .B0(n66), .Y(n61) );
  INVX2 U115 ( .A(n67), .Y(n65) );
  NOR2BXL U116 ( .AN(n125), .B(n118), .Y(n134) );
  NAND2XL U117 ( .A(n123), .B(n120), .Y(n130) );
  INVXL U118 ( .A(n125), .Y(n133) );
  NOR2BXL U119 ( .AN(n98), .B(n96), .Y(n108) );
  NAND2X2 U120 ( .A(n140), .B(n141), .Y(n117) );
  OAI2BB1X2 U121 ( .A0N(n101), .A1N(n107), .B0(n98), .Y(n105) );
  AOI2BB1X2 U122 ( .A0N(n17), .A1N(n48), .B0(n231), .Y(n230) );
  NAND2BX4 U123 ( .AN(n10), .B(n235), .Y(n38) );
  NOR2BXL U124 ( .AN(n150), .B(n146), .Y(n161) );
  XOR2X4 U125 ( .A(n57), .B(n58), .Y(SUM[5]) );
  INVX1 U126 ( .A(n66), .Y(n15) );
  NOR2BXL U127 ( .AN(n28), .B(n29), .Y(n27) );
  NOR2BX1 U128 ( .AN(n99), .B(n91), .Y(n90) );
  NAND2X1 U129 ( .A(n69), .B(n72), .Y(n11) );
  NOR2BXL U130 ( .AN(n129), .B(n23), .Y(n137) );
  XOR2X2 U131 ( .A(n202), .B(n203), .Y(SUM[12]) );
  XOR2XL U132 ( .A(n81), .B(n74), .Y(SUM[29]) );
  NAND2XL U133 ( .A(n173), .B(n192), .Y(n193) );
  NOR2XL U134 ( .A(n38), .B(n33), .Y(n224) );
  NAND2XL U135 ( .A(n71), .B(n72), .Y(n70) );
  NOR2XL U136 ( .A(n23), .B(n24), .Y(n116) );
  NAND2X4 U137 ( .A(B[0]), .B(A[0]), .Y(n159) );
  NOR2BX1 U138 ( .AN(n159), .B(n12), .Y(SUM[0]) );
  NOR2XL U139 ( .A(A[0]), .B(B[0]), .Y(n12) );
  OR2X4 U140 ( .A(A[9]), .B(B[9]), .Y(n216) );
  NOR2XL U141 ( .A(A[12]), .B(B[12]), .Y(n21) );
  NAND2XL U142 ( .A(B[18]), .B(A[18]), .Y(n152) );
  NAND2XL U143 ( .A(B[11]), .B(A[11]), .Y(n208) );
  NAND2XL U144 ( .A(B[15]), .B(A[15]), .Y(n173) );
  NOR2XL U145 ( .A(A[16]), .B(B[16]), .Y(n22) );
  NAND2XL U146 ( .A(B[21]), .B(A[21]), .Y(n129) );
  NAND2XL U147 ( .A(B[19]), .B(A[19]), .Y(n150) );
  NOR2XL U148 ( .A(A[20]), .B(B[20]), .Y(n24) );
  NAND2XL U149 ( .A(B[25]), .B(A[25]), .Y(n98) );
  AND2X2 U150 ( .A(n181), .B(n182), .Y(n13) );
  NAND2XL U151 ( .A(n186), .B(n187), .Y(n184) );
  NOR2X1 U152 ( .A(n29), .B(n213), .Y(n209) );
  NOR2X1 U153 ( .A(n145), .B(n146), .Y(n142) );
  NOR2BX1 U154 ( .AN(n178), .B(n16), .Y(n200) );
  NOR2BX1 U155 ( .AN(n208), .B(n18), .Y(n218) );
  INVX1 U156 ( .A(n56), .Y(n55) );
  OAI21X2 U157 ( .A0(n207), .A1(n18), .B0(n208), .Y(n185) );
  AOI21X1 U158 ( .A0(n209), .A1(n210), .B0(n211), .Y(n207) );
  INVX1 U159 ( .A(n212), .Y(n211) );
  NAND2X1 U160 ( .A(n28), .B(n32), .Y(n210) );
  XOR2X1 U161 ( .A(n163), .B(n164), .Y(n236) );
  NOR2BX1 U162 ( .AN(n152), .B(n145), .Y(n164) );
  INVX1 U163 ( .A(n166), .Y(n165) );
  INVX1 U164 ( .A(n117), .Y(n138) );
  INVX1 U165 ( .A(n32), .Y(n227) );
  NOR2BX1 U166 ( .AN(n196), .B(n191), .Y(n197) );
  INVX1 U167 ( .A(n54), .Y(n60) );
  INVX1 U168 ( .A(n174), .Y(n191) );
  NOR2BX1 U169 ( .AN(n41), .B(n17), .Y(n40) );
  OAI21X2 U170 ( .A0(n42), .A1(n43), .B0(n44), .Y(n39) );
  NAND2X1 U171 ( .A(n49), .B(n50), .Y(n43) );
  XOR2X1 U172 ( .A(n166), .B(n167), .Y(SUM[17]) );
  NOR2BX1 U173 ( .AN(n156), .B(n20), .Y(n167) );
  INVX1 U174 ( .A(n163), .Y(n162) );
  NOR2BX1 U175 ( .AN(n32), .B(n33), .Y(n31) );
  OAI2BB1X1 U176 ( .A0N(n34), .A1N(n35), .B0(n36), .Y(n30) );
  INVX1 U177 ( .A(n38), .Y(n34) );
  NOR2BX1 U178 ( .AN(n66), .B(n19), .Y(n77) );
  NOR2BX1 U179 ( .AN(n177), .B(n21), .Y(n203) );
  OAI21XL U180 ( .A0(n171), .A1(n172), .B0(n173), .Y(n170) );
  NAND2X1 U181 ( .A(n212), .B(n220), .Y(n222) );
  AOI21X1 U182 ( .A0(n147), .A1(n148), .B0(n149), .Y(n140) );
  NAND3X1 U183 ( .A(n142), .B(n143), .C(n144), .Y(n141) );
  INVX1 U184 ( .A(n150), .Y(n149) );
  INVX1 U185 ( .A(n48), .Y(n47) );
  INVX1 U186 ( .A(n159), .Y(n79) );
  INVX1 U187 ( .A(n41), .Y(n231) );
  NAND2X1 U188 ( .A(n189), .B(n190), .Y(n179) );
  NOR2X1 U189 ( .A(n172), .B(n191), .Y(n190) );
  NOR2X1 U190 ( .A(n16), .B(n21), .Y(n189) );
  OAI21XL U191 ( .A0(n88), .A1(n89), .B0(n90), .Y(n82) );
  NAND3BX1 U192 ( .AN(n25), .B(n100), .C(n101), .Y(n89) );
  XOR2X1 U193 ( .A(n105), .B(n106), .Y(SUM[26]) );
  NOR2BX1 U194 ( .AN(n93), .B(n94), .Y(n106) );
  INVX1 U195 ( .A(n192), .Y(n172) );
  INVX1 U196 ( .A(n28), .Y(n221) );
  INVX1 U197 ( .A(n148), .Y(n146) );
  XOR2X1 U198 ( .A(n82), .B(n86), .Y(SUM[28]) );
  NOR2BX1 U199 ( .AN(n85), .B(n87), .Y(n86) );
  INVX1 U200 ( .A(n83), .Y(n87) );
  XOR2X1 U201 ( .A(n136), .B(n137), .Y(SUM[21]) );
  XOR2X1 U202 ( .A(n117), .B(n139), .Y(SUM[20]) );
  NOR2BX1 U203 ( .AN(n128), .B(n24), .Y(n139) );
  XOR2X1 U204 ( .A(n144), .B(n168), .Y(SUM[16]) );
  NOR2BX1 U205 ( .AN(n155), .B(n22), .Y(n168) );
  NOR2BX1 U206 ( .AN(n99), .B(n25), .Y(n103) );
  XOR2X1 U207 ( .A(n109), .B(n111), .Y(SUM[24]) );
  NOR2BX1 U208 ( .AN(n97), .B(n112), .Y(n111) );
  INVX1 U209 ( .A(n110), .Y(n112) );
  XOR2X1 U210 ( .A(n107), .B(n108), .Y(SUM[25]) );
  AOI21X1 U211 ( .A0(n121), .A1(n120), .B0(n122), .Y(n113) );
  INVX1 U212 ( .A(n123), .Y(n122) );
  NOR2X1 U213 ( .A(n20), .B(n22), .Y(n143) );
  NAND2X1 U214 ( .A(n88), .B(n97), .Y(n107) );
  NAND2X1 U215 ( .A(n151), .B(n152), .Y(n147) );
  NAND2X1 U216 ( .A(n153), .B(n154), .Y(n151) );
  OAI21XL U217 ( .A0(n20), .A1(n155), .B0(n156), .Y(n154) );
  INVX1 U218 ( .A(n63), .Y(n188) );
  AOI21X1 U219 ( .A0(n82), .A1(n83), .B0(n84), .Y(n74) );
  INVX1 U220 ( .A(n85), .Y(n84) );
  OAI21XL U221 ( .A0(n73), .A1(n74), .B0(n75), .Y(n71) );
  INVX1 U222 ( .A(n76), .Y(n73) );
  INVX1 U223 ( .A(n126), .Y(n118) );
  NAND2X1 U224 ( .A(n124), .B(n125), .Y(n121) );
  NAND2X1 U225 ( .A(n126), .B(n127), .Y(n124) );
  OAI21XL U226 ( .A0(n23), .A1(n128), .B0(n129), .Y(n127) );
  NAND2X1 U227 ( .A(n75), .B(n76), .Y(n81) );
  NOR2X1 U228 ( .A(n118), .B(n119), .Y(n115) );
  INVX1 U229 ( .A(n120), .Y(n119) );
  NAND2X1 U230 ( .A(n69), .B(n70), .Y(n68) );
  INVX1 U231 ( .A(n100), .Y(n94) );
  INVX1 U232 ( .A(n101), .Y(n96) );
  AOI21X1 U233 ( .A0(n92), .A1(n93), .B0(n25), .Y(n91) );
  NAND2BX1 U234 ( .AN(n94), .B(n95), .Y(n92) );
  OAI21XL U235 ( .A0(n96), .A1(n97), .B0(n98), .Y(n95) );
  XOR3X2 U236 ( .A(B[31]), .B(A[31]), .C(n68), .Y(SUM[31]) );
  OR2X2 U237 ( .A(A[14]), .B(B[14]), .Y(n174) );
  NAND2X1 U238 ( .A(B[14]), .B(A[14]), .Y(n196) );
  OR2X2 U239 ( .A(A[8]), .B(B[8]), .Y(n226) );
  NAND2X1 U240 ( .A(B[16]), .B(A[16]), .Y(n155) );
  OR2X2 U241 ( .A(A[19]), .B(B[19]), .Y(n148) );
  OR2X2 U242 ( .A(A[18]), .B(B[18]), .Y(n153) );
  OR2X2 U243 ( .A(A[15]), .B(B[15]), .Y(n192) );
  NOR2X1 U244 ( .A(A[21]), .B(B[21]), .Y(n23) );
  NAND2X1 U245 ( .A(B[20]), .B(A[20]), .Y(n128) );
  NAND2X1 U246 ( .A(B[22]), .B(A[22]), .Y(n125) );
  NAND2X1 U247 ( .A(B[23]), .B(A[23]), .Y(n123) );
  OR2X2 U248 ( .A(A[24]), .B(B[24]), .Y(n110) );
  NOR2X1 U249 ( .A(A[27]), .B(B[27]), .Y(n25) );
  NAND2X1 U250 ( .A(B[26]), .B(A[26]), .Y(n93) );
  OR2X2 U251 ( .A(A[25]), .B(B[25]), .Y(n101) );
  NAND2X1 U252 ( .A(B[27]), .B(A[27]), .Y(n99) );
  OR2X2 U253 ( .A(A[28]), .B(B[28]), .Y(n83) );
  OR2X2 U254 ( .A(A[26]), .B(B[26]), .Y(n100) );
  NAND2X1 U255 ( .A(B[29]), .B(A[29]), .Y(n75) );
  NAND2X1 U256 ( .A(B[28]), .B(A[28]), .Y(n85) );
  OR2X2 U257 ( .A(A[30]), .B(B[30]), .Y(n72) );
  OR2X2 U258 ( .A(A[29]), .B(B[29]), .Y(n76) );
  NAND2X1 U259 ( .A(B[30]), .B(A[30]), .Y(n69) );
  NAND3BX4 U260 ( .AN(n14), .B(n63), .C(n187), .Y(n35) );
  XOR2X4 U261 ( .A(n39), .B(n40), .Y(SUM[7]) );
  XOR2X4 U262 ( .A(n51), .B(n52), .Y(SUM[6]) );
  AOI21X4 U263 ( .A0(n35), .A1(n54), .B0(n55), .Y(n42) );
  AOI21X4 U264 ( .A0(n35), .A1(n54), .B0(n55), .Y(n58) );
  XOR2X4 U265 ( .A(n195), .B(n197), .Y(SUM[14]) );
  OAI21X4 U266 ( .A0(n198), .A1(n16), .B0(n178), .Y(n195) );
  OAI21X4 U267 ( .A0(n21), .A1(n201), .B0(n177), .Y(n199) );
  CLKINVX3 U268 ( .A(n234), .Y(n64) );
endmodule


module hash_core_DW01_add_32 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n273, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272;

  NAND2X4 U2 ( .A(n65), .B(n62), .Y(n64) );
  NAND3BX4 U3 ( .AN(n54), .B(n55), .C(n35), .Y(n53) );
  NAND2X4 U4 ( .A(n55), .B(n35), .Y(n77) );
  BUFX16 U5 ( .A(n56), .Y(n35) );
  NAND2X2 U6 ( .A(n251), .B(n42), .Y(n259) );
  OAI21X4 U7 ( .A0(n4), .A1(n140), .B0(n139), .Y(n148) );
  OAI21X2 U8 ( .A0(n207), .A1(n208), .B0(n209), .Y(n204) );
  CLKINVX8 U9 ( .A(n101), .Y(n87) );
  NAND2X1 U10 ( .A(B[14]), .B(A[14]), .Y(n206) );
  OAI2BB1X4 U11 ( .A0N(n172), .A1N(n180), .B0(n169), .Y(n178) );
  NOR2X4 U12 ( .A(n267), .B(n63), .Y(n265) );
  INVX4 U13 ( .A(n49), .Y(n267) );
  NAND3X2 U14 ( .A(n264), .B(n265), .C(n266), .Y(n210) );
  INVX4 U15 ( .A(n75), .Y(n14) );
  INVX8 U16 ( .A(n47), .Y(n230) );
  INVXL U17 ( .A(n86), .Y(n174) );
  NOR2X4 U18 ( .A(n39), .B(n248), .Y(n242) );
  INVX12 U19 ( .A(n251), .Y(n39) );
  AOI21X1 U20 ( .A0(n46), .A1(n35), .B0(n198), .Y(n263) );
  CLKINVX8 U21 ( .A(n191), .Y(n46) );
  AOI21X1 U22 ( .A0(n197), .A1(n198), .B0(n199), .Y(n187) );
  OAI2BB1X4 U23 ( .A0N(n198), .A1N(n31), .B0(n260), .Y(n256) );
  BUFX3 U24 ( .A(n273), .Y(SUM[25]) );
  NAND2X4 U25 ( .A(n210), .B(n50), .Y(n198) );
  XOR2X4 U26 ( .A(n239), .B(n240), .Y(SUM[12]) );
  NOR2X2 U27 ( .A(n193), .B(n192), .Y(n197) );
  XOR2X2 U28 ( .A(n180), .B(n181), .Y(SUM[17]) );
  NAND2X2 U29 ( .A(n4), .B(n151), .Y(n7) );
  INVX1 U30 ( .A(n151), .Y(n5) );
  INVX1 U31 ( .A(n170), .Y(n161) );
  INVX2 U32 ( .A(n198), .Y(n252) );
  OR2X2 U33 ( .A(A[25]), .B(B[25]), .Y(n110) );
  INVX1 U34 ( .A(n146), .Y(n140) );
  NAND2XL U35 ( .A(n202), .B(n218), .Y(n220) );
  NOR2BXL U36 ( .AN(n164), .B(n165), .Y(n179) );
  NOR2BXL U37 ( .AN(n144), .B(n142), .Y(n154) );
  NAND2BX1 U38 ( .AN(n45), .B(n46), .Y(n40) );
  NAND2X2 U39 ( .A(n215), .B(n216), .Y(n192) );
  INVX1 U40 ( .A(n208), .Y(n235) );
  OAI21X2 U41 ( .A0(n200), .A1(n201), .B0(n202), .Y(n199) );
  INVX1 U42 ( .A(n206), .Y(n205) );
  NOR2BX1 U43 ( .AN(n74), .B(n195), .Y(n194) );
  INVX1 U44 ( .A(n192), .Y(n212) );
  NAND3BX1 U45 ( .AN(n33), .B(n171), .C(n172), .Y(n160) );
  OR2X2 U46 ( .A(n161), .B(n162), .Y(n28) );
  OAI21XL U47 ( .A0(n142), .A1(n143), .B0(n144), .Y(n141) );
  OR2X2 U48 ( .A(A[21]), .B(B[21]), .Y(n147) );
  NAND2X2 U49 ( .A(n69), .B(n18), .Y(n264) );
  NAND3X2 U50 ( .A(n62), .B(n18), .C(n57), .Y(n266) );
  OR2X2 U51 ( .A(A[9]), .B(B[9]), .Y(n251) );
  NOR2X1 U52 ( .A(A[19]), .B(B[19]), .Y(n33) );
  CLKINVX3 U53 ( .A(n59), .Y(n63) );
  INVX1 U54 ( .A(n89), .Y(n88) );
  INVX1 U55 ( .A(n229), .Y(n3) );
  NOR2BX1 U56 ( .AN(n209), .B(n207), .Y(n229) );
  NOR2BX1 U57 ( .AN(n208), .B(n219), .Y(n240) );
  NAND2X1 U58 ( .A(n115), .B(n111), .Y(n122) );
  NAND2X1 U59 ( .A(n110), .B(n127), .Y(n126) );
  XOR2X2 U60 ( .A(n148), .B(n149), .Y(SUM[23]) );
  OR2X2 U61 ( .A(A[7]), .B(B[7]), .Y(n49) );
  INVX1 U62 ( .A(n76), .Y(n15) );
  AND2X2 U63 ( .A(n100), .B(n89), .Y(n30) );
  OAI21X2 U64 ( .A0(n66), .A1(n67), .B0(n68), .Y(n65) );
  INVX4 U65 ( .A(n72), .Y(n270) );
  CLKINVX3 U66 ( .A(n150), .Y(n4) );
  NAND2X1 U67 ( .A(B[13]), .B(A[13]), .Y(n209) );
  NAND2X1 U68 ( .A(n85), .B(n84), .Y(n99) );
  NOR2X2 U69 ( .A(n69), .B(n70), .Y(n68) );
  NAND3X1 U70 ( .A(n2), .B(n87), .C(n86), .Y(n100) );
  OR2XL U71 ( .A(A[0]), .B(B[0]), .Y(n2) );
  OAI21X2 U72 ( .A0(n263), .A1(n259), .B0(n260), .Y(n261) );
  INVX1 U73 ( .A(n259), .Y(n31) );
  NAND2X4 U74 ( .A(n109), .B(n120), .Y(n127) );
  NAND2X4 U75 ( .A(n129), .B(n130), .Y(n109) );
  INVXL U76 ( .A(n44), .Y(n43) );
  OAI2BB1X1 U77 ( .A0N(n38), .A1N(n44), .B0(n251), .Y(n260) );
  NAND2X1 U78 ( .A(n38), .B(n44), .Y(n243) );
  NAND2X1 U79 ( .A(B[8]), .B(A[8]), .Y(n44) );
  NOR2BX4 U80 ( .AN(n74), .B(n81), .Y(n80) );
  AOI21X2 U81 ( .A0(n227), .A1(n223), .B0(n228), .Y(n226) );
  AOI21X2 U82 ( .A0(n222), .A1(n223), .B0(n224), .Y(n221) );
  NAND2X4 U83 ( .A(B[1]), .B(A[1]), .Y(n89) );
  NOR3BX4 U84 ( .AN(n35), .B(n259), .C(n191), .Y(n257) );
  AND2X4 U85 ( .A(n86), .B(n87), .Y(n13) );
  OAI21X4 U86 ( .A0(n230), .A1(n193), .B0(n213), .Y(n239) );
  CLKINVX4 U87 ( .A(n73), .Y(n195) );
  AOI21X1 U88 ( .A0(n198), .A1(n42), .B0(n43), .Y(n41) );
  INVX4 U89 ( .A(n196), .Y(n71) );
  AOI2BB1X2 U90 ( .A0N(n233), .A1N(n234), .B0(n235), .Y(n232) );
  INVX4 U91 ( .A(n35), .Y(n78) );
  XNOR2X4 U92 ( .A(n223), .B(n3), .Y(SUM[13]) );
  NOR3X2 U93 ( .A(n191), .B(n192), .C(n193), .Y(n190) );
  XOR2X4 U94 ( .A(n153), .B(n154), .Y(SUM[21]) );
  NAND2X2 U95 ( .A(n150), .B(n5), .Y(n6) );
  NAND2X4 U96 ( .A(n6), .B(n7), .Y(SUM[22]) );
  NAND2X4 U97 ( .A(n122), .B(n9), .Y(n10) );
  NAND2X1 U98 ( .A(n8), .B(n123), .Y(n11) );
  NAND2X4 U99 ( .A(n10), .B(n11), .Y(SUM[27]) );
  INVXL U100 ( .A(n122), .Y(n8) );
  INVX2 U101 ( .A(n123), .Y(n9) );
  AOI21X2 U102 ( .A0(n112), .A1(n124), .B0(n125), .Y(n123) );
  OR2X4 U103 ( .A(n256), .B(n257), .Y(n12) );
  NAND2X4 U104 ( .A(n12), .B(n258), .Y(n255) );
  NOR2X4 U105 ( .A(n13), .B(n88), .Y(n82) );
  OAI21X4 U106 ( .A0(n82), .A1(n83), .B0(n84), .Y(n79) );
  NAND2X2 U107 ( .A(n75), .B(n76), .Y(n16) );
  NAND2X4 U108 ( .A(n14), .B(n15), .Y(n17) );
  NAND2X4 U109 ( .A(n17), .B(n16), .Y(SUM[5]) );
  NAND2X4 U110 ( .A(n77), .B(n57), .Y(n75) );
  BUFX8 U111 ( .A(n60), .Y(n18) );
  AND3X4 U112 ( .A(n51), .B(n52), .C(n53), .Y(n29) );
  AOI21X2 U113 ( .A0(n203), .A1(n204), .B0(n205), .Y(n200) );
  NAND2X4 U114 ( .A(B[12]), .B(A[12]), .Y(n208) );
  OAI21XL U115 ( .A0(n217), .A1(n209), .B0(n206), .Y(n224) );
  NOR2BX2 U116 ( .AN(n101), .B(n26), .Y(SUM[0]) );
  NAND2X4 U117 ( .A(n133), .B(n143), .Y(n153) );
  OAI21X4 U118 ( .A0(n133), .A1(n134), .B0(n135), .Y(n129) );
  XNOR2X2 U119 ( .A(n124), .B(n20), .Y(SUM[26]) );
  CLKINVX8 U120 ( .A(n27), .Y(n155) );
  XOR2XL U121 ( .A(n102), .B(n96), .Y(SUM[29]) );
  NAND2X2 U122 ( .A(B[5]), .B(A[5]), .Y(n62) );
  NAND2X2 U123 ( .A(B[20]), .B(A[20]), .Y(n143) );
  OR2XL U124 ( .A(A[20]), .B(B[20]), .Y(n156) );
  AOI2BB1X4 U125 ( .A0N(n159), .A1N(n160), .B0(n28), .Y(n27) );
  NAND2X1 U126 ( .A(n117), .B(n112), .Y(n20) );
  INVXL U127 ( .A(n178), .Y(n177) );
  NOR2BXL U128 ( .AN(n170), .B(n33), .Y(n176) );
  NAND2XL U129 ( .A(B[18]), .B(A[18]), .Y(n164) );
  NAND2X1 U130 ( .A(B[17]), .B(A[17]), .Y(n169) );
  NAND2X1 U131 ( .A(B[21]), .B(A[21]), .Y(n144) );
  NAND2X1 U132 ( .A(B[24]), .B(A[24]), .Y(n120) );
  NAND2X1 U133 ( .A(B[25]), .B(A[25]), .Y(n121) );
  NOR2X4 U134 ( .A(n69), .B(n70), .Y(n271) );
  NOR2X4 U135 ( .A(n267), .B(n63), .Y(n272) );
  NAND2X2 U136 ( .A(n189), .B(n190), .Y(n188) );
  XOR2X4 U137 ( .A(n78), .B(n19), .Y(SUM[4]) );
  NAND2XL U138 ( .A(n57), .B(n55), .Y(n19) );
  NAND3BXL U139 ( .AN(n34), .B(n146), .C(n147), .Y(n134) );
  INVXL U140 ( .A(n117), .Y(n125) );
  NAND2X2 U141 ( .A(n126), .B(n121), .Y(n124) );
  NAND2X4 U142 ( .A(n155), .B(n156), .Y(n133) );
  OAI21X1 U143 ( .A0(n167), .A1(n168), .B0(n169), .Y(n166) );
  NOR2BX2 U144 ( .AN(n245), .B(n246), .Y(n244) );
  XOR2X2 U145 ( .A(n93), .B(n32), .Y(SUM[30]) );
  XNOR2X1 U146 ( .A(n103), .B(n22), .Y(SUM[28]) );
  NAND2X1 U147 ( .A(n106), .B(n104), .Y(n22) );
  NOR2BXL U148 ( .AN(n169), .B(n167), .Y(n181) );
  XNOR2X4 U149 ( .A(n29), .B(n23), .Y(SUM[7]) );
  AND2X1 U150 ( .A(n49), .B(n50), .Y(n23) );
  AND2X1 U151 ( .A(n247), .B(n236), .Y(n24) );
  XOR2X4 U152 ( .A(n178), .B(n179), .Y(SUM[18]) );
  AND2X1 U153 ( .A(n18), .B(n59), .Y(n25) );
  NOR2BXL U154 ( .AN(n145), .B(n34), .Y(n149) );
  INVXL U155 ( .A(n245), .Y(n254) );
  NAND2XL U156 ( .A(n93), .B(n94), .Y(n92) );
  NAND2X4 U157 ( .A(B[0]), .B(A[0]), .Y(n101) );
  NOR2XL U158 ( .A(A[0]), .B(B[0]), .Y(n26) );
  NAND2X2 U159 ( .A(B[16]), .B(A[16]), .Y(n168) );
  NAND2X1 U160 ( .A(B[6]), .B(A[6]), .Y(n60) );
  OR2X4 U161 ( .A(A[17]), .B(B[17]), .Y(n172) );
  OR2X4 U162 ( .A(A[18]), .B(B[18]), .Y(n171) );
  NAND2XL U163 ( .A(B[22]), .B(A[22]), .Y(n139) );
  NAND2XL U164 ( .A(B[19]), .B(A[19]), .Y(n170) );
  OR2XL U165 ( .A(A[16]), .B(B[16]), .Y(n183) );
  NAND2XL U166 ( .A(B[23]), .B(A[23]), .Y(n145) );
  NAND2BX1 U167 ( .AN(n219), .B(n214), .Y(n231) );
  INVXL U168 ( .A(n193), .Y(n214) );
  NOR2XL U169 ( .A(n207), .B(n217), .Y(n222) );
  INVXL U170 ( .A(n238), .Y(n233) );
  NAND2XL U171 ( .A(n206), .B(n203), .Y(n225) );
  INVX1 U172 ( .A(n209), .Y(n228) );
  OAI21XL U173 ( .A0(n71), .A1(n72), .B0(n194), .Y(n189) );
  NOR2X1 U174 ( .A(n136), .B(n137), .Y(n135) );
  INVX1 U175 ( .A(n145), .Y(n136) );
  INVX1 U176 ( .A(n171), .Y(n165) );
  INVX1 U177 ( .A(n172), .Y(n167) );
  NOR2BXL U178 ( .AN(n44), .B(n45), .Y(n48) );
  NOR2BXL U179 ( .AN(n38), .B(n39), .Y(n37) );
  XOR2X1 U180 ( .A(n155), .B(n157), .Y(SUM[20]) );
  NOR2BX1 U181 ( .AN(n143), .B(n158), .Y(n157) );
  INVX1 U182 ( .A(n156), .Y(n158) );
  XOR2X1 U183 ( .A(n182), .B(n184), .Y(SUM[16]) );
  NOR2BX1 U184 ( .AN(n168), .B(n185), .Y(n184) );
  INVX1 U185 ( .A(n183), .Y(n185) );
  NOR2BXL U186 ( .AN(n245), .B(n248), .Y(n262) );
  XOR2X1 U187 ( .A(n127), .B(n128), .Y(n273) );
  NOR2BX1 U188 ( .AN(n121), .B(n119), .Y(n128) );
  NOR2BX1 U189 ( .AN(n139), .B(n140), .Y(n151) );
  XNOR2X4 U190 ( .A(n101), .B(n173), .Y(SUM[1]) );
  XOR2X4 U191 ( .A(n30), .B(n99), .Y(SUM[2]) );
  NAND2XL U192 ( .A(n57), .B(n74), .Y(n66) );
  AOI21X1 U193 ( .A0(n163), .A1(n164), .B0(n33), .Y(n162) );
  NAND2BX1 U194 ( .AN(n165), .B(n166), .Y(n163) );
  INVXL U195 ( .A(n269), .Y(n81) );
  NOR2BX1 U196 ( .AN(n18), .B(n61), .Y(n51) );
  NOR2XL U197 ( .A(n62), .B(n63), .Y(n61) );
  NAND2XL U198 ( .A(n58), .B(n59), .Y(n54) );
  INVXL U199 ( .A(n85), .Y(n83) );
  INVX1 U200 ( .A(n247), .Y(n246) );
  OR2XL U201 ( .A(n54), .B(n57), .Y(n52) );
  NAND2XL U202 ( .A(n58), .B(n62), .Y(n76) );
  NAND2XL U203 ( .A(n236), .B(n237), .Y(n234) );
  AOI21X1 U204 ( .A0(n103), .A1(n104), .B0(n105), .Y(n96) );
  INVX1 U205 ( .A(n106), .Y(n105) );
  OAI21XL U206 ( .A0(n95), .A1(n96), .B0(n97), .Y(n93) );
  INVX1 U207 ( .A(n98), .Y(n95) );
  INVX1 U208 ( .A(n147), .Y(n142) );
  XOR2X1 U209 ( .A(n129), .B(n131), .Y(SUM[24]) );
  NOR2BX1 U210 ( .AN(n120), .B(n132), .Y(n131) );
  INVX1 U211 ( .A(n130), .Y(n132) );
  NAND2X1 U212 ( .A(n97), .B(n98), .Y(n102) );
  NAND2X1 U213 ( .A(n107), .B(n108), .Y(n103) );
  AOI21X1 U214 ( .A0(n113), .A1(n111), .B0(n114), .Y(n107) );
  NAND4BXL U215 ( .AN(n109), .B(n110), .C(n111), .D(n112), .Y(n108) );
  INVX1 U216 ( .A(n115), .Y(n114) );
  AOI21X1 U217 ( .A0(n138), .A1(n139), .B0(n34), .Y(n137) );
  NAND2BX1 U218 ( .AN(n140), .B(n141), .Y(n138) );
  AND2X2 U219 ( .A(n91), .B(n94), .Y(n32) );
  INVX1 U220 ( .A(n110), .Y(n119) );
  NAND2X1 U221 ( .A(n91), .B(n92), .Y(n90) );
  NAND2X1 U222 ( .A(n116), .B(n117), .Y(n113) );
  NAND2X1 U223 ( .A(n112), .B(n118), .Y(n116) );
  OAI21XL U224 ( .A0(n119), .A1(n120), .B0(n121), .Y(n118) );
  NAND2XL U225 ( .A(B[7]), .B(A[7]), .Y(n50) );
  NAND2XL U226 ( .A(B[9]), .B(A[9]), .Y(n38) );
  NAND2XL U227 ( .A(B[10]), .B(A[10]), .Y(n245) );
  NAND2XL U228 ( .A(B[15]), .B(A[15]), .Y(n202) );
  NAND2XL U229 ( .A(B[11]), .B(A[11]), .Y(n247) );
  XOR3X2 U230 ( .A(B[31]), .B(A[31]), .C(n90), .Y(SUM[31]) );
  OR2X2 U231 ( .A(A[22]), .B(B[22]), .Y(n146) );
  NOR2X1 U232 ( .A(A[23]), .B(B[23]), .Y(n34) );
  OR2X2 U233 ( .A(A[24]), .B(B[24]), .Y(n130) );
  OR2X2 U234 ( .A(A[26]), .B(B[26]), .Y(n112) );
  NAND2X1 U235 ( .A(B[26]), .B(A[26]), .Y(n117) );
  OR2X2 U236 ( .A(A[27]), .B(B[27]), .Y(n111) );
  NAND2X1 U237 ( .A(B[27]), .B(A[27]), .Y(n115) );
  NAND2X1 U238 ( .A(B[28]), .B(A[28]), .Y(n106) );
  OR2X2 U239 ( .A(A[28]), .B(B[28]), .Y(n104) );
  NAND2X1 U240 ( .A(B[30]), .B(A[30]), .Y(n91) );
  NAND2X1 U241 ( .A(B[29]), .B(A[29]), .Y(n97) );
  OR2X2 U242 ( .A(A[30]), .B(B[30]), .Y(n94) );
  OR2X2 U243 ( .A(A[29]), .B(B[29]), .Y(n98) );
  NAND3BX4 U244 ( .AN(n195), .B(n268), .C(n74), .Y(n56) );
  NAND3X4 U245 ( .A(n187), .B(n188), .C(n186), .Y(n182) );
  NAND2X2 U246 ( .A(B[2]), .B(A[2]), .Y(n84) );
  INVX8 U247 ( .A(n58), .Y(n69) );
  OAI21X2 U248 ( .A0(n78), .A1(n40), .B0(n41), .Y(n36) );
  NAND2X2 U249 ( .A(B[3]), .B(A[3]), .Y(n74) );
  NAND2X4 U250 ( .A(n270), .B(n196), .Y(n268) );
  XOR2X4 U251 ( .A(n47), .B(n48), .Y(SUM[8]) );
  OAI2BB1X4 U252 ( .A0N(B[0]), .A1N(A[0]), .B0(n89), .Y(n196) );
  OAI21X2 U253 ( .A0(n71), .A1(n72), .B0(n73), .Y(n67) );
  XOR2X4 U254 ( .A(n36), .B(n37), .Y(SUM[9]) );
  XOR2X4 U255 ( .A(n64), .B(n25), .Y(SUM[6]) );
  XOR2X4 U256 ( .A(n79), .B(n80), .Y(SUM[3]) );
  NAND2X4 U257 ( .A(n152), .B(n144), .Y(n150) );
  NAND2X4 U258 ( .A(n147), .B(n153), .Y(n152) );
  NOR2BX4 U259 ( .AN(n89), .B(n174), .Y(n173) );
  XOR2X4 U260 ( .A(n175), .B(n176), .Y(SUM[19]) );
  OAI21X4 U261 ( .A0(n177), .A1(n165), .B0(n164), .Y(n175) );
  NAND2X4 U262 ( .A(n159), .B(n168), .Y(n180) );
  NAND2X4 U263 ( .A(n182), .B(n183), .Y(n159) );
  NAND2X4 U264 ( .A(n211), .B(n212), .Y(n186) );
  CLKINVX3 U265 ( .A(n213), .Y(n211) );
  NOR2X4 U266 ( .A(n201), .B(n217), .Y(n216) );
  CLKINVX3 U267 ( .A(n218), .Y(n201) );
  NOR2X4 U268 ( .A(n207), .B(n219), .Y(n215) );
  XOR2X4 U269 ( .A(n221), .B(n220), .Y(SUM[15]) );
  CLKINVX3 U270 ( .A(n203), .Y(n217) );
  OR2X4 U271 ( .A(A[15]), .B(B[15]), .Y(n218) );
  XOR2X4 U272 ( .A(n225), .B(n226), .Y(SUM[14]) );
  OR2X4 U273 ( .A(A[14]), .B(B[14]), .Y(n203) );
  CLKINVX3 U274 ( .A(n227), .Y(n207) );
  OR2X4 U275 ( .A(A[13]), .B(B[13]), .Y(n227) );
  OAI21X4 U276 ( .A0(n230), .A1(n231), .B0(n232), .Y(n223) );
  CLKINVX3 U277 ( .A(n237), .Y(n219) );
  OR2X4 U278 ( .A(A[12]), .B(B[12]), .Y(n237) );
  NAND2BX4 U279 ( .AN(n241), .B(n238), .Y(n213) );
  OAI2BB1X4 U280 ( .A0N(n242), .A1N(n243), .B0(n244), .Y(n238) );
  NAND2X4 U281 ( .A(n249), .B(n250), .Y(n193) );
  NOR2X4 U282 ( .A(n45), .B(n39), .Y(n250) );
  CLKINVX3 U283 ( .A(n42), .Y(n45) );
  NOR2X4 U284 ( .A(n248), .B(n241), .Y(n249) );
  CLKINVX3 U285 ( .A(n236), .Y(n241) );
  OAI21X4 U286 ( .A0(n78), .A1(n191), .B0(n252), .Y(n47) );
  XOR2X4 U287 ( .A(n253), .B(n24), .Y(SUM[11]) );
  OR2X4 U288 ( .A(A[11]), .B(B[11]), .Y(n236) );
  NAND2BX4 U289 ( .AN(n254), .B(n255), .Y(n253) );
  XOR2X4 U290 ( .A(n261), .B(n262), .Y(SUM[10]) );
  CLKINVX3 U291 ( .A(n258), .Y(n248) );
  OR2X4 U292 ( .A(A[10]), .B(B[10]), .Y(n258) );
  OR2X4 U293 ( .A(A[8]), .B(B[8]), .Y(n42) );
  NAND2X4 U294 ( .A(B[4]), .B(A[4]), .Y(n57) );
  NAND3X4 U295 ( .A(n85), .B(n269), .C(n86), .Y(n72) );
  OR2X4 U296 ( .A(B[1]), .B(A[1]), .Y(n86) );
  OR2X4 U297 ( .A(A[2]), .B(B[2]), .Y(n85) );
  NAND2BX4 U298 ( .AN(n84), .B(n269), .Y(n73) );
  OR2X4 U299 ( .A(A[3]), .B(B[3]), .Y(n269) );
  NAND2X4 U300 ( .A(n271), .B(n272), .Y(n191) );
  OR2X4 U301 ( .A(A[6]), .B(B[6]), .Y(n59) );
  CLKINVX3 U302 ( .A(n55), .Y(n70) );
  OR2X4 U303 ( .A(A[4]), .B(B[4]), .Y(n55) );
  OR2X4 U304 ( .A(A[5]), .B(B[5]), .Y(n58) );
endmodule


module hash_core_DW01_add_38 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n278, n279, n280, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277;

  NOR2X4 U2 ( .A(n85), .B(n276), .Y(n273) );
  NOR2X1 U3 ( .A(n123), .B(n124), .Y(n122) );
  NAND2X2 U4 ( .A(n116), .B(n117), .Y(n114) );
  NAND3BX2 U5 ( .AN(n61), .B(n78), .C(B[5]), .Y(n277) );
  NOR3BX2 U6 ( .AN(n211), .B(n216), .C(n220), .Y(n219) );
  AND2X4 U7 ( .A(n79), .B(n56), .Y(n24) );
  INVX8 U8 ( .A(n170), .Y(n149) );
  NAND2X1 U9 ( .A(B[19]), .B(A[19]), .Y(n184) );
  AOI21X4 U10 ( .A0(n211), .A1(n206), .B0(n245), .Y(n244) );
  NAND2X4 U11 ( .A(n1), .B(n204), .Y(n261) );
  AND2X2 U12 ( .A(n70), .B(n215), .Y(n1) );
  OR2X4 U13 ( .A(A[1]), .B(B[1]), .Y(n111) );
  INVX8 U14 ( .A(n220), .Y(n265) );
  DLY1X1 U15 ( .A(n204), .Y(n18) );
  BUFX12 U16 ( .A(n278), .Y(SUM[26]) );
  CLKINVX3 U17 ( .A(n279), .Y(n2) );
  INVX4 U18 ( .A(n2), .Y(SUM[20]) );
  XOR2X2 U19 ( .A(n116), .B(n118), .Y(SUM[28]) );
  BUFX3 U20 ( .A(n164), .Y(n4) );
  NAND2BX4 U21 ( .AN(n258), .B(n259), .Y(n257) );
  AOI21X4 U22 ( .A0(n112), .A1(n187), .B0(n186), .Y(n267) );
  NAND2X2 U23 ( .A(n79), .B(n274), .Y(n87) );
  NOR2BX4 U24 ( .AN(n211), .B(n216), .Y(n242) );
  AOI21X4 U25 ( .A0(n273), .A1(n52), .B0(n275), .Y(n272) );
  CLKINVX4 U26 ( .A(B[12]), .Y(n13) );
  OAI21X2 U27 ( .A0(n120), .A1(n121), .B0(n122), .Y(n116) );
  NOR4X2 U28 ( .A(n50), .B(n49), .C(n176), .D(n177), .Y(n175) );
  OAI21X1 U29 ( .A0(n176), .A1(n182), .B0(n183), .Y(n181) );
  INVX2 U30 ( .A(n195), .Y(n176) );
  NAND2X2 U31 ( .A(n174), .B(n175), .Y(n173) );
  XOR2X2 U32 ( .A(n144), .B(n146), .Y(SUM[24]) );
  INVX4 U33 ( .A(n110), .Y(n30) );
  NOR2BX4 U34 ( .AN(n98), .B(n53), .Y(n110) );
  BUFX8 U35 ( .A(n82), .Y(n57) );
  NAND2X2 U36 ( .A(n82), .B(n276), .Y(n81) );
  NAND2X2 U37 ( .A(B[5]), .B(A[5]), .Y(n82) );
  NOR2X4 U38 ( .A(A[19]), .B(B[19]), .Y(n50) );
  NOR2BX2 U39 ( .AN(n112), .B(n186), .Y(n185) );
  CLKINVX4 U40 ( .A(n276), .Y(n88) );
  NOR2BX4 U41 ( .AN(n276), .B(n93), .Y(n92) );
  OAI2BB1X4 U42 ( .A0N(n79), .A1N(n56), .B0(n276), .Y(n89) );
  NAND2X4 U43 ( .A(B[4]), .B(A[4]), .Y(n276) );
  NAND2X2 U44 ( .A(B[6]), .B(A[6]), .Y(n76) );
  INVX4 U45 ( .A(n111), .Y(n186) );
  NAND2X2 U46 ( .A(B[17]), .B(A[17]), .Y(n183) );
  OR2X4 U47 ( .A(A[17]), .B(B[17]), .Y(n195) );
  NAND2X4 U48 ( .A(n31), .B(n32), .Y(SUM[2]) );
  XOR2X2 U49 ( .A(n36), .B(n185), .Y(SUM[1]) );
  OAI21X2 U50 ( .A0(n29), .A1(n53), .B0(n98), .Y(n94) );
  NOR2BXL U51 ( .AN(n132), .B(n130), .Y(n143) );
  INVX1 U52 ( .A(n206), .Y(n12) );
  NAND2X1 U53 ( .A(B[14]), .B(A[14]), .Y(n229) );
  CLKINVX2 U54 ( .A(n15), .Y(n256) );
  INVX4 U55 ( .A(n240), .Y(n238) );
  NAND2XL U56 ( .A(B[27]), .B(A[27]), .Y(n133) );
  INVX2 U57 ( .A(n167), .Y(n43) );
  NOR2BXL U58 ( .AN(n76), .B(n85), .Y(n84) );
  INVX1 U59 ( .A(n76), .Y(n275) );
  INVX1 U60 ( .A(n209), .Y(n223) );
  NOR2X2 U61 ( .A(B[7]), .B(A[7]), .Y(n270) );
  INVX1 U62 ( .A(n246), .Y(n245) );
  NOR2X2 U63 ( .A(n213), .B(n212), .Y(n203) );
  NAND2X2 U64 ( .A(n10), .B(n230), .Y(n225) );
  NAND2X1 U65 ( .A(n40), .B(n27), .Y(n28) );
  OR2X2 U66 ( .A(A[23]), .B(B[23]), .Y(n162) );
  NAND2X1 U67 ( .A(B[16]), .B(A[16]), .Y(n182) );
  INVX1 U68 ( .A(n65), .Y(n264) );
  AOI21X2 U69 ( .A0(n65), .A1(n69), .B0(n15), .Y(n249) );
  OR2X2 U70 ( .A(A[16]), .B(B[16]), .Y(n196) );
  NOR2X2 U71 ( .A(A[21]), .B(B[21]), .Y(n48) );
  INVX4 U72 ( .A(n78), .Y(n85) );
  INVX1 U73 ( .A(n133), .Y(n123) );
  NAND2X1 U74 ( .A(B[24]), .B(A[24]), .Y(n131) );
  OAI2BB1X2 U75 ( .A0N(n111), .A1N(n36), .B0(n112), .Y(n99) );
  NAND2BX2 U76 ( .AN(n60), .B(A[3]), .Y(n96) );
  NAND2X2 U77 ( .A(B[1]), .B(A[1]), .Y(n112) );
  AND2X2 U78 ( .A(B[0]), .B(A[0]), .Y(n36) );
  NOR2BX2 U79 ( .AN(n235), .B(n237), .Y(n236) );
  NOR2BX1 U80 ( .AN(n180), .B(n49), .Y(n192) );
  INVX1 U81 ( .A(n141), .Y(n130) );
  NAND2X1 U82 ( .A(n29), .B(n110), .Y(n32) );
  NAND2X1 U83 ( .A(n99), .B(n30), .Y(n31) );
  XOR2X2 U84 ( .A(n103), .B(n105), .Y(SUM[30]) );
  OAI21X2 U85 ( .A0(n138), .A1(n128), .B0(n126), .Y(n136) );
  NOR2X1 U86 ( .A(n48), .B(n51), .Y(n160) );
  AND2X2 U87 ( .A(n227), .B(n209), .Y(n5) );
  AND2X2 U88 ( .A(n195), .B(n196), .Y(n6) );
  AND2X2 U89 ( .A(A[12]), .B(n14), .Y(n7) );
  AND2X2 U90 ( .A(n253), .B(n254), .Y(n8) );
  AND2X2 U91 ( .A(n70), .B(n56), .Y(n9) );
  CLKINVX3 U92 ( .A(n99), .Y(n29) );
  AND2X2 U93 ( .A(n33), .B(n229), .Y(n10) );
  AND2X2 U94 ( .A(n28), .B(n158), .Y(n11) );
  NOR3X4 U95 ( .A(n12), .B(n207), .C(n208), .Y(n205) );
  INVX1 U96 ( .A(n227), .Y(n226) );
  CLKINVX3 U97 ( .A(n13), .Y(n14) );
  AND2X1 U98 ( .A(n246), .B(n211), .Y(n45) );
  INVX3 U99 ( .A(n232), .Y(n21) );
  OAI21X4 U100 ( .A0(n165), .A1(n156), .B0(n154), .Y(n163) );
  INVX3 U101 ( .A(n166), .Y(n165) );
  NOR2X4 U102 ( .A(n247), .B(n206), .Y(n38) );
  OAI2BB1X2 U103 ( .A0N(A[7]), .A1N(B[7]), .B0(n277), .Y(n271) );
  INVXL U104 ( .A(B[7]), .Y(n58) );
  OR2X4 U105 ( .A(A[5]), .B(B[5]), .Y(n52) );
  OR2X2 U106 ( .A(A[5]), .B(B[5]), .Y(n274) );
  NOR2X4 U107 ( .A(A[9]), .B(B[9]), .Y(n15) );
  INVX1 U108 ( .A(n214), .Y(n237) );
  NOR2X4 U109 ( .A(A[11]), .B(B[11]), .Y(n17) );
  AOI21X4 U110 ( .A0(n67), .A1(n35), .B0(n216), .Y(n247) );
  NAND2BX4 U111 ( .AN(n73), .B(n204), .Y(n67) );
  INVX4 U112 ( .A(n191), .Y(n190) );
  NAND2X2 U113 ( .A(B[11]), .B(A[11]), .Y(n253) );
  NOR2X2 U114 ( .A(n16), .B(n17), .Y(n248) );
  INVX3 U115 ( .A(n253), .Y(n252) );
  AOI21X4 U116 ( .A0(n196), .A1(n174), .B0(n198), .Y(n197) );
  OAI2BB1X2 U117 ( .A0N(n215), .A1N(n204), .B0(n35), .Y(n243) );
  NOR2X2 U118 ( .A(n88), .B(n56), .Y(n86) );
  OAI21X4 U119 ( .A0(n86), .A1(n87), .B0(n57), .Y(n83) );
  NOR2X2 U120 ( .A(B[10]), .B(A[10]), .Y(n16) );
  NAND2X1 U121 ( .A(B[25]), .B(A[25]), .Y(n132) );
  NOR2BX2 U122 ( .AN(n187), .B(n39), .Y(SUM[0]) );
  NAND3X4 U123 ( .A(n201), .B(n202), .C(n200), .Y(n19) );
  NAND3X4 U124 ( .A(n217), .B(n218), .C(n219), .Y(n201) );
  OAI21X4 U125 ( .A0(n238), .A1(n239), .B0(n33), .Y(n20) );
  NOR2BX1 U126 ( .AN(n65), .B(n15), .Y(n64) );
  NAND2X2 U127 ( .A(n14), .B(A[12]), .Y(n246) );
  NAND3X1 U128 ( .A(n160), .B(n161), .C(n162), .Y(n148) );
  INVX2 U129 ( .A(n161), .Y(n156) );
  XOR2X2 U130 ( .A(n142), .B(n143), .Y(SUM[25]) );
  NAND2X2 U131 ( .A(n7), .B(n210), .Y(n230) );
  NAND2X2 U132 ( .A(n209), .B(n210), .Y(n208) );
  NAND2BX4 U133 ( .AN(n5), .B(n21), .Y(n22) );
  OR2X4 U134 ( .A(A[5]), .B(B[5]), .Y(n77) );
  INVX4 U135 ( .A(n210), .Y(n239) );
  NOR2X4 U136 ( .A(n97), .B(n53), .Y(n268) );
  INVX8 U137 ( .A(n269), .Y(n97) );
  CLKINVX8 U138 ( .A(n25), .Y(n26) );
  NAND2X2 U139 ( .A(B[10]), .B(A[10]), .Y(n251) );
  AOI21X4 U140 ( .A0(n203), .A1(n18), .B0(n205), .Y(n202) );
  INVX4 U141 ( .A(n139), .Y(n138) );
  NAND2X2 U142 ( .A(n265), .B(n56), .Y(n68) );
  OR2X4 U143 ( .A(A[27]), .B(B[27]), .Y(n135) );
  NAND2X2 U144 ( .A(n232), .B(n5), .Y(n23) );
  NAND2X4 U145 ( .A(n22), .B(n23), .Y(SUM[15]) );
  NOR2X4 U146 ( .A(n24), .B(n81), .Y(n74) );
  OAI21X4 U147 ( .A0(n74), .A1(n75), .B0(n76), .Y(n71) );
  NAND2X4 U148 ( .A(n69), .B(n261), .Y(n25) );
  NAND2X4 U149 ( .A(n26), .B(n262), .Y(n63) );
  NAND2X4 U150 ( .A(n9), .B(n265), .Y(n262) );
  CLKINVX3 U151 ( .A(n157), .Y(n27) );
  NAND2X4 U152 ( .A(n19), .B(n6), .Y(n194) );
  XOR2X4 U153 ( .A(n109), .B(n113), .Y(SUM[29]) );
  NAND2X4 U154 ( .A(n114), .B(n115), .Y(n109) );
  OAI21X4 U155 ( .A0(n51), .A1(n149), .B0(n157), .Y(n168) );
  INVX2 U156 ( .A(n79), .Y(n93) );
  CLKBUFX8 U157 ( .A(n228), .Y(n33) );
  NAND4BX4 U158 ( .AN(n270), .B(n77), .C(n78), .D(n79), .Y(n220) );
  OAI21X4 U159 ( .A0(n54), .A1(n107), .B0(n108), .Y(n103) );
  NAND3X1 U160 ( .A(n69), .B(n261), .C(n262), .Y(n260) );
  AOI21X4 U161 ( .A0(n214), .A1(n20), .B0(n234), .Y(n232) );
  XOR2X2 U162 ( .A(n168), .B(n169), .Y(SUM[21]) );
  OAI21X2 U163 ( .A0(n130), .A1(n131), .B0(n132), .Y(n129) );
  XOR2X4 U164 ( .A(n139), .B(n140), .Y(n278) );
  XOR2X2 U165 ( .A(n56), .B(n92), .Y(SUM[4]) );
  XOR2X4 U166 ( .A(n89), .B(n90), .Y(SUM[5]) );
  NOR2BX2 U167 ( .AN(n154), .B(n156), .Y(n167) );
  NAND2X2 U168 ( .A(B[0]), .B(A[0]), .Y(n187) );
  NOR2X1 U169 ( .A(A[0]), .B(B[0]), .Y(n39) );
  BUFX8 U170 ( .A(n68), .Y(n35) );
  NAND2X1 U171 ( .A(B[21]), .B(A[21]), .Y(n158) );
  OR2XL U172 ( .A(A[24]), .B(B[24]), .Y(n145) );
  OAI21X1 U173 ( .A0(B[14]), .A1(A[14]), .B0(n211), .Y(n207) );
  NAND2XL U174 ( .A(B[13]), .B(A[13]), .Y(n228) );
  XNOR2X4 U175 ( .A(n83), .B(n62), .Y(SUM[6]) );
  INVX2 U176 ( .A(n162), .Y(n155) );
  NOR2BXL U177 ( .AN(n159), .B(n155), .Y(n164) );
  NAND2X1 U178 ( .A(B[18]), .B(A[18]), .Y(n180) );
  XNOR2X4 U179 ( .A(n166), .B(n43), .Y(SUM[22]) );
  NOR2BX4 U180 ( .AN(n33), .B(n239), .Y(n241) );
  NOR2BXL U181 ( .AN(n133), .B(n127), .Y(n137) );
  NOR2BX1 U182 ( .AN(n184), .B(n50), .Y(n189) );
  NAND2X2 U183 ( .A(B[8]), .B(A[8]), .Y(n69) );
  NOR2X4 U184 ( .A(A[18]), .B(B[18]), .Y(n49) );
  NOR2X2 U185 ( .A(n151), .B(n152), .Y(n150) );
  INVX4 U186 ( .A(n95), .Y(n37) );
  NOR2BX1 U187 ( .AN(n157), .B(n51), .Y(n171) );
  XOR2X4 U188 ( .A(n191), .B(n192), .Y(SUM[18]) );
  AOI21X2 U189 ( .A0(n179), .A1(n180), .B0(n50), .Y(n178) );
  INVX1 U190 ( .A(n135), .Y(n127) );
  NOR2X4 U191 ( .A(B[2]), .B(A[2]), .Y(n53) );
  XNOR2X4 U192 ( .A(n94), .B(n37), .Y(SUM[3]) );
  NOR2BX4 U193 ( .AN(n57), .B(n91), .Y(n90) );
  INVX4 U194 ( .A(n77), .Y(n91) );
  BUFX12 U195 ( .A(n80), .Y(n56) );
  INVX4 U196 ( .A(n221), .Y(n266) );
  INVX4 U197 ( .A(n134), .Y(n128) );
  INVXL U198 ( .A(n117), .Y(n119) );
  NOR2BXL U199 ( .AN(n126), .B(n128), .Y(n140) );
  OR2X4 U200 ( .A(n156), .B(n11), .Y(n153) );
  NAND2XL U201 ( .A(n103), .B(n104), .Y(n102) );
  INVX4 U202 ( .A(n41), .Y(SUM[17]) );
  XNOR2X4 U203 ( .A(n45), .B(n38), .Y(SUM[12]) );
  INVX1 U204 ( .A(n48), .Y(n40) );
  NOR2BX2 U205 ( .AN(n184), .B(n178), .Y(n172) );
  NOR2XL U206 ( .A(n182), .B(n176), .Y(n193) );
  NOR2BXL U207 ( .AN(n182), .B(n177), .Y(n199) );
  OR2X4 U208 ( .A(A[4]), .B(B[4]), .Y(n79) );
  OR2X4 U209 ( .A(A[22]), .B(B[22]), .Y(n161) );
  NAND2XL U210 ( .A(B[22]), .B(A[22]), .Y(n154) );
  OR2X4 U211 ( .A(A[13]), .B(B[13]), .Y(n210) );
  NAND2X2 U212 ( .A(B[20]), .B(A[20]), .Y(n157) );
  NAND2XL U213 ( .A(B[30]), .B(A[30]), .Y(n101) );
  NAND2XL U214 ( .A(B[28]), .B(A[28]), .Y(n115) );
  NAND2XL U215 ( .A(B[23]), .B(A[23]), .Y(n159) );
  INVXL U216 ( .A(A[7]), .Y(n59) );
  INVXL U217 ( .A(A[5]), .Y(n61) );
  INVX1 U218 ( .A(n84), .Y(n62) );
  INVX1 U219 ( .A(n109), .Y(n107) );
  NAND3BX1 U220 ( .AN(n130), .B(n134), .C(n135), .Y(n121) );
  OAI2BB1X4 U221 ( .A0N(n168), .A1N(n40), .B0(n158), .Y(n166) );
  XOR2X2 U222 ( .A(n42), .B(n197), .Y(n41) );
  AND2X1 U223 ( .A(n183), .B(n195), .Y(n42) );
  INVX1 U224 ( .A(n235), .Y(n234) );
  OAI21XL U225 ( .A0(n16), .A1(n65), .B0(n251), .Y(n258) );
  INVX1 U226 ( .A(n196), .Y(n177) );
  NAND2BX1 U227 ( .AN(n49), .B(n181), .Y(n179) );
  XOR2X4 U228 ( .A(n44), .B(n66), .Y(SUM[8]) );
  AND2X1 U229 ( .A(n69), .B(n70), .Y(n44) );
  NOR2BX1 U230 ( .AN(n131), .B(n147), .Y(n146) );
  INVX1 U231 ( .A(n145), .Y(n147) );
  NOR2BX1 U232 ( .AN(n101), .B(n106), .Y(n105) );
  INVX1 U233 ( .A(n104), .Y(n106) );
  NOR2BX1 U234 ( .AN(n115), .B(n119), .Y(n118) );
  NOR2BX1 U235 ( .AN(n158), .B(n48), .Y(n169) );
  XOR2X1 U236 ( .A(n170), .B(n171), .Y(n279) );
  NOR2BX1 U237 ( .AN(n108), .B(n54), .Y(n113) );
  AOI21X1 U238 ( .A0(n125), .A1(n126), .B0(n127), .Y(n124) );
  NAND2BX1 U239 ( .AN(n128), .B(n129), .Y(n125) );
  AOI21X2 U240 ( .A0(n153), .A1(n154), .B0(n155), .Y(n152) );
  XNOR2X4 U241 ( .A(n263), .B(n46), .Y(SUM[10]) );
  AND2X1 U242 ( .A(n251), .B(n255), .Y(n46) );
  NOR2BX2 U243 ( .AN(n209), .B(n231), .Y(n224) );
  NOR2X2 U244 ( .A(n231), .B(n239), .Y(n218) );
  NAND2X2 U245 ( .A(n47), .B(n260), .Y(n259) );
  AND2X1 U246 ( .A(n255), .B(n256), .Y(n47) );
  INVX1 U247 ( .A(n159), .Y(n151) );
  INVX1 U248 ( .A(n182), .Y(n198) );
  NOR2X1 U249 ( .A(A[20]), .B(B[20]), .Y(n51) );
  NAND2X2 U250 ( .A(B[9]), .B(A[9]), .Y(n65) );
  NAND2XL U251 ( .A(B[15]), .B(A[15]), .Y(n227) );
  NAND2XL U252 ( .A(B[14]), .B(A[14]), .Y(n235) );
  OR2X2 U253 ( .A(A[26]), .B(B[26]), .Y(n134) );
  OR2X2 U254 ( .A(A[25]), .B(B[25]), .Y(n141) );
  NAND2X1 U255 ( .A(B[26]), .B(A[26]), .Y(n126) );
  NOR2X1 U256 ( .A(A[29]), .B(B[29]), .Y(n54) );
  NAND2X1 U257 ( .A(B[29]), .B(A[29]), .Y(n108) );
  OR2X2 U258 ( .A(A[28]), .B(B[28]), .Y(n117) );
  OR2X2 U259 ( .A(A[30]), .B(B[30]), .Y(n104) );
  XOR3X2 U260 ( .A(B[31]), .B(A[31]), .C(n100), .Y(SUM[31]) );
  NAND2X1 U261 ( .A(n101), .B(n102), .Y(n100) );
  NAND3BX4 U262 ( .AN(n266), .B(n96), .C(n222), .Y(n80) );
  NAND3X4 U263 ( .A(n201), .B(n202), .C(n200), .Y(n174) );
  NOR2X2 U264 ( .A(B[14]), .B(A[14]), .Y(n231) );
  NAND2X1 U265 ( .A(n274), .B(n78), .Y(n75) );
  BUFX4 U266 ( .A(n280), .Y(SUM[16]) );
  AOI2BB1X4 U267 ( .A0N(n58), .A1N(n59), .B0(n73), .Y(n72) );
  NAND3BX2 U268 ( .AN(n216), .B(n210), .C(n211), .Y(n212) );
  INVXL U269 ( .A(B[3]), .Y(n60) );
  XOR2X1 U270 ( .A(n19), .B(n199), .Y(n280) );
  XOR2X4 U271 ( .A(n63), .B(n64), .Y(SUM[9]) );
  NAND2X4 U272 ( .A(n67), .B(n35), .Y(n66) );
  XOR2X4 U273 ( .A(n71), .B(n72), .Y(SUM[7]) );
  NOR2BX4 U274 ( .AN(n96), .B(n97), .Y(n95) );
  XOR2X4 U275 ( .A(n136), .B(n137), .Y(SUM[27]) );
  OAI2BB1X4 U276 ( .A0N(n141), .A1N(n142), .B0(n132), .Y(n139) );
  NAND2X4 U277 ( .A(n120), .B(n131), .Y(n142) );
  NAND2X4 U278 ( .A(n144), .B(n145), .Y(n120) );
  OAI21X4 U279 ( .A0(n148), .A1(n149), .B0(n150), .Y(n144) );
  XOR2X4 U280 ( .A(n163), .B(n4), .Y(SUM[23]) );
  NAND2X4 U281 ( .A(n172), .B(n173), .Y(n170) );
  XOR2X4 U282 ( .A(n188), .B(n189), .Y(SUM[19]) );
  OAI21X4 U283 ( .A0(n190), .A1(n49), .B0(n180), .Y(n188) );
  NAND3BX4 U284 ( .AN(n193), .B(n183), .C(n194), .Y(n191) );
  NAND3X4 U285 ( .A(n209), .B(n214), .C(n215), .Y(n213) );
  AOI31X2 U286 ( .A0(n96), .A1(n221), .A2(n222), .B0(n223), .Y(n217) );
  AOI21X4 U287 ( .A0(n224), .A1(n225), .B0(n226), .Y(n200) );
  OR2X4 U288 ( .A(A[15]), .B(B[15]), .Y(n209) );
  XOR2X4 U289 ( .A(n233), .B(n236), .Y(SUM[14]) );
  OR2X4 U290 ( .A(B[14]), .B(A[14]), .Y(n214) );
  OAI21X4 U291 ( .A0(n238), .A1(n239), .B0(n33), .Y(n233) );
  XOR2X4 U292 ( .A(n240), .B(n241), .Y(SUM[13]) );
  OAI2BB1X4 U293 ( .A0N(n242), .A1N(n243), .B0(n244), .Y(n240) );
  OAI2BB1X4 U294 ( .A0N(n248), .A1N(n249), .B0(n250), .Y(n206) );
  AOI2BB1X4 U295 ( .A0N(n17), .A1N(n251), .B0(n252), .Y(n250) );
  NAND4BX4 U296 ( .AN(n15), .B(n70), .C(n254), .D(n255), .Y(n216) );
  CLKINVX3 U297 ( .A(n215), .Y(n73) );
  OR2X4 U298 ( .A(A[12]), .B(B[12]), .Y(n211) );
  XOR2X4 U299 ( .A(n257), .B(n8), .Y(SUM[11]) );
  OR2X4 U300 ( .A(B[11]), .B(A[11]), .Y(n254) );
  AOI21X4 U301 ( .A0(n256), .A1(n63), .B0(n264), .Y(n263) );
  NAND2X4 U302 ( .A(n267), .B(n268), .Y(n222) );
  NAND2BX4 U303 ( .AN(n98), .B(n269), .Y(n221) );
  OR2X4 U304 ( .A(A[3]), .B(B[3]), .Y(n269) );
  NAND2X4 U305 ( .A(B[2]), .B(A[2]), .Y(n98) );
  NAND2BX4 U306 ( .AN(n271), .B(n272), .Y(n204) );
  OR2X4 U307 ( .A(A[6]), .B(B[6]), .Y(n78) );
  OR2X4 U308 ( .A(A[7]), .B(B[7]), .Y(n215) );
  OR2X4 U309 ( .A(B[8]), .B(A[8]), .Y(n70) );
  OR2X4 U310 ( .A(B[10]), .B(A[10]), .Y(n255) );
endmodule


module hash_core ( clk, reset, Wt, inner_busy, first_block, output_enable, 
        digest );
  input [31:0] Wt;
  output [7:0] digest;
  input clk, reset, inner_busy, first_block, output_enable;
  wire   N145, N146, N147, N148, N149, N150, N151, N819, N820, N821, N822,
         N823, N824, N825, N826, N827, N828, N829, N830, N831, N832, N833,
         N834, N835, N836, N837, N838, N839, N840, N841, N842, N843, N844,
         N845, N846, N847, N848, N849, N850, N851, N852, N853, N854, N855,
         N856, N857, N858, N859, N860, N861, N862, N863, N864, N865, N866,
         N867, N868, N869, N870, N871, N872, N873, N874, N875, N876, N877,
         N878, N879, N880, N881, N882, N883, N884, N885, N886, N887, N888,
         N889, N890, N891, N892, N893, N894, N895, N896, N897, N898, N899,
         N900, N901, N902, N903, N904, N905, N906, N907, N908, N909, N910,
         N911, N912, N913, N914, N915, N916, N917, N918, N919, N920, N921,
         N922, N923, N924, N925, N926, N927, N928, N929, N930, N931, N932,
         N933, N934, N935, N936, N937, N938, N939, N940, N941, N942, N943,
         N944, N945, N946, N947, N948, N949, N950, N951, N952, N953, N954,
         N955, N956, N957, N958, N959, N960, N961, N962, N963, N964, N965,
         N966, N967, N968, N969, N970, N971, N972, N973, N974, N975, N976,
         N977, N978, N979, N980, N981, N982, N983, N984, N985, N986, N987,
         N988, N989, N990, N991, N992, N993, N994, N995, N996, N997, N998,
         N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008,
         N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1017, N1018,
         N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028,
         N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036, N1037, N1038,
         N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046, N1047, N1048,
         N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056, N1057, N1058,
         N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066, N1067, N1068,
         N1069, N1070, N1071, N1072, N1073, N1074, N2970, N2971, N2972, N2973,
         N2974, N2975, N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983,
         N2984, N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993,
         N2994, N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3180, N3181,
         N3182, N3183, N3189, N3190, N3191, N3192, N3193, N3194, N3195, N3196,
         N3197, N3198, N3199, N3200, N3201, n1370, n1383, n1388, n1396, n1433,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1455, n1456,
         n1457, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1486, n1487, n1488, n1489,
         n1490, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1610, n1611, n1614, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1630, n1631,
         n1632, n1634, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1719, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1754, n1755, n1756, n1757, n1758, n1759, n1762, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1784, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1848, n1858, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1877, n1974, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2193, n2194, n2195, n2196, n2198, n2199, n2201, n2202, n2203,
         n2204, n2205, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, T2_32_9_, T2_32_8_,
         T2_32_7_, T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_, T2_32_31_,
         T2_32_30_, T2_32_2_, T2_32_29_, T2_32_28_, T2_32_27_, T2_32_26_,
         T2_32_25_, T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_, T2_32_20_,
         T2_32_1_, T2_32_19_, T2_32_18_, T2_32_17_, T2_32_16_, T2_32_15_,
         T2_32_14_, T2_32_13_, T2_32_12_, T2_32_11_, T2_32_10_, T2_32_0_, N99,
         N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85,
         N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71,
         N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57,
         N56, N55, N54, N53, N52, N51, N50, N49, N48, N143, N142, N141, N140,
         N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129,
         N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118,
         N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107,
         N106, N105, N104, N103, N102, N101, N100, n10, n11, n12, n13, n14,
         n15, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985;
  wire   [31:0] f1_EFG_32;
  wire   [31:0] f2_ABC_32;
  wire   [31:0] f3_A_32;
  wire   [31:0] f4_E_32;
  wire   [31:0] Kt;
  wire   [31:0] T1_32;
  wire   [31:0] next_E;
  wire   [31:0] next_A;
  wire   [255:0] SHA256_result;
  wire   [6:2] round;
  wire   [31:0] H0;
  wire   [31:1] H1;
  wire   [31:0] H2;
  wire   [31:1] H3;
  wire   [31:0] H4;
  wire   [31:0] H5;
  wire   [31:0] H6;
  wire   [31:0] H7;
  wire   [4:0] read_counter;

  DFFHQX4 B_reg_0_ ( .D(n2908), .CK(clk), .Q(SHA256_result[192]) );
  DFFHQX4 E_reg_1_ ( .D(n2810), .CK(clk), .Q(SHA256_result[97]) );
  DFFHQX4 E_reg_2_ ( .D(n2809), .CK(clk), .Q(SHA256_result[98]) );
  DFFHQX4 E_reg_4_ ( .D(n2807), .CK(clk), .Q(SHA256_result[100]) );
  DFFHQX4 E_reg_7_ ( .D(n2804), .CK(clk), .Q(SHA256_result[103]) );
  DFFHQX4 E_reg_11_ ( .D(n2800), .CK(clk), .Q(SHA256_result[107]) );
  DFFHQX4 E_reg_13_ ( .D(n2798), .CK(clk), .Q(SHA256_result[109]) );
  DFFHQX4 F_reg_0_ ( .D(n2779), .CK(clk), .Q(SHA256_result[64]) );
  DFFHQX4 F_reg_3_ ( .D(n2776), .CK(clk), .Q(SHA256_result[67]) );
  DFFHQX4 G_reg_2_ ( .D(n2586), .CK(clk), .Q(SHA256_result[34]) );
  DFFHQX4 G_reg_3_ ( .D(n2585), .CK(clk), .Q(SHA256_result[35]) );
  DFFHQX4 Kt_reg_13_ ( .D(N2983), .CK(clk), .Q(Kt[13]) );
  DFFHQX4 Kt_reg_12_ ( .D(N2982), .CK(clk), .Q(Kt[12]) );
  DFFHQX4 Kt_reg_10_ ( .D(N2980), .CK(clk), .Q(Kt[10]) );
  DFFHQX4 Kt_reg_6_ ( .D(N2976), .CK(clk), .Q(Kt[6]) );
  DFFHQX4 Kt_reg_3_ ( .D(N2973), .CK(clk), .Q(Kt[3]) );
  DFFHQX4 Kt_reg_2_ ( .D(N2972), .CK(clk), .Q(Kt[2]) );
  DFFHQX4 Kt_reg_1_ ( .D(N2971), .CK(clk), .Q(Kt[1]) );
  DFFHQX4 Kt_reg_0_ ( .D(N2970), .CK(clk), .Q(Kt[0]) );
  AND2X2 U1356 ( .A(n2164), .B(n2165), .Y(n1987) );
  AND2X2 U1357 ( .A(n2166), .B(n2165), .Y(n1986) );
  AND2X2 U1359 ( .A(n2164), .B(n2167), .Y(n1989) );
  AND2X2 U1360 ( .A(n2166), .B(n2167), .Y(n1988) );
  AND2X2 U1362 ( .A(n2164), .B(n2168), .Y(n1991) );
  AND2X2 U1363 ( .A(n2166), .B(n2168), .Y(n1990) );
  AND2X2 U1365 ( .A(n2164), .B(n2169), .Y(n1993) );
  AND2X2 U1366 ( .A(n2166), .B(n2169), .Y(n1992) );
  AND2X2 U1369 ( .A(n2164), .B(n2174), .Y(n1999) );
  AND2X2 U1370 ( .A(n2166), .B(n2174), .Y(n1998) );
  AND2X2 U1372 ( .A(n2164), .B(n2175), .Y(n2001) );
  AND2X2 U1373 ( .A(n2166), .B(n2175), .Y(n2000) );
  AND2X2 U1375 ( .A(n2164), .B(n2176), .Y(n2003) );
  AND2X2 U1376 ( .A(n2166), .B(n2176), .Y(n2002) );
  AND2X2 U1378 ( .A(n2164), .B(n2177), .Y(n2005) );
  AND2X2 U1379 ( .A(read_counter[4]), .B(read_counter[0]), .Y(n2164) );
  AND2X2 U1380 ( .A(n2166), .B(n2177), .Y(n2004) );
  AND2X2 U1381 ( .A(read_counter[4]), .B(n983), .Y(n2166) );
  AND2X2 U1384 ( .A(n2165), .B(n2182), .Y(n2011) );
  AND2X2 U1385 ( .A(n2165), .B(n2183), .Y(n2010) );
  AND2X2 U1386 ( .A(n2184), .B(n985), .Y(n2165) );
  AND2X2 U1388 ( .A(n2167), .B(n2182), .Y(n2013) );
  AND2X2 U1389 ( .A(n2167), .B(n2183), .Y(n2012) );
  AND2X2 U1390 ( .A(read_counter[3]), .B(n2185), .Y(n2167) );
  AND2X2 U1392 ( .A(n2168), .B(n2182), .Y(n2015) );
  AND2X2 U1393 ( .A(n2168), .B(n2183), .Y(n2014) );
  AND2X2 U1394 ( .A(n2184), .B(read_counter[2]), .Y(n2168) );
  AND2X2 U1395 ( .A(read_counter[3]), .B(n984), .Y(n2184) );
  AND2X2 U1397 ( .A(n2169), .B(n2182), .Y(n2017) );
  AND2X2 U1398 ( .A(n2169), .B(n2183), .Y(n2016) );
  AND2X2 U1402 ( .A(n2182), .B(n2174), .Y(n2022) );
  AND2X2 U1406 ( .A(n2175), .B(n2182), .Y(n2024) );
  AND2X2 U1407 ( .A(n2175), .B(n2183), .Y(n2023) );
  AND2X2 U1411 ( .A(n2176), .B(n2182), .Y(n2026) );
  AND2X2 U1412 ( .A(n2176), .B(n2183), .Y(n2025) );
  AND2X2 U1413 ( .A(n2190), .B(n984), .Y(n2176) );
  AND2X2 U1415 ( .A(n2177), .B(n2182), .Y(n2028) );
  AND2X2 U1417 ( .A(n2177), .B(n2183), .Y(n2027) );
  AND2X2 U1419 ( .A(n2190), .B(read_counter[1]), .Y(n2177) );
  AND2X2 U1481 ( .A(n2309), .B(n367), .Y(n2248) );
  CLKINVX4 U2078 ( .A(reset), .Y(n1433) );
  hash_core_DW01_add_0 add_317 ( .A({SHA256_result[63:46], n12, 
        SHA256_result[44:34], n84, n88}), .B({H7[31:3], n91, n92, H7[0]}), 
        .SUM({N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, 
        N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, 
        N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, 
        N1045, N1044, N1043}) );
  hash_core_DW01_add_1 add_316 ( .A({SHA256_result[95:66], n66, 
        SHA256_result[64]}), .B(H6), .SUM({N1042, N1041, N1040, N1039, N1038, 
        N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, 
        N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, 
        N1017, N1016, N1015, N1014, N1013, N1012, N1011}) );
  hash_core_DW01_add_2 add_315 ( .A({SHA256_result[127], n143, n14, 
        SHA256_result[124:118], n144, SHA256_result[116], n145, 
        SHA256_result[114], n146, SHA256_result[112], n147, 
        SHA256_result[110:109], n148, SHA256_result[107], n149, n150, n151, 
        SHA256_result[103], n152, SHA256_result[101], n43, 
        SHA256_result[99:98], n63, n19}), .B(H5), .SUM({N1010, N1009, N1008, 
        N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, 
        N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, 
        N985, N984, N983, N982, N981, N980, N979}) );
  hash_core_DW01_add_4 add_313 ( .A({SHA256_result[191:163], n94, n121, n71}), 
        .B({H3, n108}), .SUM({N946, N945, N944, N943, N942, N941, N940, N939, 
        N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, 
        N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915}) );
  hash_core_DW01_add_5 add_312 ( .A(SHA256_result[223:192]), .B(H2), .SUM({
        N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, 
        N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, 
        N890, N889, N888, N887, N886, N885, N884, N883}) );
  hash_core_DW01_add_6 add_311 ( .A({SHA256_result[255], n153, n154, n13, n155, 
        n156, n157, n158, n159, SHA256_result[246], n160, n161, n162, n163, 
        n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
        n176, n177, n178, n179, n60, n58}), .B({H1, n90}), .SUM({N882, N881, 
        N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, 
        N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, 
        N856, N855, N854, N853, N852, N851}) );
  hash_core_DW01_inc_0 add_119 ( .A({round[6], n181, n180, round[3:2], n372, 
        n182}), .SUM({N151, N150, N149, N148, N147, N146, N145}) );
  hash_core_DW01_add_15 add_314 ( .A({next_E[31:21], n32, next_E[19:0]}), .B(
        H4), .SUM({N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, 
        N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, 
        N956, N955, N954, N953, N952, N951, N950, N949, N948, N947}) );
  hash_core_DW01_add_16 add_310 ( .A(next_A), .B(H0), .SUM({N850, N849, N848, 
        N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, 
        N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, 
        N823, N822, N821, N820, N819}) );
  hash_core_DW01_add_20 add_1_root_add_0_root_add_113 ( .A(f2_ABC_32), .B(
        f3_A_32), .SUM({T2_32_31_, T2_32_30_, T2_32_29_, T2_32_28_, T2_32_27_, 
        T2_32_26_, T2_32_25_, T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_, 
        T2_32_20_, T2_32_19_, T2_32_18_, T2_32_17_, T2_32_16_, T2_32_15_, 
        T2_32_14_, T2_32_13_, T2_32_12_, T2_32_11_, T2_32_10_, T2_32_9_, 
        T2_32_8_, T2_32_7_, T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_, T2_32_2_, 
        T2_32_1_, T2_32_0_}) );
  hash_core_DW01_add_19 add_0_root_add_0_root_add_108_4 ( .A({N143, N142, N141, 
        N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, 
        N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, 
        N116, N115, N114, N113, N112}), .B({N111, N110, N109, N108, N107, N106, 
        N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, 
        N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80}), 
        .SUM(T1_32) );
  hash_core_DW01_add_26 add_112 ( .A(SHA256_result[159:128]), .B({T1_32[31:14], 
        n10, T1_32[12:8], n31, T1_32[6:0]}), .SUM(next_E) );
  hash_core_DW01_add_27 add_0_root_add_0_root_add_113 ( .A({T2_32_31_, 
        T2_32_30_, T2_32_29_, T2_32_28_, T2_32_27_, T2_32_26_, T2_32_25_, 
        T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_, T2_32_20_, T2_32_19_, 
        T2_32_18_, T2_32_17_, T2_32_16_, T2_32_15_, T2_32_14_, T2_32_13_, 
        T2_32_12_, T2_32_11_, T2_32_10_, T2_32_9_, T2_32_8_, T2_32_7_, 
        T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_, T2_32_2_, T2_32_1_, T2_32_0_}), 
        .B({T1_32[31:14], n10, T1_32[12:8], n31, T1_32[6:0]}), .SUM(next_A) );
  hash_core_DW01_add_30 add_2_root_add_0_root_add_108_4 ( .A(
        SHA256_result[31:0]), .B({f1_EFG_32[31:5], n27, f1_EFG_32[3:0]}), 
        .SUM({N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, 
        N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, 
        N120, N119, N118, N117, N116, N115, N114, N113, N112}) );
  hash_core_DW01_add_32 add_3_root_add_0_root_add_108_4 ( .A(Kt), .B(Wt), 
        .SUM({N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, 
        N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, 
        N52, N51, N50, N49, N48}) );
  hash_core_DW01_add_38 add_1_root_add_0_root_add_108_4 ( .A(f4_E_32), .B({N79, 
        N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, 
        N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, 
        N50, N49, N48}), .SUM({N111, N110, N109, N108, N107, N106, N105, N104, 
        N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, 
        N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80}) );
  DFFHQXL A_reg_30_ ( .D(n2942), .CK(clk), .Q(SHA256_result[254]) );
  DFFHQX1 read_counter_reg_4_ ( .D(N3201), .CK(clk), .Q(read_counter[4]) );
  DFFHQX1 read_counter_reg_0_ ( .D(N3197), .CK(clk), .Q(read_counter[0]) );
  DFFHQX1 read_counter_reg_1_ ( .D(N3198), .CK(clk), .Q(read_counter[1]) );
  DFFHQX1 read_counter_reg_2_ ( .D(N3199), .CK(clk), .Q(read_counter[2]) );
  DFFHQX1 read_counter_reg_3_ ( .D(N3200), .CK(clk), .Q(read_counter[3]) );
  DFFHQX1 Kt_reg_31_ ( .D(N3001), .CK(clk), .Q(Kt[31]) );
  DFFHQX1 Kt_reg_30_ ( .D(N3000), .CK(clk), .Q(Kt[30]) );
  DFFHQX1 Kt_reg_29_ ( .D(N2999), .CK(clk), .Q(Kt[29]) );
  DFFHQX1 Kt_reg_28_ ( .D(N2998), .CK(clk), .Q(Kt[28]) );
  DFFHQX1 Kt_reg_27_ ( .D(N2997), .CK(clk), .Q(Kt[27]) );
  DFFHQX1 Kt_reg_26_ ( .D(N2996), .CK(clk), .Q(Kt[26]) );
  DFFHQX1 Kt_reg_25_ ( .D(N2995), .CK(clk), .Q(Kt[25]) );
  DFFHQX1 Kt_reg_24_ ( .D(N2994), .CK(clk), .Q(Kt[24]) );
  DFFHQX1 Kt_reg_23_ ( .D(N2993), .CK(clk), .Q(Kt[23]) );
  DFFHQX1 H_reg_16_ ( .D(n2540), .CK(clk), .Q(SHA256_result[16]) );
  DFFHQX1 H_reg_18_ ( .D(n2538), .CK(clk), .Q(SHA256_result[18]) );
  DFFHQX1 C_reg_10_ ( .D(n2865), .CK(clk), .Q(SHA256_result[170]) );
  DFFHQX1 C_reg_13_ ( .D(n2862), .CK(clk), .Q(SHA256_result[173]) );
  DFFHQX1 B_reg_12_ ( .D(n2896), .CK(clk), .Q(SHA256_result[204]) );
  DFFHQX1 B_reg_13_ ( .D(n2895), .CK(clk), .Q(SHA256_result[205]) );
  DFFHQX1 B_reg_14_ ( .D(n2894), .CK(clk), .Q(SHA256_result[206]) );
  DFFHQX1 F_reg_20_ ( .D(n2759), .CK(clk), .Q(SHA256_result[84]) );
  DFFHQX1 F_reg_21_ ( .D(n2758), .CK(clk), .Q(SHA256_result[85]) );
  DFFHQX1 G_reg_20_ ( .D(n2568), .CK(clk), .Q(SHA256_result[52]) );
  DFFHQX1 A_reg_6_ ( .D(n2966), .CK(clk), .Q(SHA256_result[230]) );
  DFFHQX1 A_reg_7_ ( .D(n2965), .CK(clk), .Q(SHA256_result[231]) );
  DFFHQX1 A_reg_23_ ( .D(n2949), .CK(clk), .Q(SHA256_result[247]) );
  DFFHQX1 A_reg_24_ ( .D(n2948), .CK(clk), .Q(SHA256_result[248]) );
  DFFHQXL A_reg_25_ ( .D(n2947), .CK(clk), .Q(SHA256_result[249]) );
  DFFHQXL A_reg_26_ ( .D(n2946), .CK(clk), .Q(SHA256_result[250]) );
  DFFHQXL A_reg_27_ ( .D(n2945), .CK(clk), .Q(SHA256_result[251]) );
  DFFHQXL A_reg_29_ ( .D(n2943), .CK(clk), .Q(SHA256_result[253]) );
  DFFHQX1 Kt_reg_22_ ( .D(N2992), .CK(clk), .Q(Kt[22]) );
  DFFHQX1 Kt_reg_21_ ( .D(N2991), .CK(clk), .Q(Kt[21]) );
  DFFHQX1 Kt_reg_20_ ( .D(N2990), .CK(clk), .Q(Kt[20]) );
  DFFHQX1 Kt_reg_19_ ( .D(N2989), .CK(clk), .Q(Kt[19]) );
  DFFHQX1 H6_reg_4_ ( .D(n2615), .CK(clk), .Q(H6[4]) );
  DFFHQX1 F_reg_15_ ( .D(n2764), .CK(clk), .Q(SHA256_result[79]) );
  DFFHQX1 F_reg_16_ ( .D(n2763), .CK(clk), .Q(SHA256_result[80]) );
  DFFHQX1 F_reg_17_ ( .D(n2762), .CK(clk), .Q(SHA256_result[81]) );
  DFFHQX1 G_reg_15_ ( .D(n2573), .CK(clk), .Q(SHA256_result[47]) );
  DFFHQX1 H_reg_15_ ( .D(n2541), .CK(clk), .Q(SHA256_result[15]) );
  DFFHQX1 H_reg_17_ ( .D(n2539), .CK(clk), .Q(SHA256_result[17]) );
  DFFHQX1 C_reg_8_ ( .D(n2867), .CK(clk), .Q(SHA256_result[168]) );
  DFFHQX1 C_reg_5_ ( .D(n2870), .CK(clk), .Q(SHA256_result[165]) );
  DFFHQX1 B_reg_8_ ( .D(n2900), .CK(clk), .Q(SHA256_result[200]) );
  DFFHQX1 B_reg_9_ ( .D(n2899), .CK(clk), .Q(SHA256_result[201]) );
  DFFHQX1 F_reg_18_ ( .D(n2761), .CK(clk), .Q(SHA256_result[82]) );
  DFFHQX1 B_reg_5_ ( .D(n2903), .CK(clk), .Q(SHA256_result[197]) );
  DFFHQX1 A_reg_2_ ( .D(n2970), .CK(clk), .Q(SHA256_result[226]) );
  DFFHQX1 A_reg_3_ ( .D(n2969), .CK(clk), .Q(SHA256_result[227]) );
  DFFHQX1 A_reg_4_ ( .D(n2968), .CK(clk), .Q(SHA256_result[228]) );
  DFFHQX1 A_reg_5_ ( .D(n2967), .CK(clk), .Q(SHA256_result[229]) );
  DFFHQX1 E_reg_19_ ( .D(n2792), .CK(clk), .Q(SHA256_result[115]) );
  DFFHQXL E_reg_30_ ( .D(n2781), .CK(clk), .Q(SHA256_result[126]) );
  DFFHQX1 Kt_reg_18_ ( .D(N2988), .CK(clk), .Q(Kt[18]) );
  DFFHQX1 Kt_reg_17_ ( .D(N2987), .CK(clk), .Q(Kt[17]) );
  DFFHQX1 Kt_reg_16_ ( .D(N2986), .CK(clk), .Q(Kt[16]) );
  DFFHQX1 H3_reg_2_ ( .D(n2681), .CK(clk), .Q(H3[2]) );
  DFFHQX1 H2_reg_2_ ( .D(n2650), .CK(clk), .Q(H2[2]) );
  DFFHQX1 H5_reg_2_ ( .D(n2745), .CK(clk), .Q(H5[2]) );
  DFFHQX1 H6_reg_2_ ( .D(n2617), .CK(clk), .Q(H6[2]) );
  DFFHQX1 H6_reg_3_ ( .D(n2616), .CK(clk), .Q(H6[3]) );
  DFFHQX1 H_reg_3_ ( .D(n2553), .CK(clk), .Q(SHA256_result[3]) );
  DFFHQX1 C_reg_4_ ( .D(n2871), .CK(clk), .Q(SHA256_result[164]) );
  DFFHQX1 B_reg_4_ ( .D(n2904), .CK(clk), .Q(SHA256_result[196]) );
  DFFHQX1 digest_reg_7_ ( .D(N3196), .CK(clk), .Q(digest[7]) );
  DFFHQX1 digest_reg_6_ ( .D(N3195), .CK(clk), .Q(digest[6]) );
  DFFHQX1 digest_reg_5_ ( .D(N3194), .CK(clk), .Q(digest[5]) );
  DFFHQX1 digest_reg_4_ ( .D(N3193), .CK(clk), .Q(digest[4]) );
  DFFHQX1 digest_reg_3_ ( .D(N3192), .CK(clk), .Q(digest[3]) );
  DFFHQX1 digest_reg_2_ ( .D(N3191), .CK(clk), .Q(digest[2]) );
  DFFHQX1 digest_reg_1_ ( .D(N3190), .CK(clk), .Q(digest[1]) );
  DFFHQX1 digest_reg_0_ ( .D(N3189), .CK(clk), .Q(digest[0]) );
  DFFHQX4 E_reg_25_ ( .D(n2786), .CK(clk), .Q(SHA256_result[121]) );
  DFFHQXL H3_reg_11_ ( .D(n2672), .CK(clk), .Q(H3[11]) );
  DFFHQXL H5_reg_10_ ( .D(n2737), .CK(clk), .Q(H5[10]) );
  DFFHQXL H2_reg_10_ ( .D(n2642), .CK(clk), .Q(H2[10]) );
  DFFHQXL H3_reg_10_ ( .D(n2673), .CK(clk), .Q(H3[10]) );
  DFFHQXL H_reg_23_ ( .D(n2533), .CK(clk), .Q(SHA256_result[23]) );
  DFFHQXL D_reg_1_ ( .D(n2842), .CK(clk), .Q(SHA256_result[129]) );
  DFFHQXL D_reg_0_ ( .D(n2843), .CK(clk), .Q(SHA256_result[128]) );
  DFFHQXL D_reg_2_ ( .D(n2841), .CK(clk), .Q(SHA256_result[130]) );
  DFFHQXL E_reg_21_ ( .D(n2790), .CK(clk), .Q(SHA256_result[117]) );
  DFFHQXL A_reg_12_ ( .D(n2960), .CK(clk), .Q(SHA256_result[236]) );
  DFFHQXL H3_reg_9_ ( .D(n2674), .CK(clk), .Q(H3[9]) );
  DFFHQXL H1_reg_8_ ( .D(n2932), .CK(clk), .Q(H1[8]) );
  DFFHQXL H2_reg_7_ ( .D(n2645), .CK(clk), .Q(H2[7]) );
  DFFHQXL H3_reg_7_ ( .D(n2676), .CK(clk), .Q(H3[7]) );
  DFFHQXL H2_reg_9_ ( .D(n2643), .CK(clk), .Q(H2[9]) );
  DFFHQXL H2_reg_8_ ( .D(n2644), .CK(clk), .Q(H2[8]) );
  DFFHQXL H3_reg_8_ ( .D(n2675), .CK(clk), .Q(H3[8]) );
  DFFHQXL A_reg_21_ ( .D(n2951), .CK(clk), .Q(SHA256_result[245]) );
  DFFHQXL A_reg_10_ ( .D(n2962), .CK(clk), .Q(SHA256_result[234]) );
  DFFHQXL A_reg_11_ ( .D(n2961), .CK(clk), .Q(SHA256_result[235]) );
  DFFHQXL A_reg_9_ ( .D(n2963), .CK(clk), .Q(SHA256_result[233]) );
  DFFHQXL A_reg_20_ ( .D(n2952), .CK(clk), .Q(SHA256_result[244]) );
  DFFHQXL A_reg_18_ ( .D(n2954), .CK(clk), .Q(SHA256_result[242]) );
  DFFHQXL A_reg_17_ ( .D(n2955), .CK(clk), .Q(SHA256_result[241]) );
  DFFHQXL A_reg_8_ ( .D(n2964), .CK(clk), .Q(SHA256_result[232]) );
  DFFHQXL A_reg_19_ ( .D(n2953), .CK(clk), .Q(SHA256_result[243]) );
  DFFHQXL A_reg_16_ ( .D(n2956), .CK(clk), .Q(SHA256_result[240]) );
  DFFHQXL E_reg_17_ ( .D(n2794), .CK(clk), .Q(SHA256_result[113]) );
  DFFHQXL A_reg_15_ ( .D(n2957), .CK(clk), .Q(SHA256_result[239]) );
  DFFHQXL H5_reg_6_ ( .D(n2741), .CK(clk), .Q(H5[6]) );
  DFFHQXL H1_reg_6_ ( .D(n2934), .CK(clk), .Q(H1[6]) );
  DFFHQXL H7_reg_5_ ( .D(n2519), .CK(clk), .Q(H7[5]) );
  DFFHQXL H2_reg_6_ ( .D(n2646), .CK(clk), .Q(H2[6]) );
  DFFHQXL H2_reg_5_ ( .D(n2647), .CK(clk), .Q(H2[5]) );
  DFFHQXL H3_reg_5_ ( .D(n2678), .CK(clk), .Q(H3[5]) );
  DFFHQXL H5_reg_4_ ( .D(n2743), .CK(clk), .Q(H5[4]) );
  DFFHQXL A_reg_13_ ( .D(n2959), .CK(clk), .Q(SHA256_result[237]) );
  DFFHQXL A_reg_14_ ( .D(n2958), .CK(clk), .Q(SHA256_result[238]) );
  DFFHQXL E_reg_15_ ( .D(n2796), .CK(clk), .Q(SHA256_result[111]) );
  DFFHQXL H2_reg_4_ ( .D(n2648), .CK(clk), .Q(H2[4]) );
  DFFHQXL H3_reg_4_ ( .D(n2679), .CK(clk), .Q(H3[4]) );
  DFFHQXL H2_reg_3_ ( .D(n2649), .CK(clk), .Q(H2[3]) );
  DFFHQX1 C_reg_11_ ( .D(n2864), .CK(clk), .Q(SHA256_result[171]) );
  DFFHQX1 G_reg_18_ ( .D(n2570), .CK(clk), .Q(SHA256_result[50]) );
  DFFHQX1 G_reg_19_ ( .D(n2569), .CK(clk), .Q(SHA256_result[51]) );
  DFFHQX1 H3_reg_6_ ( .D(n2677), .CK(clk), .Q(H3[6]) );
  DFFHQX1 H5_reg_5_ ( .D(n2742), .CK(clk), .Q(H5[5]) );
  DFFHQX1 H7_reg_4_ ( .D(n2520), .CK(clk), .Q(H7[4]) );
  DFFHQX1 H_reg_12_ ( .D(n2544), .CK(clk), .Q(SHA256_result[12]) );
  DFFHQX1 H_reg_7_ ( .D(n2549), .CK(clk), .Q(SHA256_result[7]) );
  DFFHQX1 H_reg_5_ ( .D(n2551), .CK(clk), .Q(SHA256_result[5]) );
  DFFHQX1 H1_reg_3_ ( .D(n2937), .CK(clk), .Q(H1[3]) );
  DFFHQX1 H3_reg_3_ ( .D(n2680), .CK(clk), .Q(H3[3]) );
  DFFHQX1 H5_reg_3_ ( .D(n2744), .CK(clk), .Q(H5[3]) );
  DFFHQX1 G_reg_10_ ( .D(n2578), .CK(clk), .Q(SHA256_result[42]) );
  DFFHQX1 B_reg_11_ ( .D(n2897), .CK(clk), .Q(SHA256_result[203]) );
  DFFHQX1 H_reg_8_ ( .D(n2548), .CK(clk), .Q(SHA256_result[8]) );
  DFFHQX1 H_reg_14_ ( .D(n2542), .CK(clk), .Q(SHA256_result[14]) );
  DFFHQX1 H_reg_11_ ( .D(n2545), .CK(clk), .Q(SHA256_result[11]) );
  DFFHQX1 F_reg_14_ ( .D(n2765), .CK(clk), .Q(SHA256_result[78]) );
  DFFHQX1 G_reg_14_ ( .D(n2574), .CK(clk), .Q(SHA256_result[46]) );
  DFFHQX1 C_reg_9_ ( .D(n2866), .CK(clk), .Q(SHA256_result[169]) );
  DFFHQX1 G_reg_16_ ( .D(n2572), .CK(clk), .Q(SHA256_result[48]) );
  DFFHQX1 B_reg_10_ ( .D(n2898), .CK(clk), .Q(SHA256_result[202]) );
  DFFHQX1 H_reg_4_ ( .D(n2552), .CK(clk), .Q(SHA256_result[4]) );
  DFFHQX1 F_reg_8_ ( .D(n2771), .CK(clk), .Q(SHA256_result[72]) );
  DFFHQX1 G_reg_8_ ( .D(n2580), .CK(clk), .Q(SHA256_result[40]) );
  DFFHQX1 G_reg_11_ ( .D(n2577), .CK(clk), .Q(SHA256_result[43]) );
  DFFHQXL D_reg_31_ ( .D(n2812), .CK(clk), .Q(SHA256_result[159]) );
  DFFHQXL B_reg_30_ ( .D(n2878), .CK(clk), .Q(SHA256_result[222]) );
  DFFHQXL C_reg_30_ ( .D(n2845), .CK(clk), .Q(SHA256_result[190]) );
  DFFHQXL C_reg_29_ ( .D(n2846), .CK(clk), .Q(SHA256_result[189]) );
  DFFHQX1 H3_reg_19_ ( .D(n2664), .CK(clk), .Q(H3[19]) );
  DFFHQXL H0_reg_31_ ( .D(n2973), .CK(clk), .Q(H0[31]) );
  DFFHQXL H1_reg_30_ ( .D(n2910), .CK(clk), .Q(H1[30]) );
  DFFHQXL H6_reg_30_ ( .D(n2589), .CK(clk), .Q(H6[30]) );
  DFFHQXL H2_reg_30_ ( .D(n2622), .CK(clk), .Q(H2[30]) );
  DFFHQXL H7_reg_30_ ( .D(n2494), .CK(clk), .Q(H7[30]) );
  DFFHQXL H4_reg_31_ ( .D(n2684), .CK(clk), .Q(H4[31]) );
  DFFHQXL H5_reg_30_ ( .D(n2717), .CK(clk), .Q(H5[30]) );
  DFFHQXL H3_reg_30_ ( .D(n2653), .CK(clk), .Q(H3[30]) );
  DFFHQXL H2_reg_31_ ( .D(n2621), .CK(clk), .Q(H2[31]) );
  DFFHQXL H6_reg_31_ ( .D(n2588), .CK(clk), .Q(H6[31]) );
  DFFHQXL H7_reg_31_ ( .D(n2493), .CK(clk), .Q(H7[31]) );
  DFFHQXL H1_reg_31_ ( .D(n2909), .CK(clk), .Q(H1[31]) );
  DFFHQXL H5_reg_31_ ( .D(n2716), .CK(clk), .Q(H5[31]) );
  DFFHQXL H3_reg_31_ ( .D(n2652), .CK(clk), .Q(H3[31]) );
  DFFHQXL H0_reg_28_ ( .D(n2976), .CK(clk), .Q(H0[28]) );
  DFFHQXL H4_reg_28_ ( .D(n2687), .CK(clk), .Q(H4[28]) );
  DFFHQXL H0_reg_29_ ( .D(n2975), .CK(clk), .Q(H0[29]) );
  DFFHQXL H4_reg_29_ ( .D(n2686), .CK(clk), .Q(H4[29]) );
  DFFHQXL H0_reg_30_ ( .D(n2974), .CK(clk), .Q(H0[30]) );
  DFFHQXL H4_reg_30_ ( .D(n2685), .CK(clk), .Q(H4[30]) );
  DFFHQXL H3_reg_27_ ( .D(n2656), .CK(clk), .Q(H3[27]) );
  DFFHQXL H5_reg_29_ ( .D(n2718), .CK(clk), .Q(H5[29]) );
  DFFHQXL H1_reg_27_ ( .D(n2913), .CK(clk), .Q(H1[27]) );
  DFFHQXL H1_reg_28_ ( .D(n2912), .CK(clk), .Q(H1[28]) );
  DFFHQXL H2_reg_28_ ( .D(n2624), .CK(clk), .Q(H2[28]) );
  DFFHQXL H3_reg_29_ ( .D(n2654), .CK(clk), .Q(H3[29]) );
  DFFHQXL H5_reg_28_ ( .D(n2719), .CK(clk), .Q(H5[28]) );
  DFFHQXL H6_reg_28_ ( .D(n2591), .CK(clk), .Q(H6[28]) );
  DFFHQXL H7_reg_27_ ( .D(n2497), .CK(clk), .Q(H7[27]) );
  DFFHQXL H7_reg_28_ ( .D(n2496), .CK(clk), .Q(H7[28]) );
  DFFHQXL H1_reg_29_ ( .D(n2911), .CK(clk), .Q(H1[29]) );
  DFFHQXL H2_reg_27_ ( .D(n2625), .CK(clk), .Q(H2[27]) );
  DFFHQXL H2_reg_29_ ( .D(n2623), .CK(clk), .Q(H2[29]) );
  DFFHQXL H0_reg_21_ ( .D(n2983), .CK(clk), .Q(H0[21]) );
  DFFHQXL H4_reg_23_ ( .D(n2692), .CK(clk), .Q(H4[23]) );
  DFFHQXL H4_reg_21_ ( .D(n2694), .CK(clk), .Q(H4[21]) );
  DFFHQXL H0_reg_23_ ( .D(n2981), .CK(clk), .Q(H0[23]) );
  DFFHQXL H0_reg_22_ ( .D(n2982), .CK(clk), .Q(H0[22]) );
  DFFHQXL H4_reg_26_ ( .D(n2689), .CK(clk), .Q(H4[26]) );
  DFFHQXL H4_reg_27_ ( .D(n2688), .CK(clk), .Q(H4[27]) );
  DFFHQXL H0_reg_27_ ( .D(n2977), .CK(clk), .Q(H0[27]) );
  DFFHQXL H0_reg_20_ ( .D(n2984), .CK(clk), .Q(H0[20]) );
  DFFHQXL D_reg_30_ ( .D(n2813), .CK(clk), .Q(SHA256_result[158]) );
  DFFHQXL H4_reg_22_ ( .D(n2693), .CK(clk), .Q(H4[22]) );
  DFFHQXL H4_reg_20_ ( .D(n2695), .CK(clk), .Q(H4[20]) );
  DFFHQXL H0_reg_26_ ( .D(n2978), .CK(clk), .Q(H0[26]) );
  DFFHQXL H0_reg_25_ ( .D(n2979), .CK(clk), .Q(H0[25]) );
  DFFHQXL H4_reg_24_ ( .D(n2691), .CK(clk), .Q(H4[24]) );
  DFFHQXL H0_reg_24_ ( .D(n2980), .CK(clk), .Q(H0[24]) );
  DFFHQXL H4_reg_25_ ( .D(n2690), .CK(clk), .Q(H4[25]) );
  DFFHQXL H2_reg_24_ ( .D(n2628), .CK(clk), .Q(H2[24]) );
  DFFHQXL H5_reg_26_ ( .D(n2721), .CK(clk), .Q(H5[26]) );
  DFFHQXL H1_reg_24_ ( .D(n2916), .CK(clk), .Q(H1[24]) );
  DFFHQXL H1_reg_25_ ( .D(n2915), .CK(clk), .Q(H1[25]) );
  DFFHQXL H2_reg_26_ ( .D(n2626), .CK(clk), .Q(H2[26]) );
  DFFHQXL H3_reg_24_ ( .D(n2659), .CK(clk), .Q(H3[24]) );
  DFFHQXL H3_reg_26_ ( .D(n2657), .CK(clk), .Q(H3[26]) );
  DFFHQXL H6_reg_26_ ( .D(n2593), .CK(clk), .Q(H6[26]) );
  DFFHQXL H7_reg_25_ ( .D(n2499), .CK(clk), .Q(H7[25]) );
  DFFHQXL H1_reg_26_ ( .D(n2914), .CK(clk), .Q(H1[26]) );
  DFFHQXL H3_reg_25_ ( .D(n2658), .CK(clk), .Q(H3[25]) );
  DFFHQXL H7_reg_24_ ( .D(n2500), .CK(clk), .Q(H7[24]) );
  DFFHQXL H5_reg_25_ ( .D(n2722), .CK(clk), .Q(H5[25]) );
  DFFHQXL H6_reg_25_ ( .D(n2594), .CK(clk), .Q(H6[25]) );
  DFFHQXL H4_reg_15_ ( .D(n2700), .CK(clk), .Q(H4[15]) );
  DFFHQXL H0_reg_17_ ( .D(n2987), .CK(clk), .Q(H0[17]) );
  DFFHQXL H0_reg_12_ ( .D(n2992), .CK(clk), .Q(H0[12]) );
  DFFHQXL H0_reg_15_ ( .D(n2989), .CK(clk), .Q(H0[15]) );
  DFFHQXL H4_reg_13_ ( .D(n2702), .CK(clk), .Q(H4[13]) );
  DFFHQXL H4_reg_16_ ( .D(n2699), .CK(clk), .Q(H4[16]) );
  DFFHQXL H4_reg_17_ ( .D(n2698), .CK(clk), .Q(H4[17]) );
  DFFHQXL H4_reg_19_ ( .D(n2696), .CK(clk), .Q(H4[19]) );
  DFFHQXL H4_reg_12_ ( .D(n2703), .CK(clk), .Q(H4[12]) );
  DFFHQXL H0_reg_18_ ( .D(n2986), .CK(clk), .Q(H0[18]) );
  DFFHQXL H4_reg_14_ ( .D(n2701), .CK(clk), .Q(H4[14]) );
  DFFHQXL H4_reg_18_ ( .D(n2697), .CK(clk), .Q(H4[18]) );
  DFFHQXL H0_reg_19_ ( .D(n2985), .CK(clk), .Q(H0[19]) );
  DFFHQXL H0_reg_14_ ( .D(n2990), .CK(clk), .Q(H0[14]) );
  DFFHQXL H0_reg_16_ ( .D(n2988), .CK(clk), .Q(H0[16]) );
  DFFHQXL D_reg_29_ ( .D(n2814), .CK(clk), .Q(SHA256_result[157]) );
  DFFHQXL H0_reg_13_ ( .D(n2991), .CK(clk), .Q(H0[13]) );
  DFFHQXL D_reg_25_ ( .D(n2818), .CK(clk), .Q(SHA256_result[153]) );
  DFFHQXL D_reg_28_ ( .D(n2815), .CK(clk), .Q(SHA256_result[156]) );
  DFFHQXL D_reg_26_ ( .D(n2817), .CK(clk), .Q(SHA256_result[154]) );
  DFFHQXL D_reg_27_ ( .D(n2816), .CK(clk), .Q(SHA256_result[155]) );
  DFFHQXL H5_reg_23_ ( .D(n2724), .CK(clk), .Q(H5[23]) );
  DFFHQXL H2_reg_22_ ( .D(n2630), .CK(clk), .Q(H2[22]) );
  DFFHQXL H3_reg_22_ ( .D(n2661), .CK(clk), .Q(H3[22]) );
  DFFHQXL H7_reg_23_ ( .D(n2501), .CK(clk), .Q(H7[23]) );
  DFFHQXL H1_reg_22_ ( .D(n2918), .CK(clk), .Q(H1[22]) );
  DFFHQXL H5_reg_24_ ( .D(n2723), .CK(clk), .Q(H5[24]) );
  DFFHQXL H6_reg_23_ ( .D(n2596), .CK(clk), .Q(H6[23]) );
  DFFHQXL H1_reg_23_ ( .D(n2917), .CK(clk), .Q(H1[23]) );
  DFFHQXL H2_reg_23_ ( .D(n2629), .CK(clk), .Q(H2[23]) );
  DFFHQXL H3_reg_23_ ( .D(n2660), .CK(clk), .Q(H3[23]) );
  DFFHQXL H4_reg_4_ ( .D(n2711), .CK(clk), .Q(H4[4]) );
  DFFHQXL H4_reg_3_ ( .D(n2712), .CK(clk), .Q(H4[3]) );
  DFFHQXL H4_reg_8_ ( .D(n2707), .CK(clk), .Q(H4[8]) );
  DFFHQXL H0_reg_6_ ( .D(n2998), .CK(clk), .Q(H0[6]) );
  DFFHQXL H0_reg_8_ ( .D(n2996), .CK(clk), .Q(H0[8]) );
  DFFHQXL H4_reg_11_ ( .D(n2704), .CK(clk), .Q(H4[11]) );
  DFFHQXL H0_reg_11_ ( .D(n2993), .CK(clk), .Q(H0[11]) );
  DFFHQXL H_reg_31_ ( .D(n2525), .CK(clk), .Q(SHA256_result[31]) );
  DFFHQXL H0_reg_9_ ( .D(n2995), .CK(clk), .Q(H0[9]) );
  DFFHQXL H0_reg_10_ ( .D(n2994), .CK(clk), .Q(H0[10]) );
  DFFHQXL H4_reg_10_ ( .D(n2705), .CK(clk), .Q(H4[10]) );
  DFFHQXL D_reg_23_ ( .D(n2820), .CK(clk), .Q(SHA256_result[151]) );
  DFFHQXL D_reg_22_ ( .D(n2821), .CK(clk), .Q(SHA256_result[150]) );
  DFFHQXL D_reg_21_ ( .D(n2822), .CK(clk), .Q(SHA256_result[149]) );
  DFFHQXL D_reg_20_ ( .D(n2823), .CK(clk), .Q(SHA256_result[148]) );
  DFFHQXL D_reg_24_ ( .D(n2819), .CK(clk), .Q(SHA256_result[152]) );
  DFFHQXL H1_reg_20_ ( .D(n2920), .CK(clk), .Q(H1[20]) );
  DFFHQXL H5_reg_20_ ( .D(n2727), .CK(clk), .Q(H5[20]) );
  DFFHQXL H6_reg_20_ ( .D(n2599), .CK(clk), .Q(H6[20]) );
  DFFHQXL H7_reg_20_ ( .D(n2504), .CK(clk), .Q(H7[20]) );
  DFFHQXL H3_reg_20_ ( .D(n2663), .CK(clk), .Q(H3[20]) );
  DFFHQXL H5_reg_22_ ( .D(n2725), .CK(clk), .Q(H5[22]) );
  DFFHQXL H6_reg_22_ ( .D(n2597), .CK(clk), .Q(H6[22]) );
  DFFHQXL H2_reg_21_ ( .D(n2631), .CK(clk), .Q(H2[21]) );
  DFFHQXL H7_reg_22_ ( .D(n2502), .CK(clk), .Q(H7[22]) );
  DFFHQXL H2_reg_19_ ( .D(n2633), .CK(clk), .Q(H2[19]) );
  DFFHQXL H2_reg_20_ ( .D(n2632), .CK(clk), .Q(H2[20]) );
  DFFHQXL H5_reg_21_ ( .D(n2726), .CK(clk), .Q(H5[21]) );
  DFFHQXL H6_reg_21_ ( .D(n2598), .CK(clk), .Q(H6[21]) );
  DFFHQXL H7_reg_19_ ( .D(n2505), .CK(clk), .Q(H7[19]) );
  DFFHQXL H1_reg_21_ ( .D(n2919), .CK(clk), .Q(H1[21]) );
  DFFHQXL H0_reg_0_ ( .D(n3004), .CK(clk), .Q(H0[0]) );
  DFFHQXL H0_reg_4_ ( .D(n3000), .CK(clk), .Q(H0[4]) );
  DFFHQXL H4_reg_0_ ( .D(n2715), .CK(clk), .Q(H4[0]) );
  DFFHQXL H4_reg_1_ ( .D(n2714), .CK(clk), .Q(H4[1]) );
  DFFHQXL H4_reg_5_ ( .D(n2710), .CK(clk), .Q(H4[5]) );
  DFFHQXL H0_reg_3_ ( .D(n3001), .CK(clk), .Q(H0[3]) );
  DFFHQXL H0_reg_7_ ( .D(n2997), .CK(clk), .Q(H0[7]) );
  DFFHQXL H4_reg_7_ ( .D(n2708), .CK(clk), .Q(H4[7]) );
  DFFHQXL H0_reg_2_ ( .D(n3002), .CK(clk), .Q(H0[2]) );
  DFFHQXL H4_reg_2_ ( .D(n2713), .CK(clk), .Q(H4[2]) );
  DFFHQXL H_reg_30_ ( .D(n2526), .CK(clk), .Q(SHA256_result[30]) );
  DFFHQXL D_reg_17_ ( .D(n2826), .CK(clk), .Q(SHA256_result[145]) );
  DFFHQXL D_reg_18_ ( .D(n2825), .CK(clk), .Q(SHA256_result[146]) );
  DFFHQXL D_reg_19_ ( .D(n2824), .CK(clk), .Q(SHA256_result[147]) );
  DFFHQXL D_reg_13_ ( .D(n2830), .CK(clk), .Q(SHA256_result[141]) );
  DFFHQXL D_reg_10_ ( .D(n2833), .CK(clk), .Q(SHA256_result[138]) );
  DFFHQXL D_reg_11_ ( .D(n2832), .CK(clk), .Q(SHA256_result[139]) );
  DFFHQXL D_reg_16_ ( .D(n2827), .CK(clk), .Q(SHA256_result[144]) );
  DFFHQXL B_reg_29_ ( .D(n2879), .CK(clk), .Q(SHA256_result[221]) );
  DFFHQXL B_reg_28_ ( .D(n2880), .CK(clk), .Q(SHA256_result[220]) );
  DFFHQXL D_reg_15_ ( .D(n2828), .CK(clk), .Q(SHA256_result[143]) );
  DFFHQXL H6_reg_18_ ( .D(n2601), .CK(clk), .Q(H6[18]) );
  DFFHQXL H7_reg_17_ ( .D(n2507), .CK(clk), .Q(H7[17]) );
  DFFHQXL H7_reg_18_ ( .D(n2506), .CK(clk), .Q(H7[18]) );
  DFFHQXL H1_reg_16_ ( .D(n2924), .CK(clk), .Q(H1[16]) );
  DFFHQXL H1_reg_18_ ( .D(n2922), .CK(clk), .Q(H1[18]) );
  DFFHQXL H6_reg_17_ ( .D(n2602), .CK(clk), .Q(H6[17]) );
  DFFHQXL H2_reg_17_ ( .D(n2635), .CK(clk), .Q(H2[17]) );
  DFFHQXL H2_reg_18_ ( .D(n2634), .CK(clk), .Q(H2[18]) );
  DFFHQXL H5_reg_18_ ( .D(n2729), .CK(clk), .Q(H5[18]) );
  DFFHQXL H3_reg_18_ ( .D(n2665), .CK(clk), .Q(H3[18]) );
  DFFHQXL H5_reg_17_ ( .D(n2730), .CK(clk), .Q(H5[17]) );
  DFFHQXL H5_reg_19_ ( .D(n2728), .CK(clk), .Q(H5[19]) );
  DFFHQXL H_reg_28_ ( .D(n2528), .CK(clk), .Q(SHA256_result[28]) );
  DFFHQXL H_reg_29_ ( .D(n2527), .CK(clk), .Q(SHA256_result[29]) );
  DFFHQXL D_reg_9_ ( .D(n2834), .CK(clk), .Q(SHA256_result[137]) );
  DFFHQXL D_reg_14_ ( .D(n2829), .CK(clk), .Q(SHA256_result[142]) );
  DFFHQXL D_reg_8_ ( .D(n2835), .CK(clk), .Q(SHA256_result[136]) );
  DFFHQXL C_reg_26_ ( .D(n2849), .CK(clk), .Q(SHA256_result[186]) );
  DFFHQXL C_reg_24_ ( .D(n2851), .CK(clk), .Q(SHA256_result[184]) );
  DFFHQXL G_reg_30_ ( .D(n2558), .CK(clk), .Q(SHA256_result[62]) );
  DFFHQXL D_reg_12_ ( .D(n2831), .CK(clk), .Q(SHA256_result[140]) );
  DFFHQXL B_reg_27_ ( .D(n2881), .CK(clk), .Q(SHA256_result[219]) );
  DFFHQXL B_reg_26_ ( .D(n2882), .CK(clk), .Q(SHA256_result[218]) );
  DFFHQXL C_reg_27_ ( .D(n2848), .CK(clk), .Q(SHA256_result[187]) );
  DFFHQXL F_reg_30_ ( .D(n2749), .CK(clk), .Q(SHA256_result[94]) );
  DFFHQXL H7_reg_16_ ( .D(n2508), .CK(clk), .Q(H7[16]) );
  DFFHQXL H1_reg_15_ ( .D(n2925), .CK(clk), .Q(H1[15]) );
  DFFHQXL H5_reg_16_ ( .D(n2731), .CK(clk), .Q(H5[16]) );
  DFFHQXL H6_reg_15_ ( .D(n2604), .CK(clk), .Q(H6[15]) );
  DFFHQXL H6_reg_16_ ( .D(n2603), .CK(clk), .Q(H6[16]) );
  DFFHQXL H7_reg_14_ ( .D(n2510), .CK(clk), .Q(H7[14]) );
  DFFHQXL H7_reg_15_ ( .D(n2509), .CK(clk), .Q(H7[15]) );
  DFFHQXL H2_reg_15_ ( .D(n2637), .CK(clk), .Q(H2[15]) );
  DFFHQXL H3_reg_16_ ( .D(n2667), .CK(clk), .Q(H3[16]) );
  DFFHQXL H1_reg_14_ ( .D(n2926), .CK(clk), .Q(H1[14]) );
  DFFHQXL H2_reg_16_ ( .D(n2636), .CK(clk), .Q(H2[16]) );
  DFFHQXL H5_reg_15_ ( .D(n2732), .CK(clk), .Q(H5[15]) );
  DFFHQXL H_reg_24_ ( .D(n2532), .CK(clk), .Q(SHA256_result[24]) );
  DFFHQXL H_reg_26_ ( .D(n2530), .CK(clk), .Q(SHA256_result[26]) );
  DFFHQXL D_reg_4_ ( .D(n2839), .CK(clk), .Q(SHA256_result[132]) );
  DFFHQXL H_reg_27_ ( .D(n2529), .CK(clk), .Q(SHA256_result[27]) );
  DFFHQXL D_reg_5_ ( .D(n2838), .CK(clk), .Q(SHA256_result[133]) );
  DFFHQXL G_reg_28_ ( .D(n2560), .CK(clk), .Q(SHA256_result[60]) );
  DFFHQXL G_reg_27_ ( .D(n2561), .CK(clk), .Q(SHA256_result[59]) );
  DFFHQXL D_reg_7_ ( .D(n2836), .CK(clk), .Q(SHA256_result[135]) );
  DFFHQXL D_reg_6_ ( .D(n2837), .CK(clk), .Q(SHA256_result[134]) );
  DFFHQXL C_reg_22_ ( .D(n2853), .CK(clk), .Q(SHA256_result[182]) );
  DFFHQXL C_reg_25_ ( .D(n2850), .CK(clk), .Q(SHA256_result[185]) );
  DFFHQXL B_reg_22_ ( .D(n2886), .CK(clk), .Q(SHA256_result[214]) );
  DFFHQXL F_reg_28_ ( .D(n2751), .CK(clk), .Q(SHA256_result[92]) );
  DFFHQXL C_reg_23_ ( .D(n2852), .CK(clk), .Q(SHA256_result[183]) );
  DFFHQXL C_reg_20_ ( .D(n2855), .CK(clk), .Q(SHA256_result[180]) );
  DFFHQXL B_reg_23_ ( .D(n2885), .CK(clk), .Q(SHA256_result[215]) );
  DFFHQXL B_reg_24_ ( .D(n2884), .CK(clk), .Q(SHA256_result[216]) );
  DFFHQXL B_reg_20_ ( .D(n2888), .CK(clk), .Q(SHA256_result[212]) );
  DFFTRX1 round_reg_0_ ( .D(N145), .RN(n141), .CK(clk), .Q(n366), .QN(n1396)
         );
  DFFHQXL H5_reg_12_ ( .D(n2735), .CK(clk), .Q(H5[12]) );
  DFFHQXL H6_reg_13_ ( .D(n2606), .CK(clk), .Q(H6[13]) );
  DFFHQXL H7_reg_12_ ( .D(n2512), .CK(clk), .Q(H7[12]) );
  DFFHQXL H1_reg_11_ ( .D(n2929), .CK(clk), .Q(H1[11]) );
  DFFHQXL H1_reg_13_ ( .D(n2927), .CK(clk), .Q(H1[13]) );
  DFFHQXL H5_reg_14_ ( .D(n2733), .CK(clk), .Q(H5[14]) );
  DFFHQXL H6_reg_12_ ( .D(n2607), .CK(clk), .Q(H6[12]) );
  DFFHQXL H6_reg_14_ ( .D(n2605), .CK(clk), .Q(H6[14]) );
  DFFHQXL H2_reg_13_ ( .D(n2639), .CK(clk), .Q(H2[13]) );
  DFFHQXL H2_reg_14_ ( .D(n2638), .CK(clk), .Q(H2[14]) );
  DFFHQXL H3_reg_14_ ( .D(n2669), .CK(clk), .Q(H3[14]) );
  DFFHQXL H3_reg_15_ ( .D(n2668), .CK(clk), .Q(H3[15]) );
  DFFHQXL H3_reg_12_ ( .D(n2671), .CK(clk), .Q(H3[12]) );
  DFFHQXL H1_reg_12_ ( .D(n2928), .CK(clk), .Q(H1[12]) );
  DFFHQXL H_reg_25_ ( .D(n2531), .CK(clk), .Q(SHA256_result[25]) );
  DFFHQXL H_reg_20_ ( .D(n2536), .CK(clk), .Q(SHA256_result[20]) );
  DFFHQXL H_reg_21_ ( .D(n2535), .CK(clk), .Q(SHA256_result[21]) );
  DFFHQXL C_reg_18_ ( .D(n2857), .CK(clk), .Q(SHA256_result[178]) );
  DFFHQXL D_reg_3_ ( .D(n2840), .CK(clk), .Q(SHA256_result[131]) );
  DFFHQXL H_reg_22_ ( .D(n2534), .CK(clk), .Q(SHA256_result[22]) );
  DFFHQXL G_reg_24_ ( .D(n2564), .CK(clk), .Q(SHA256_result[56]) );
  DFFHQXL F_reg_26_ ( .D(n2753), .CK(clk), .Q(SHA256_result[90]) );
  DFFHQXL G_reg_25_ ( .D(n2563), .CK(clk), .Q(SHA256_result[57]) );
  DFFHQXL B_reg_18_ ( .D(n2890), .CK(clk), .Q(SHA256_result[210]) );
  DFFHQXL B_reg_19_ ( .D(n2889), .CK(clk), .Q(SHA256_result[211]) );
  DFFHQXL F_reg_25_ ( .D(n2754), .CK(clk), .Q(SHA256_result[89]) );
  DFFHQXL B_reg_21_ ( .D(n2887), .CK(clk), .Q(SHA256_result[213]) );
  DFFHQXL E_reg_10_ ( .D(n2801), .CK(clk), .Q(SHA256_result[106]) );
  DFFHQXL H4_reg_6_ ( .D(n2709), .CK(clk), .Q(H4[6]) );
  DFFHQXL H4_reg_9_ ( .D(n2706), .CK(clk), .Q(H4[9]) );
  DFFHQXL H0_reg_1_ ( .D(n3003), .CK(clk), .Q(H0[1]) );
  DFFHQXL H0_reg_5_ ( .D(n2999), .CK(clk), .Q(H0[5]) );
  DFFHQX1 H_reg_13_ ( .D(n2543), .CK(clk), .Q(SHA256_result[13]) );
  DFFHQX1 H_reg_9_ ( .D(n2547), .CK(clk), .Q(SHA256_result[9]) );
  DFFHQX1 H_reg_2_ ( .D(n2554), .CK(clk), .Q(SHA256_result[2]) );
  DFFHQX1 G_reg_17_ ( .D(n2571), .CK(clk), .Q(SHA256_result[49]) );
  DFFX4 C_reg_1_ ( .D(n2874), .CK(clk), .Q(n121), .QN(n122) );
  DFFHQXL H2_reg_11_ ( .D(n2641), .CK(clk), .Q(H2[11]) );
  DFFHQXL H7_reg_11_ ( .D(n2513), .CK(clk), .Q(H7[11]) );
  DFFHQXL H5_reg_11_ ( .D(n2736), .CK(clk), .Q(H5[11]) );
  DFFHQXL H3_reg_13_ ( .D(n2670), .CK(clk), .Q(H3[13]) );
  DFFHQXL H2_reg_12_ ( .D(n2640), .CK(clk), .Q(H2[12]) );
  DFFHQXL H_reg_19_ ( .D(n2537), .CK(clk), .Q(SHA256_result[19]) );
  DFFHQXL C_reg_15_ ( .D(n2860), .CK(clk), .Q(SHA256_result[175]) );
  DFFHQXL F_reg_23_ ( .D(n2756), .CK(clk), .Q(SHA256_result[87]) );
  DFFHQXL G_reg_23_ ( .D(n2565), .CK(clk), .Q(SHA256_result[55]) );
  DFFHQXL C_reg_16_ ( .D(n2859), .CK(clk), .Q(SHA256_result[176]) );
  DFFHQXL B_reg_17_ ( .D(n2891), .CK(clk), .Q(SHA256_result[209]) );
  DFFHQXL B_reg_15_ ( .D(n2893), .CK(clk), .Q(SHA256_result[207]) );
  DFFHQXL B_reg_16_ ( .D(n2892), .CK(clk), .Q(SHA256_result[208]) );
  DFFHQX1 G_reg_12_ ( .D(n2576), .CK(clk), .Q(SHA256_result[44]) );
  DFFHQX4 B_reg_1_ ( .D(n2907), .CK(clk), .Q(SHA256_result[193]) );
  DFFHQXL C_reg_31_ ( .D(n2844), .CK(clk), .Q(SHA256_result[191]) );
  DFFHQX1 H7_reg_3_ ( .D(n2521), .CK(clk), .Q(H7[3]) );
  DFFHQX1 H6_reg_27_ ( .D(n2592), .CK(clk), .Q(H6[27]) );
  DFFHQX1 F_reg_27_ ( .D(n2752), .CK(clk), .Q(SHA256_result[91]) );
  DFFHQX1 G_reg_31_ ( .D(n2557), .CK(clk), .Q(SHA256_result[63]) );
  DFFHQXL F_reg_31_ ( .D(n2748), .CK(clk), .Q(SHA256_result[95]) );
  DFFHQX4 H7_reg_0_ ( .D(n2524), .CK(clk), .Q(H7[0]) );
  DFFX4 H3_reg_0_ ( .D(n2683), .CK(clk), .Q(n108) );
  DFFX4 A_reg_1_ ( .D(n2971), .CK(clk), .Q(n106), .QN(n107) );
  DFFHQXL B_reg_31_ ( .D(n2877), .CK(clk), .Q(SHA256_result[223]) );
  DFFX4 A_reg_0_ ( .D(n2972), .CK(clk), .Q(n97), .QN(n98) );
  DFFHQX1 H3_reg_17_ ( .D(n2666), .CK(clk), .Q(H3[17]) );
  DFFHQXL H6_reg_10_ ( .D(n2609), .CK(clk), .Q(H6[10]) );
  DFFX4 H7_reg_1_ ( .D(n2523), .CK(clk), .Q(n92) );
  DFFHQX1 H7_reg_21_ ( .D(n2503), .CK(clk), .Q(H7[21]) );
  DFFHQX1 H6_reg_24_ ( .D(n2595), .CK(clk), .Q(H6[24]) );
  DFFHQXL H5_reg_9_ ( .D(n2738), .CK(clk), .Q(H5[9]) );
  DFFHQX1 G_reg_21_ ( .D(n2567), .CK(clk), .Q(SHA256_result[53]) );
  DFFTRX1 round_reg_5_ ( .D(N150), .RN(n141), .CK(clk), .Q(round[5]), .QN(
        n1370) );
  DFFHQX1 H5_reg_8_ ( .D(n2739), .CK(clk), .Q(H5[8]) );
  DFFHQX1 H6_reg_9_ ( .D(n2610), .CK(clk), .Q(H6[9]) );
  DFFHQX1 H7_reg_9_ ( .D(n2515), .CK(clk), .Q(H7[9]) );
  DFFHQX1 H1_reg_7_ ( .D(n2933), .CK(clk), .Q(H1[7]) );
  DFFHQX1 H1_reg_9_ ( .D(n2931), .CK(clk), .Q(H1[9]) );
  DFFHQX1 H5_reg_7_ ( .D(n2740), .CK(clk), .Q(H5[7]) );
  DFFHQX1 H6_reg_8_ ( .D(n2611), .CK(clk), .Q(H6[8]) );
  DFFHQX1 H7_reg_8_ ( .D(n2516), .CK(clk), .Q(H7[8]) );
  DFFHQX1 H7_reg_10_ ( .D(n2514), .CK(clk), .Q(H7[10]) );
  DFFHQX1 G_reg_22_ ( .D(n2566), .CK(clk), .Q(SHA256_result[54]) );
  DFFHQX1 F_reg_22_ ( .D(n2757), .CK(clk), .Q(SHA256_result[86]) );
  DFFHQX1 E_reg_24_ ( .D(n2787), .CK(clk), .Q(SHA256_result[120]) );
  DFFHQX1 H1_reg_5_ ( .D(n2935), .CK(clk), .Q(H1[5]) );
  DFFHQX1 H6_reg_6_ ( .D(n2613), .CK(clk), .Q(H6[6]) );
  DFFHQX1 H7_reg_6_ ( .D(n2518), .CK(clk), .Q(H7[6]) );
  DFFHQX1 H7_reg_7_ ( .D(n2517), .CK(clk), .Q(H7[7]) );
  DFFHQX1 H6_reg_7_ ( .D(n2612), .CK(clk), .Q(H6[7]) );
  DFFHQX1 H_reg_6_ ( .D(n2550), .CK(clk), .Q(SHA256_result[6]) );
  DFFHQX1 C_reg_7_ ( .D(n2868), .CK(clk), .Q(SHA256_result[167]) );
  DFFHQX1 H_reg_1_ ( .D(n2555), .CK(clk), .Q(SHA256_result[1]) );
  DFFHQX1 C_reg_14_ ( .D(n2861), .CK(clk), .Q(SHA256_result[174]) );
  DFFHQX1 E_reg_22_ ( .D(n2789), .CK(clk), .Q(SHA256_result[118]) );
  DFFHQX1 E_reg_9_ ( .D(n2802), .CK(clk), .Q(SHA256_result[105]) );
  DFFHQX1 C_reg_6_ ( .D(n2869), .CK(clk), .Q(SHA256_result[166]) );
  DFFHQX1 B_reg_7_ ( .D(n2901), .CK(clk), .Q(SHA256_result[199]) );
  DFFHQX1 E_reg_6_ ( .D(n2805), .CK(clk), .Q(SHA256_result[102]) );
  DFFHQX1 E_reg_12_ ( .D(n2799), .CK(clk), .Q(SHA256_result[108]) );
  DFFHQX1 E_reg_8_ ( .D(n2803), .CK(clk), .Q(SHA256_result[104]) );
  DFFHQX4 H6_reg_0_ ( .D(n2619), .CK(clk), .Q(H6[0]) );
  DFFHQX4 H6_reg_1_ ( .D(n2618), .CK(clk), .Q(H6[1]) );
  DFFHQX4 H3_reg_1_ ( .D(n2682), .CK(clk), .Q(H3[1]) );
  DFFX4 G_reg_0_ ( .D(n2620), .CK(clk), .Q(n88), .QN(n87) );
  DFFX4 G_reg_1_ ( .D(n2587), .CK(clk), .Q(n84), .QN(n83) );
  DFFX4 C_reg_0_ ( .D(n2875), .CK(clk), .Q(n71), .QN(n70) );
  DFFX4 F_reg_1_ ( .D(n2778), .CK(clk), .Q(n66), .QN(n67) );
  DFFHQX4 H2_reg_0_ ( .D(n2876), .CK(clk), .Q(H2[0]) );
  DFFX4 E_reg_0_ ( .D(n2811), .CK(clk), .Q(n65), .QN(n64) );
  DFFHQX4 F_reg_4_ ( .D(n2775), .CK(clk), .Q(SHA256_result[68]) );
  DFFHQX2 H2_reg_1_ ( .D(n2651), .CK(clk), .Q(H2[1]) );
  DFFHQX4 E_reg_31_ ( .D(n2780), .CK(clk), .Q(SHA256_result[127]) );
  DFFHQX4 A_reg_31_ ( .D(n2941), .CK(clk), .Q(SHA256_result[255]) );
  DFFHQXL C_reg_28_ ( .D(n2847), .CK(clk), .Q(SHA256_result[188]) );
  DFFHQXL C_reg_19_ ( .D(n2856), .CK(clk), .Q(SHA256_result[179]) );
  DFFHQXL H_reg_10_ ( .D(n2546), .CK(clk), .Q(SHA256_result[10]) );
  DFFHQX1 G_reg_7_ ( .D(n2581), .CK(clk), .Q(SHA256_result[39]) );
  DFFHQX1 F_reg_13_ ( .D(n2766), .CK(clk), .Q(SHA256_result[77]) );
  DFFHQXL C_reg_21_ ( .D(n2854), .CK(clk), .Q(SHA256_result[181]) );
  DFFHQXL C_reg_17_ ( .D(n2858), .CK(clk), .Q(SHA256_result[177]) );
  DFFHQXL F_reg_24_ ( .D(n2755), .CK(clk), .Q(SHA256_result[88]) );
  DFFHQXL C_reg_12_ ( .D(n2863), .CK(clk), .Q(SHA256_result[172]) );
  DFFTRX1 round_reg_4_ ( .D(N149), .RN(n141), .CK(clk), .Q(n371), .QN(n369) );
  DFFTRX1 round_reg_1_ ( .D(N146), .RN(n141), .CK(clk), .Q(n368), .QN(n373) );
  DFFTRX2 round_reg_3_ ( .D(N148), .RN(n141), .CK(clk), .Q(round[3]), .QN(
        n1383) );
  DFFTRX2 round_reg_2_ ( .D(N147), .RN(n141), .CK(clk), .Q(round[2]), .QN(
        n1388) );
  DFFHQX2 B_reg_2_ ( .D(n2906), .CK(clk), .Q(SHA256_result[194]) );
  DFFHQX1 B_reg_3_ ( .D(n2905), .CK(clk), .Q(SHA256_result[195]) );
  DFFHQX2 E_reg_16_ ( .D(n2795), .CK(clk), .Q(SHA256_result[112]) );
  DFFHQX2 E_reg_26_ ( .D(n2785), .CK(clk), .Q(SHA256_result[122]) );
  DFFHQX2 E_reg_28_ ( .D(n2783), .CK(clk), .Q(SHA256_result[124]) );
  DFFHQX2 F_reg_2_ ( .D(n2777), .CK(clk), .Q(SHA256_result[66]) );
  DFFHQX2 G_reg_5_ ( .D(n2583), .CK(clk), .Q(SHA256_result[37]) );
  DFFHQX2 Kt_reg_15_ ( .D(N2985), .CK(clk), .Q(Kt[15]) );
  DFFHQX2 Kt_reg_14_ ( .D(N2984), .CK(clk), .Q(Kt[14]) );
  DFFHQX2 Kt_reg_11_ ( .D(N2981), .CK(clk), .Q(Kt[11]) );
  DFFHQX2 Kt_reg_9_ ( .D(N2979), .CK(clk), .Q(Kt[9]) );
  DFFHQX2 Kt_reg_8_ ( .D(N2978), .CK(clk), .Q(Kt[8]) );
  DFFHQX2 Kt_reg_7_ ( .D(N2977), .CK(clk), .Q(Kt[7]) );
  DFFHQX2 Kt_reg_5_ ( .D(N2975), .CK(clk), .Q(Kt[5]) );
  DFFHQX2 Kt_reg_4_ ( .D(N2974), .CK(clk), .Q(Kt[4]) );
  DFFHQX1 H_reg_0_ ( .D(n2556), .CK(clk), .Q(SHA256_result[0]) );
  DFFX2 C_reg_2_ ( .D(n2873), .CK(clk), .Q(n94), .QN(n95) );
  DFFHQX1 E_reg_23_ ( .D(n2788), .CK(clk), .Q(SHA256_result[119]) );
  DFFX2 H7_reg_2_ ( .D(n2522), .CK(clk), .Q(n91) );
  DFFX2 H1_reg_0_ ( .D(n2940), .CK(clk), .Q(n90) );
  DFFHQX1 H1_reg_17_ ( .D(n2923), .CK(clk), .Q(H1[17]) );
  DFFHQX1 B_reg_6_ ( .D(n2902), .CK(clk), .Q(SHA256_result[198]) );
  DFFHQX1 H6_reg_5_ ( .D(n2614), .CK(clk), .Q(H6[5]) );
  DFFHQX1 H5_reg_27_ ( .D(n2720), .CK(clk), .Q(H5[27]) );
  DFFHQX2 E_reg_27_ ( .D(n2784), .CK(clk), .Q(SHA256_result[123]) );
  DFFHQX1 H5_reg_13_ ( .D(n2734), .CK(clk), .Q(H5[13]) );
  DFFHQX1 H7_reg_29_ ( .D(n2495), .CK(clk), .Q(H7[29]) );
  DFFHQXL G_reg_29_ ( .D(n2559), .CK(clk), .Q(SHA256_result[61]) );
  DFFHQX1 H1_reg_10_ ( .D(n2930), .CK(clk), .Q(H1[10]) );
  DFFHQX1 H6_reg_19_ ( .D(n2600), .CK(clk), .Q(H6[19]) );
  DFFHQX1 F_reg_19_ ( .D(n2760), .CK(clk), .Q(SHA256_result[83]) );
  DFFHQX1 H7_reg_26_ ( .D(n2498), .CK(clk), .Q(H7[26]) );
  DFFHQX1 G_reg_26_ ( .D(n2562), .CK(clk), .Q(SHA256_result[58]) );
  DFFHQX1 H6_reg_29_ ( .D(n2590), .CK(clk), .Q(H6[29]) );
  DFFHQX1 F_reg_29_ ( .D(n2750), .CK(clk), .Q(SHA256_result[93]) );
  DFFHQX2 A_reg_22_ ( .D(n2950), .CK(clk), .Q(SHA256_result[246]) );
  DFFHQX1 F_reg_9_ ( .D(n2770), .CK(clk), .Q(SHA256_result[73]) );
  DFFHQX2 G_reg_4_ ( .D(n2584), .CK(clk), .Q(SHA256_result[36]) );
  DFFHQX2 H1_reg_1_ ( .D(n2939), .CK(clk), .Q(H1[1]) );
  DFFHQX1 H1_reg_2_ ( .D(n2938), .CK(clk), .Q(H1[2]) );
  DFFHQX1 H2_reg_25_ ( .D(n2627), .CK(clk), .Q(H2[25]) );
  DFFHQX1 B_reg_25_ ( .D(n2883), .CK(clk), .Q(SHA256_result[217]) );
  DFFHQX1 H7_reg_13_ ( .D(n2511), .CK(clk), .Q(H7[13]) );
  DFFHQX1 H3_reg_21_ ( .D(n2662), .CK(clk), .Q(H3[21]) );
  DFFHQX1 H1_reg_19_ ( .D(n2921), .CK(clk), .Q(H1[19]) );
  DFFHQX1 H3_reg_28_ ( .D(n2655), .CK(clk), .Q(H3[28]) );
  DFFHQX1 H1_reg_4_ ( .D(n2936), .CK(clk), .Q(H1[4]) );
  DFFHQX1 H6_reg_11_ ( .D(n2608), .CK(clk), .Q(H6[11]) );
  DFFHQX2 F_reg_11_ ( .D(n2768), .CK(clk), .Q(SHA256_result[75]) );
  DFFHQX1 G_reg_9_ ( .D(n2579), .CK(clk), .Q(SHA256_result[41]) );
  EDFFTRX1 round_reg_6_ ( .RN(N151), .D(n141), .E(1'b1), .CK(clk), .Q(round[6]), .QN(n380) );
  DFFHQX1 E_reg_20_ ( .D(n2791), .CK(clk), .Q(SHA256_result[116]) );
  DFFHQX2 H5_reg_1_ ( .D(n2746), .CK(clk), .Q(H5[1]) );
  DFFHQX4 F_reg_6_ ( .D(n2773), .CK(clk), .Q(SHA256_result[70]) );
  DFFHQX4 H5_reg_0_ ( .D(n2747), .CK(clk), .Q(H5[0]) );
  DFFHQXL E_reg_29_ ( .D(n2782), .CK(clk), .Q(SHA256_result[125]) );
  DFFHQX4 F_reg_10_ ( .D(n2769), .CK(clk), .Q(SHA256_result[74]) );
  DFFHQX2 C_reg_3_ ( .D(n2872), .CK(clk), .Q(SHA256_result[163]) );
  DFFHQX4 E_reg_5_ ( .D(n2806), .CK(clk), .Q(SHA256_result[101]) );
  DFFHQXL A_reg_28_ ( .D(n2944), .CK(clk), .Q(SHA256_result[252]) );
  DFFHQX4 E_reg_3_ ( .D(n2808), .CK(clk), .Q(SHA256_result[99]) );
  DFFHQX4 F_reg_5_ ( .D(n2774), .CK(clk), .Q(SHA256_result[69]) );
  DFFHQXL G_reg_13_ ( .D(n2575), .CK(clk), .Q(SHA256_result[45]) );
  DFFHQX4 F_reg_12_ ( .D(n2767), .CK(clk), .Q(SHA256_result[76]) );
  DFFHQX4 G_reg_6_ ( .D(n2582), .CK(clk), .Q(SHA256_result[38]) );
  DFFHQX2 F_reg_7_ ( .D(n2772), .CK(clk), .Q(SHA256_result[71]) );
  DFFHQX4 E_reg_14_ ( .D(n2797), .CK(clk), .Q(SHA256_result[110]) );
  DFFHQX2 E_reg_18_ ( .D(n2793), .CK(clk), .Q(SHA256_result[114]) );
  CLKINVX3 U3 ( .A(SHA256_result[98]), .Y(n76) );
  INVX1 U4 ( .A(SHA256_result[37]), .Y(n436) );
  INVX2 U5 ( .A(n1436), .Y(n46) );
  AOI21XL U15 ( .A0(N887), .A1(n237), .B0(n272), .Y(n1749) );
  AOI21XL U16 ( .A0(N888), .A1(n234), .B0(n272), .Y(n1748) );
  AOI21XL U17 ( .A0(N864), .A1(n238), .B0(n272), .Y(n1772) );
  AOI21XL U18 ( .A0(N878), .A1(n11), .B0(n272), .Y(n1758) );
  AOI21XL U19 ( .A0(N872), .A1(n11), .B0(n272), .Y(n1764) );
  XNOR3X2 U20 ( .A(n15), .B(SHA256_result[109]), .C(n892), .Y(f4_E_32[7]) );
  INVX1 U21 ( .A(SHA256_result[114]), .Y(n892) );
  OAI2BB1X4 U22 ( .A0N(N973), .A1N(n238), .B0(n462), .Y(n2785) );
  INVXL U23 ( .A(n179), .Y(n701) );
  OAI2BB1X1 U24 ( .A0N(SHA256_result[194]), .A1N(n179), .B0(n607), .Y(
        f2_ABC_32[2]) );
  NAND3X2 U25 ( .A(n454), .B(n453), .C(n452), .Y(n2783) );
  NAND2X2 U26 ( .A(N975), .B(n241), .Y(n452) );
  OAI211XL U27 ( .A0(n361), .A1(n440), .B0(n48), .C0(n1538), .Y(n2616) );
  INVX1 U28 ( .A(SHA256_result[35]), .Y(n440) );
  BUFX12 U29 ( .A(T1_32[13]), .Y(n10) );
  OAI2BB1X4 U30 ( .A0N(N974), .A1N(n234), .B0(n458), .Y(n2784) );
  NAND2X4 U31 ( .A(n40), .B(n41), .Y(f1_EFG_32[7]) );
  OAI211X4 U32 ( .A0(n337), .A1(n39), .B0(n415), .C0(n414), .Y(n2772) );
  INVX12 U33 ( .A(n245), .Y(n11) );
  INVX20 U34 ( .A(n710), .Y(n713) );
  INVX2 U35 ( .A(n246), .Y(n232) );
  INVX12 U36 ( .A(n245), .Y(n235) );
  INVX12 U37 ( .A(n244), .Y(n242) );
  INVX2 U38 ( .A(n38), .Y(n236) );
  INVX3 U39 ( .A(n244), .Y(n243) );
  INVX12 U40 ( .A(n245), .Y(n234) );
  CLKINVX3 U41 ( .A(n38), .Y(n241) );
  INVX4 U42 ( .A(n245), .Y(n231) );
  INVX4 U43 ( .A(n245), .Y(n240) );
  INVX2 U44 ( .A(n244), .Y(n238) );
  MX2X4 U45 ( .A(SHA256_result[42]), .B(SHA256_result[74]), .S0(n149), .Y(
        f1_EFG_32[10]) );
  BUFX8 U46 ( .A(SHA256_result[106]), .Y(n149) );
  OAI211X4 U47 ( .A0(n337), .A1(n441), .B0(n401), .C0(n400), .Y(n2586) );
  NAND2XL U48 ( .A(n441), .B(SHA256_result[98]), .Y(n78) );
  OAI211XL U49 ( .A0(n361), .A1(n441), .B0(n48), .C0(n1608), .Y(n2745) );
  INVX4 U50 ( .A(SHA256_result[66]), .Y(n441) );
  MX2X4 U51 ( .A(SHA256_result[44]), .B(SHA256_result[76]), .S0(n148), .Y(
        f1_EFG_32[12]) );
  CLKBUFX8 U52 ( .A(SHA256_result[45]), .Y(n12) );
  OAI21X1 U53 ( .A0(n183), .A1(n923), .B0(n1611), .Y(n2750) );
  INVX8 U54 ( .A(SHA256_result[69]), .Y(n435) );
  XOR2X4 U55 ( .A(SHA256_result[127]), .B(n42), .Y(f4_E_32[6]) );
  NAND2X4 U56 ( .A(n24), .B(n1754), .Y(n2877) );
  MXI2X4 U57 ( .A(n440), .B(n439), .S0(SHA256_result[99]), .Y(f1_EFG_32[3]) );
  INVX12 U58 ( .A(n1455), .Y(n280) );
  INVX2 U59 ( .A(n1455), .Y(n281) );
  INVX16 U60 ( .A(n279), .Y(n353) );
  INVX12 U61 ( .A(n279), .Y(n352) );
  INVX8 U62 ( .A(n339), .Y(n340) );
  INVX12 U63 ( .A(n278), .Y(n342) );
  INVX8 U64 ( .A(n276), .Y(n347) );
  INVX12 U65 ( .A(n277), .Y(n349) );
  INVX2 U66 ( .A(n275), .Y(n341) );
  INVX12 U67 ( .A(n275), .Y(n345) );
  INVX2 U68 ( .A(n275), .Y(n343) );
  INVX12 U69 ( .A(n277), .Y(n348) );
  INVX12 U70 ( .A(n278), .Y(n350) );
  INVX12 U71 ( .A(n278), .Y(n351) );
  INVX3 U72 ( .A(n292), .Y(n287) );
  INVX3 U73 ( .A(n293), .Y(n284) );
  INVX4 U74 ( .A(n291), .Y(n290) );
  INVX3 U75 ( .A(n292), .Y(n289) );
  INVX4 U76 ( .A(n294), .Y(n288) );
  INVX4 U77 ( .A(n294), .Y(n286) );
  INVX4 U78 ( .A(n293), .Y(n285) );
  INVX4 U79 ( .A(n295), .Y(n283) );
  OR3X1 U80 ( .A(n1848), .B(n378), .C(n377), .Y(n1455) );
  INVX4 U81 ( .A(n280), .Y(n279) );
  CLKINVX2 U82 ( .A(n280), .Y(n278) );
  CLKINVX3 U83 ( .A(n282), .Y(n339) );
  INVX4 U84 ( .A(n281), .Y(n276) );
  INVX4 U85 ( .A(n281), .Y(n277) );
  INVX4 U86 ( .A(n281), .Y(n275) );
  CLKINVX3 U87 ( .A(n353), .Y(n291) );
  CLKINVX3 U88 ( .A(n353), .Y(n292) );
  CLKINVX3 U89 ( .A(n353), .Y(n293) );
  CLKINVX3 U90 ( .A(n352), .Y(n294) );
  CLKINVX3 U91 ( .A(n352), .Y(n295) );
  CLKINVX3 U92 ( .A(n340), .Y(n338) );
  CLKINVX3 U93 ( .A(n340), .Y(n337) );
  CLKINVX3 U94 ( .A(n351), .Y(n299) );
  CLKINVX3 U95 ( .A(n351), .Y(n298) );
  CLKINVX3 U96 ( .A(n347), .Y(n315) );
  CLKINVX3 U97 ( .A(n347), .Y(n316) );
  CLKINVX3 U98 ( .A(n347), .Y(n317) );
  CLKINVX3 U99 ( .A(n349), .Y(n309) );
  CLKINVX3 U100 ( .A(n349), .Y(n308) );
  CLKINVX3 U101 ( .A(n349), .Y(n307) );
  CLKINVX3 U102 ( .A(n288), .Y(n96) );
  CLKINVX3 U103 ( .A(n341), .Y(n334) );
  CLKINVX3 U104 ( .A(n341), .Y(n335) );
  CLKINVX3 U105 ( .A(n341), .Y(n336) );
  CLKINVX3 U106 ( .A(n345), .Y(n324) );
  CLKINVX3 U107 ( .A(n345), .Y(n325) );
  CLKINVX3 U108 ( .A(n345), .Y(n326) );
  INVXL U109 ( .A(n346), .Y(n323) );
  CLKINVX3 U110 ( .A(n348), .Y(n311) );
  CLKINVX3 U111 ( .A(n348), .Y(n310) );
  CLKBUFX8 U112 ( .A(SHA256_result[252]), .Y(n13) );
  AOI22X1 U113 ( .A0(N1021), .A1(n239), .B0(SHA256_result[74]), .B1(n342), .Y(
        n1513) );
  CLKBUFX8 U114 ( .A(SHA256_result[125]), .Y(n14) );
  XOR3X4 U115 ( .A(n151), .B(SHA256_result[109]), .C(SHA256_result[123]), .Y(
        f4_E_32[2]) );
  MX2X4 U116 ( .A(SHA256_result[40]), .B(SHA256_result[72]), .S0(n151), .Y(
        f1_EFG_32[8]) );
  CLKBUFX8 U117 ( .A(SHA256_result[104]), .Y(n151) );
  OAI211X4 U118 ( .A0(n307), .A1(n62), .B0(n428), .C0(n427), .Y(n2778) );
  OAI211X4 U119 ( .A0(n360), .A1(n62), .B0(n51), .C0(n1594), .Y(n2714) );
  INVX8 U120 ( .A(n62), .Y(n63) );
  CLKINVX8 U121 ( .A(SHA256_result[97]), .Y(n62) );
  MX2X4 U122 ( .A(SHA256_result[38]), .B(SHA256_result[70]), .S0(n152), .Y(
        f1_EFG_32[6]) );
  AOI22X1 U123 ( .A0(N1017), .A1(n233), .B0(SHA256_result[70]), .B1(n349), .Y(
        n1517) );
  OAI21X4 U124 ( .A0(n186), .A1(n852), .B0(n1723), .Y(n2845) );
  NAND2X4 U125 ( .A(n119), .B(n1722), .Y(n2844) );
  INVX8 U126 ( .A(n57), .Y(n58) );
  CLKINVX8 U127 ( .A(n97), .Y(n57) );
  MXI2X4 U128 ( .A(n436), .B(n435), .S0(SHA256_result[101]), .Y(f1_EFG_32[5])
         );
  BUFX8 U129 ( .A(n20), .Y(n15) );
  BUFX20 U130 ( .A(n63), .Y(n61) );
  INVX8 U131 ( .A(n18), .Y(n19) );
  INVXL U132 ( .A(n18), .Y(n20) );
  CLKINVX8 U133 ( .A(n65), .Y(n18) );
  INVX1 U134 ( .A(n388), .Y(n1456) );
  OAI211X1 U135 ( .A0(n356), .A1(n930), .B0(n48), .C0(n1534), .Y(n2608) );
  NAND2X2 U136 ( .A(N1009), .B(n232), .Y(n102) );
  XOR3X2 U137 ( .A(SHA256_result[107]), .B(SHA256_result[112]), .C(n143), .Y(
        f4_E_32[5]) );
  CLKINVX4 U138 ( .A(n79), .Y(f1_EFG_32[2]) );
  NAND2X2 U139 ( .A(n77), .B(n78), .Y(n79) );
  XOR3X2 U140 ( .A(SHA256_result[103]), .B(n148), .C(SHA256_result[122]), .Y(
        f4_E_32[1]) );
  MXI2X2 U141 ( .A(n83), .B(n67), .S0(n61), .Y(f1_EFG_32[1]) );
  NAND2X1 U142 ( .A(SHA256_result[71]), .B(SHA256_result[103]), .Y(n41) );
  NAND2X1 U143 ( .A(SHA256_result[39]), .B(n39), .Y(n40) );
  OAI2BB1X1 U144 ( .A0N(SHA256_result[192]), .A1N(n59), .B0(n609), .Y(
        f2_ABC_32[0]) );
  XOR3X2 U145 ( .A(n179), .B(n168), .C(SHA256_result[246]), .Y(f3_A_32[0]) );
  INVX1 U146 ( .A(n381), .Y(n36) );
  INVX1 U147 ( .A(first_block), .Y(n35) );
  NAND2X1 U148 ( .A(n1858), .B(n380), .Y(n378) );
  NAND2BX1 U149 ( .AN(n1848), .B(output_enable), .Y(n1490) );
  NAND2BX1 U150 ( .AN(n1858), .B(round[6]), .Y(n376) );
  INVX1 U151 ( .A(n1490), .Y(n377) );
  BUFX12 U152 ( .A(n106), .Y(n60) );
  BUFX4 U153 ( .A(SHA256_result[105]), .Y(n150) );
  CLKBUFX8 U154 ( .A(SHA256_result[102]), .Y(n152) );
  BUFX3 U155 ( .A(SHA256_result[248]), .Y(n158) );
  BUFX3 U156 ( .A(SHA256_result[247]), .Y(n159) );
  BUFX3 U157 ( .A(SHA256_result[237]), .Y(n168) );
  CLKINVX3 U158 ( .A(SHA256_result[68]), .Y(n437) );
  BUFX4 U159 ( .A(SHA256_result[243]), .Y(n162) );
  CLKBUFX8 U160 ( .A(SHA256_result[241]), .Y(n164) );
  CLKBUFX8 U161 ( .A(SHA256_result[242]), .Y(n163) );
  BUFX3 U162 ( .A(SHA256_result[244]), .Y(n161) );
  BUFX3 U163 ( .A(SHA256_result[233]), .Y(n172) );
  BUFX3 U164 ( .A(SHA256_result[235]), .Y(n170) );
  BUFX4 U165 ( .A(SHA256_result[234]), .Y(n171) );
  BUFX4 U166 ( .A(SHA256_result[245]), .Y(n160) );
  BUFX3 U167 ( .A(next_A[21]), .Y(n33) );
  BUFX3 U168 ( .A(SHA256_result[115]), .Y(n145) );
  CLKBUFX8 U169 ( .A(SHA256_result[226]), .Y(n179) );
  CLKBUFX8 U170 ( .A(SHA256_result[229]), .Y(n176) );
  CLKBUFX8 U171 ( .A(SHA256_result[232]), .Y(n173) );
  CLKBUFX8 U172 ( .A(SHA256_result[113]), .Y(n146) );
  BUFX3 U173 ( .A(SHA256_result[111]), .Y(n147) );
  INVX2 U174 ( .A(SHA256_result[36]), .Y(n438) );
  INVX8 U175 ( .A(n22), .Y(n364) );
  BUFX3 U176 ( .A(SHA256_result[231]), .Y(n174) );
  BUFX3 U177 ( .A(SHA256_result[230]), .Y(n175) );
  BUFX3 U178 ( .A(SHA256_result[117]), .Y(n144) );
  BUFX3 U179 ( .A(SHA256_result[238]), .Y(n167) );
  BUFX3 U180 ( .A(SHA256_result[236]), .Y(n169) );
  NOR2X1 U181 ( .A(n788), .B(n182), .Y(n1877) );
  NOR2X1 U182 ( .A(n793), .B(n181), .Y(n2225) );
  BUFX3 U183 ( .A(round[5]), .Y(n181) );
  OAI2BB1X1 U184 ( .A0N(n713), .A1N(N976), .B0(n450), .Y(n2782) );
  OAI221XL U185 ( .A0(n315), .A1(n920), .B0(n229), .B1(n945), .C0(n1497), .Y(
        n2562) );
  NAND2X1 U186 ( .A(H5[0]), .B(n254), .Y(n429) );
  AND2X2 U187 ( .A(n111), .B(n112), .Y(n1493) );
  NAND3X2 U188 ( .A(n68), .B(n69), .C(n1457), .Y(n2526) );
  OR2X2 U189 ( .A(n1456), .B(n982), .Y(n69) );
  OR2X2 U190 ( .A(n293), .B(n949), .Y(n68) );
  NAND2X2 U191 ( .A(n113), .B(n1453), .Y(n2525) );
  NAND2X1 U192 ( .A(n73), .B(n1755), .Y(n2878) );
  AND2X2 U193 ( .A(n74), .B(n75), .Y(n1755) );
  OAI221XL U194 ( .A0(n291), .A1(n905), .B0(n226), .B1(n930), .C0(n1512), .Y(
        n2577) );
  OAI21XL U195 ( .A0(n364), .A1(n435), .B0(n416), .Y(n2742) );
  NAND3X2 U196 ( .A(n444), .B(n445), .C(n446), .Y(n2781) );
  OAI221XL U197 ( .A0(n318), .A1(n890), .B0(n227), .B1(n910), .C0(n1624), .Y(
        n2763) );
  NAND2X1 U198 ( .A(n26), .B(n615), .Y(n2943) );
  NAND2X1 U199 ( .A(N844), .B(n11), .Y(n628) );
  OAI2BB1X1 U200 ( .A0N(N843), .A1N(n236), .B0(n634), .Y(n2948) );
  OAI221XL U201 ( .A0(n292), .A1(n808), .B0(n217), .B1(n835), .C0(n1740), .Y(
        n2862) );
  OAI2BB1X1 U202 ( .A0N(N963), .A1N(n242), .B0(n488), .Y(n2795) );
  NAND2X1 U203 ( .A(N961), .B(n11), .Y(n491) );
  NAND2X2 U204 ( .A(n23), .B(n620), .Y(n2945) );
  NAND2X4 U205 ( .A(N846), .B(n242), .Y(n620) );
  CLKINVX3 U206 ( .A(n1436), .Y(n47) );
  OR2X2 U207 ( .A(n377), .B(n129), .Y(n710) );
  CLKINVX2 U208 ( .A(n47), .Y(n55) );
  INVX1 U209 ( .A(n47), .Y(n54) );
  INVX1 U210 ( .A(n47), .Y(n56) );
  INVX1 U211 ( .A(n46), .Y(n52) );
  CLKINVX3 U212 ( .A(n246), .Y(n239) );
  INVX1 U213 ( .A(n274), .Y(n267) );
  INVX1 U214 ( .A(n206), .Y(n200) );
  INVX1 U215 ( .A(n46), .Y(n48) );
  CLKINVX3 U216 ( .A(n246), .Y(n233) );
  INVX1 U217 ( .A(n46), .Y(n49) );
  INVX1 U218 ( .A(n46), .Y(n51) );
  INVX1 U219 ( .A(n46), .Y(n50) );
  INVX1 U220 ( .A(n37), .Y(n237) );
  INVX8 U221 ( .A(n262), .Y(n258) );
  INVX1 U222 ( .A(n140), .Y(n671) );
  NOR2BX1 U223 ( .AN(first_block), .B(n1489), .Y(n140) );
  INVX1 U224 ( .A(n47), .Y(n53) );
  INVX1 U225 ( .A(n131), .Y(n765) );
  CLKINVX3 U226 ( .A(n198), .Y(n184) );
  INVX1 U227 ( .A(n273), .Y(n269) );
  NOR3X2 U228 ( .A(n1848), .B(round[6]), .C(n258), .Y(n138) );
  INVX1 U229 ( .A(n258), .Y(n247) );
  NOR2X1 U230 ( .A(n1370), .B(n369), .Y(n21) );
  NOR2X1 U231 ( .A(first_block), .B(n361), .Y(n22) );
  INVX1 U232 ( .A(n34), .Y(n199) );
  AND2X2 U233 ( .A(n621), .B(n622), .Y(n23) );
  AND2X2 U234 ( .A(n105), .B(n104), .Y(n24) );
  AND2X2 U235 ( .A(n613), .B(n614), .Y(n25) );
  AND2X2 U236 ( .A(n616), .B(n617), .Y(n26) );
  INVX1 U237 ( .A(n87), .Y(n89) );
  AND2X2 U238 ( .A(n81), .B(n82), .Y(n27) );
  INVX1 U239 ( .A(n354), .Y(n363) );
  NOR2X1 U240 ( .A(n1370), .B(n180), .Y(n28) );
  AND2X2 U241 ( .A(n2183), .B(n2174), .Y(n29) );
  INVX1 U242 ( .A(SHA256_result[103]), .Y(n39) );
  BUFX16 U243 ( .A(SHA256_result[100]), .Y(n43) );
  CLKINVX3 U244 ( .A(n43), .Y(n80) );
  INVX1 U245 ( .A(n70), .Y(n72) );
  NOR2X1 U246 ( .A(n1383), .B(round[2]), .Y(n137) );
  NOR2XL U247 ( .A(n1383), .B(n1388), .Y(n2303) );
  AOI21X1 U249 ( .A0(N896), .A1(n236), .B0(n271), .Y(n1740) );
  AOI21X1 U250 ( .A0(N897), .A1(n233), .B0(n271), .Y(n1739) );
  AOI21X1 U251 ( .A0(N892), .A1(n234), .B0(n271), .Y(n1744) );
  AOI21X1 U252 ( .A0(N891), .A1(n233), .B0(n271), .Y(n1745) );
  AOI21X1 U253 ( .A0(N889), .A1(n237), .B0(n271), .Y(n1747) );
  AOI21X1 U254 ( .A0(N993), .A1(n237), .B0(n269), .Y(n1626) );
  AOI21X1 U255 ( .A0(N992), .A1(n240), .B0(n269), .Y(n1627) );
  AOI21X1 U256 ( .A0(N1054), .A1(n242), .B0(n268), .Y(n1477) );
  AOI21X1 U257 ( .A0(N1058), .A1(n233), .B0(n268), .Y(n1473) );
  AOI21X1 U258 ( .A0(N1057), .A1(n231), .B0(n268), .Y(n1474) );
  AOI21X1 U259 ( .A0(N1051), .A1(n11), .B0(n268), .Y(n1480) );
  AOI21X1 U260 ( .A0(N1037), .A1(n240), .B0(n268), .Y(n1497) );
  NAND2X4 U261 ( .A(N946), .B(n233), .Y(n120) );
  AOI21XL U262 ( .A0(N1071), .A1(n237), .B0(n268), .Y(n1460) );
  AOI21XL U263 ( .A0(N1068), .A1(n11), .B0(n270), .Y(n1463) );
  AOI21XL U264 ( .A0(N1070), .A1(n241), .B0(n272), .Y(n1461) );
  AOI21XL U265 ( .A0(N939), .A1(n243), .B0(n269), .Y(n1697) );
  AOI21XL U266 ( .A0(N941), .A1(n242), .B0(n269), .Y(n1695) );
  AOI21XL U267 ( .A0(N937), .A1(n233), .B0(n269), .Y(n1699) );
  NAND2X2 U268 ( .A(n25), .B(n612), .Y(n2942) );
  NAND2X2 U269 ( .A(N849), .B(n11), .Y(n612) );
  AOI2BB2X4 U270 ( .B0(N914), .B1(n242), .A0N(n794), .A1N(n305), .Y(n1722) );
  AOI21XL U271 ( .A0(N1035), .A1(n235), .B0(n269), .Y(n1499) );
  AOI21XL U272 ( .A0(N997), .A1(n234), .B0(n272), .Y(n1622) );
  AOI21XL U273 ( .A0(N1003), .A1(n238), .B0(n269), .Y(n1616) );
  AOI21XL U274 ( .A0(N1026), .A1(n232), .B0(n269), .Y(n1508) );
  AOI21XL U275 ( .A0(N1036), .A1(n241), .B0(n268), .Y(n1498) );
  AOI21XL U276 ( .A0(N1038), .A1(n236), .B0(n268), .Y(n1496) );
  AOI21XL U277 ( .A0(N1039), .A1(n243), .B0(n268), .Y(n1495) );
  AOI21XL U278 ( .A0(N905), .A1(n713), .B0(n271), .Y(n1731) );
  AOI21XL U279 ( .A0(N904), .A1(n237), .B0(n271), .Y(n1732) );
  AOI21XL U280 ( .A0(N895), .A1(n235), .B0(n271), .Y(n1741) );
  BUFX8 U281 ( .A(T1_32[7]), .Y(n31) );
  AOI21X1 U282 ( .A0(n143), .A1(n208), .B0(n496), .Y(n446) );
  INVX12 U283 ( .A(SHA256_result[64]), .Y(n443) );
  AOI21XL U284 ( .A0(N995), .A1(n237), .B0(n269), .Y(n1624) );
  AOI21XL U285 ( .A0(N932), .A1(n238), .B0(n266), .Y(n1704) );
  AOI21XL U286 ( .A0(N934), .A1(n238), .B0(n270), .Y(n1702) );
  AOI21XL U287 ( .A0(N933), .A1(n238), .B0(n269), .Y(n1703) );
  AOI21XL U288 ( .A0(N931), .A1(n241), .B0(n269), .Y(n1705) );
  AOI21XL U289 ( .A0(N944), .A1(n231), .B0(n269), .Y(n1692) );
  BUFX8 U290 ( .A(next_E[20]), .Y(n32) );
  NAND2X4 U291 ( .A(N977), .B(n237), .Y(n444) );
  NAND2X4 U292 ( .A(N1041), .B(n236), .Y(n111) );
  NAND2BX1 U293 ( .AN(n361), .B(first_block), .Y(n1436) );
  CLKINVX3 U294 ( .A(n138), .Y(n361) );
  OAI211X1 U295 ( .A0(n361), .A1(n83), .B0(n51), .C0(n1539), .Y(n2618) );
  OAI211X1 U296 ( .A0(n361), .A1(n439), .B0(n49), .C0(n1607), .Y(n2744) );
  OAI211X2 U297 ( .A0(n480), .A1(n293), .B0(n479), .C0(n478), .Y(n2792) );
  AOI21X1 U298 ( .A0(n35), .A1(n36), .B0(n377), .Y(n34) );
  MX2X4 U299 ( .A(n12), .B(SHA256_result[77]), .S0(SHA256_result[109]), .Y(
        f1_EFG_32[13]) );
  INVXL U300 ( .A(n713), .Y(n37) );
  INVXL U301 ( .A(n713), .Y(n38) );
  NAND2X2 U302 ( .A(N848), .B(n241), .Y(n615) );
  OAI2BB1X4 U303 ( .A0N(n232), .A1N(N978), .B0(n549), .Y(n2780) );
  OAI2BB1X4 U304 ( .A0N(n243), .A1N(N850), .B0(n611), .Y(n2941) );
  XOR2X1 U305 ( .A(n146), .B(n148), .Y(n42) );
  NAND2X2 U306 ( .A(N913), .B(n713), .Y(n125) );
  BUFX3 U307 ( .A(n45), .Y(n44) );
  INVX1 U308 ( .A(n46), .Y(n45) );
  CLKINVX2 U309 ( .A(n57), .Y(n59) );
  NAND2XL U310 ( .A(H7[0]), .B(n256), .Y(n1452) );
  OAI211X1 U311 ( .A0(n294), .A1(n437), .B0(n396), .C0(n395), .Y(n2584) );
  MX2X4 U312 ( .A(SHA256_result[41]), .B(SHA256_result[73]), .S0(n150), .Y(
        f1_EFG_32[9]) );
  OAI21X1 U313 ( .A0(n178), .A1(SHA256_result[195]), .B0(SHA256_result[163]), 
        .Y(n606) );
  OAI2BB1X2 U314 ( .A0N(SHA256_result[195]), .A1N(n178), .B0(n606), .Y(
        f2_ABC_32[3]) );
  NOR2X1 U315 ( .A(n367), .B(n182), .Y(n131) );
  INVXL U316 ( .A(next_E[9]), .Y(n512) );
  XOR3X4 U317 ( .A(n152), .B(SHA256_result[107]), .C(SHA256_result[121]), .Y(
        f4_E_32[0]) );
  AND2X4 U318 ( .A(n116), .B(n671), .Y(n1457) );
  NAND2XL U319 ( .A(N1073), .B(n231), .Y(n116) );
  OR2X2 U320 ( .A(n184), .B(n825), .Y(n73) );
  NAND2X4 U321 ( .A(N881), .B(n11), .Y(n74) );
  NAND2XL U322 ( .A(n153), .B(n350), .Y(n75) );
  NAND2X2 U323 ( .A(n442), .B(n76), .Y(n77) );
  INVXL U324 ( .A(SHA256_result[34]), .Y(n442) );
  NAND2X4 U325 ( .A(n438), .B(n80), .Y(n81) );
  NAND2X4 U326 ( .A(n437), .B(n43), .Y(n82) );
  INVX1 U327 ( .A(n83), .Y(n85) );
  MXI2X4 U328 ( .A(n87), .B(n443), .S0(n15), .Y(f1_EFG_32[0]) );
  INVXL U329 ( .A(n443), .Y(n86) );
  NAND2X4 U330 ( .A(N1074), .B(n231), .Y(n114) );
  OAI211XL U331 ( .A0(n358), .A1(n856), .B0(n52), .C0(n1579), .Y(n2682) );
  AND2X4 U332 ( .A(n114), .B(n115), .Y(n1453) );
  NAND3X4 U333 ( .A(n127), .B(n128), .C(n1690), .Y(n2812) );
  NAND2XL U334 ( .A(N945), .B(n237), .Y(n100) );
  AOI2BB2X4 U335 ( .B0(N1042), .B1(n234), .A0N(n899), .A1N(n303), .Y(n1492) );
  INVX1 U336 ( .A(n198), .Y(n185) );
  OAI2BB1X1 U337 ( .A0N(n188), .A1N(SHA256_result[94]), .B0(n1610), .Y(n2749)
         );
  AND2X2 U338 ( .A(n102), .B(n103), .Y(n1610) );
  NAND2XL U339 ( .A(SHA256_result[63]), .B(n285), .Y(n115) );
  OAI21XL U340 ( .A0(n179), .A1(SHA256_result[194]), .B0(n94), .Y(n607) );
  NAND2X1 U341 ( .A(n99), .B(n1691), .Y(n2813) );
  AND2X2 U342 ( .A(n100), .B(n101), .Y(n1691) );
  AOI21X4 U343 ( .A0(N882), .A1(n242), .B0(n272), .Y(n1754) );
  OR2XL U344 ( .A(n185), .B(n885), .Y(n99) );
  NAND2X1 U345 ( .A(SHA256_result[190]), .B(n286), .Y(n101) );
  AOI21XL U346 ( .A0(n209), .A1(SHA256_result[95]), .B0(n266), .Y(n433) );
  NAND2XL U347 ( .A(n143), .B(n287), .Y(n103) );
  AND2X4 U348 ( .A(n125), .B(n126), .Y(n1723) );
  OR2X2 U349 ( .A(n311), .B(n735), .Y(n104) );
  OR2X2 U350 ( .A(n219), .B(n794), .Y(n105) );
  OAI211XL U351 ( .A0(n355), .A1(n952), .B0(n53), .C0(n1452), .Y(n2524) );
  NAND2X4 U352 ( .A(n1492), .B(n118), .Y(n2557) );
  NAND2X1 U353 ( .A(N912), .B(n240), .Y(n117) );
  OAI211X2 U354 ( .A0(n310), .A1(n547), .B0(n433), .C0(n432), .Y(n2748) );
  NAND2X4 U355 ( .A(N1010), .B(n235), .Y(n432) );
  OAI2BB2XL U356 ( .B0(n364), .B1(n855), .A0N(n108), .A1N(n261), .Y(n2683) );
  INVXL U357 ( .A(n34), .Y(n198) );
  NOR2XL U358 ( .A(n187), .B(n640), .Y(n641) );
  AND2X2 U359 ( .A(n117), .B(n671), .Y(n1724) );
  NAND3X1 U360 ( .A(n123), .B(n124), .C(n1724), .Y(n2846) );
  NAND2XL U361 ( .A(SHA256_result[222]), .B(n351), .Y(n126) );
  NAND2X1 U362 ( .A(n110), .B(n1493), .Y(n2558) );
  OR2XL U363 ( .A(n186), .B(n949), .Y(n110) );
  NAND2X1 U364 ( .A(SHA256_result[94]), .B(n347), .Y(n112) );
  OR2X2 U365 ( .A(n740), .B(n951), .Y(n113) );
  INVX1 U366 ( .A(n273), .Y(n270) );
  INVX1 U367 ( .A(n199), .Y(n186) );
  BUFX12 U368 ( .A(SHA256_result[228]), .Y(n177) );
  OAI2BB1X1 U369 ( .A0N(SHA256_result[193]), .A1N(n60), .B0(n608), .Y(
        f2_ABC_32[1]) );
  OAI21XL U370 ( .A0(SHA256_result[193]), .A1(n60), .B0(n121), .Y(n608) );
  OR2X2 U371 ( .A(n186), .B(n950), .Y(n118) );
  OR2X2 U372 ( .A(n186), .B(n853), .Y(n119) );
  CLKINVX3 U373 ( .A(n273), .Y(n272) );
  INVXL U374 ( .A(SHA256_result[67]), .Y(n439) );
  AND2X4 U375 ( .A(n120), .B(n671), .Y(n1690) );
  INVX1 U376 ( .A(n212), .Y(n209) );
  CLKINVX3 U377 ( .A(n363), .Y(n355) );
  INVXL U378 ( .A(n140), .Y(n274) );
  NOR2XL U379 ( .A(n131), .B(n2215), .Y(n2473) );
  NAND2X1 U380 ( .A(N834), .B(n243), .Y(n657) );
  NAND2X1 U381 ( .A(N838), .B(n240), .Y(n647) );
  OAI211X1 U382 ( .A0(n649), .A1(n304), .B0(n648), .C0(n647), .Y(n2953) );
  NAND2X1 U383 ( .A(N833), .B(n237), .Y(n660) );
  NAND2X1 U384 ( .A(N964), .B(n231), .Y(n484) );
  NAND2X1 U385 ( .A(N957), .B(n11), .Y(n505) );
  NAND2X1 U386 ( .A(N835), .B(n232), .Y(n654) );
  NAND2X1 U387 ( .A(N832), .B(n11), .Y(n663) );
  NAND2X1 U388 ( .A(N831), .B(n235), .Y(n666) );
  NAND2XL U389 ( .A(n190), .B(n169), .Y(n667) );
  NAND2X1 U390 ( .A(N828), .B(n237), .Y(n676) );
  NAND2XL U391 ( .A(N821), .B(n236), .Y(n703) );
  NAND2XL U392 ( .A(N824), .B(n233), .Y(n689) );
  NAND2XL U393 ( .A(N823), .B(n237), .Y(n693) );
  INVXL U394 ( .A(n137), .Y(n789) );
  AOI211XL U395 ( .A0(n757), .A1(round[2]), .B0(n2291), .C0(n2292), .Y(n2290)
         );
  AOI221XL U396 ( .A0(n2221), .A1(n372), .B0(n131), .B1(n21), .C0(n2292), .Y(
        n2337) );
  AOI211XL U397 ( .A0(n757), .A1(n137), .B0(n2240), .C0(n2241), .Y(n2230) );
  AOI21XL U398 ( .A0(n137), .A1(n2427), .B0(n2228), .Y(n2233) );
  AOI21XL U399 ( .A0(n209), .A1(SHA256_result[110]), .B0(n267), .Y(n492) );
  NAND2X1 U400 ( .A(N965), .B(n238), .Y(n481) );
  NAND2X1 U401 ( .A(N971), .B(n240), .Y(n467) );
  OAI2BB2X1 U402 ( .B0(n364), .B1(n861), .A0N(H3[6]), .A1N(n261), .Y(n2677) );
  AOI22X1 U403 ( .A0(N906), .A1(n232), .B0(SHA256_result[215]), .B1(n344), .Y(
        n1730) );
  BUFX8 U404 ( .A(SHA256_result[126]), .Y(n143) );
  BUFX8 U405 ( .A(SHA256_result[250]), .Y(n156) );
  NAND2XL U406 ( .A(N1012), .B(n243), .Y(n403) );
  NAND2XL U407 ( .A(N947), .B(n236), .Y(n544) );
  NAND2XL U408 ( .A(N981), .B(n239), .Y(n425) );
  NAND2XL U409 ( .A(N982), .B(n238), .Y(n423) );
  NAND2XL U410 ( .A(N984), .B(n243), .Y(n417) );
  NAND2XL U411 ( .A(N980), .B(n240), .Y(n427) );
  OAI211X1 U412 ( .A0(n295), .A1(n435), .B0(n393), .C0(n392), .Y(n2583) );
  OAI211X1 U413 ( .A0(n314), .A1(n439), .B0(n398), .C0(n397), .Y(n2585) );
  OAI21XL U414 ( .A0(SHA256_result[201]), .A1(n172), .B0(SHA256_result[169]), 
        .Y(n600) );
  BUFX8 U415 ( .A(SHA256_result[254]), .Y(n153) );
  BUFX3 U416 ( .A(n366), .Y(n182) );
  MX2X1 U417 ( .A(SHA256_result[51]), .B(SHA256_result[83]), .S0(n145), .Y(
        f1_EFG_32[19]) );
  AOI222XL U418 ( .A0(n131), .A1(n2199), .B0(n2272), .B1(n373), .C0(n2381), 
        .C1(n1396), .Y(n2434) );
  AOI211XL U419 ( .A0(n2474), .A1(n137), .B0(n2400), .C0(n2402), .Y(n2469) );
  OR2X2 U420 ( .A(n96), .B(n824), .Y(n123) );
  OR2X2 U421 ( .A(n224), .B(n851), .Y(n124) );
  OR2X2 U422 ( .A(n297), .B(n853), .Y(n127) );
  OR2X2 U423 ( .A(n229), .B(n854), .Y(n128) );
  INVXL U424 ( .A(n352), .Y(n296) );
  INVXL U425 ( .A(n354), .Y(n362) );
  INVXL U426 ( .A(n713), .Y(n244) );
  OAI2BB1X2 U427 ( .A0N(N845), .A1N(n232), .B0(n626), .Y(n2946) );
  NOR2XL U428 ( .A(n187), .B(n624), .Y(n625) );
  OAI2BB1X2 U429 ( .A0N(N842), .A1N(n243), .B0(n638), .Y(n2949) );
  NAND2XL U430 ( .A(n381), .B(n1490), .Y(n709) );
  NAND2XL U431 ( .A(n1489), .B(n1490), .Y(n388) );
  INVXL U432 ( .A(n184), .Y(n197) );
  INVXL U433 ( .A(n184), .Y(n196) );
  INVXL U434 ( .A(n1455), .Y(n282) );
  AOI222XL U435 ( .A0(n2381), .A1(n2212), .B0(n2363), .B1(n2382), .C0(n2383), 
        .C1(n370), .Y(n2375) );
  NAND2XL U436 ( .A(n131), .B(n2455), .Y(n2261) );
  AOI21XL U437 ( .A0(n209), .A1(n166), .B0(n267), .Y(n658) );
  AOI21XL U438 ( .A0(n209), .A1(n167), .B0(n267), .Y(n661) );
  AOI21XL U439 ( .A0(n209), .A1(n168), .B0(n272), .Y(n664) );
  AOI21XL U440 ( .A0(n209), .A1(n162), .B0(n267), .Y(n648) );
  AOI21XL U441 ( .A0(n209), .A1(n145), .B0(n272), .Y(n479) );
  NAND2X2 U442 ( .A(N966), .B(n241), .Y(n478) );
  AOI21XL U443 ( .A0(next_A[31]), .A1(n350), .B0(n610), .Y(n611) );
  AOI21XL U444 ( .A0(next_E[31]), .A1(n346), .B0(n548), .Y(n549) );
  AOI21XL U445 ( .A0(n209), .A1(n153), .B0(n267), .Y(n614) );
  NAND2XL U446 ( .A(n344), .B(next_A[30]), .Y(n613) );
  AOI21XL U447 ( .A0(n210), .A1(n155), .B0(n267), .Y(n622) );
  AOI21XL U448 ( .A0(n209), .A1(n154), .B0(n267), .Y(n617) );
  AOI21XL U449 ( .A0(n157), .A1(n207), .B0(n267), .Y(n630) );
  OAI2BB1X2 U450 ( .A0N(N970), .A1N(n242), .B0(n471), .Y(n2788) );
  NOR2XL U451 ( .A(n187), .B(n460), .Y(n461) );
  AOI21XL U452 ( .A0(n208), .A1(n146), .B0(n272), .Y(n485) );
  INVXL U453 ( .A(next_E[10]), .Y(n507) );
  AOI21XL U454 ( .A0(n210), .A1(n172), .B0(n672), .Y(n675) );
  AOI21XL U455 ( .A0(n209), .A1(n165), .B0(n267), .Y(n655) );
  AOI21XL U456 ( .A0(n208), .A1(n148), .B0(n496), .Y(n497) );
  AOI22XL U457 ( .A0(next_E[12]), .A1(n353), .B0(N959), .B1(n243), .Y(n498) );
  NOR2XL U458 ( .A(n187), .B(n464), .Y(n465) );
  NAND2XL U459 ( .A(N956), .B(n239), .Y(n511) );
  AOI21XL U460 ( .A0(n150), .A1(n208), .B0(n272), .Y(n510) );
  INVXL U461 ( .A(next_E[8]), .Y(n517) );
  NAND2XL U462 ( .A(N955), .B(n239), .Y(n515) );
  OR2XL U463 ( .A(n1848), .B(n376), .Y(n129) );
  AOI21XL U464 ( .A0(N1066), .A1(n234), .B0(n268), .Y(n1465) );
  AOI21XL U465 ( .A0(N1065), .A1(n231), .B0(n268), .Y(n1466) );
  AOI21XL U466 ( .A0(N1064), .A1(n241), .B0(n268), .Y(n1467) );
  AOI21XL U467 ( .A0(N1053), .A1(n11), .B0(n268), .Y(n1478) );
  AOI21XL U468 ( .A0(N869), .A1(n240), .B0(n272), .Y(n1767) );
  AOI21XL U469 ( .A0(N868), .A1(n232), .B0(n272), .Y(n1768) );
  AOI21XL U470 ( .A0(N866), .A1(n713), .B0(n272), .Y(n1770) );
  AOI21XL U471 ( .A0(N901), .A1(n233), .B0(n271), .Y(n1735) );
  AOI21XL U472 ( .A0(N900), .A1(n235), .B0(n271), .Y(n1736) );
  AOI21XL U473 ( .A0(N902), .A1(n236), .B0(n271), .Y(n1734) );
  AOI21XL U474 ( .A0(N1034), .A1(n239), .B0(n269), .Y(n1500) );
  AOI21XL U475 ( .A0(N898), .A1(n233), .B0(n271), .Y(n1738) );
  AOI21XL U476 ( .A0(N1025), .A1(n234), .B0(n266), .Y(n1509) );
  AOI21XL U477 ( .A0(N1019), .A1(n235), .B0(n272), .Y(n1515) );
  AOI21XL U478 ( .A0(N1022), .A1(n233), .B0(n272), .Y(n1512) );
  AOI21XL U479 ( .A0(N867), .A1(n232), .B0(n272), .Y(n1769) );
  AOI21XL U480 ( .A0(N862), .A1(n232), .B0(n272), .Y(n1774) );
  AOI21XL U481 ( .A0(N861), .A1(n233), .B0(n268), .Y(n1775) );
  AOI21XL U482 ( .A0(N858), .A1(n713), .B0(n272), .Y(n1778) );
  AOI21XL U483 ( .A0(N1018), .A1(n231), .B0(n266), .Y(n1516) );
  AOI21XL U484 ( .A0(N1027), .A1(n232), .B0(n266), .Y(n1507) );
  AOI21XL U485 ( .A0(N1028), .A1(n232), .B0(n266), .Y(n1506) );
  AOI21XL U486 ( .A0(N1023), .A1(n238), .B0(n272), .Y(n1511) );
  AOI22XL U487 ( .A0(N874), .A1(n243), .B0(n159), .B1(n345), .Y(n1762) );
  AOI22XL U488 ( .A0(N998), .A1(n238), .B0(n145), .B1(n343), .Y(n1621) );
  AOI22XL U489 ( .A0(N994), .A1(n235), .B0(n147), .B1(n340), .Y(n1625) );
  AOI22XL U490 ( .A0(N991), .A1(n237), .B0(n148), .B1(n341), .Y(n1628) );
  AOI22XL U491 ( .A0(N989), .A1(n241), .B0(n149), .B1(n340), .Y(n1630) );
  AOI22XL U492 ( .A0(N988), .A1(n234), .B0(n150), .B1(n351), .Y(n1631) );
  AOI22XL U493 ( .A0(N987), .A1(n240), .B0(n151), .B1(n290), .Y(n1632) );
  AOI22XL U494 ( .A0(N870), .A1(n242), .B0(n162), .B1(n282), .Y(n1766) );
  AOI22XL U495 ( .A0(N985), .A1(n11), .B0(n152), .B1(n345), .Y(n1634) );
  AOI22XL U496 ( .A0(N855), .A1(n243), .B0(n177), .B1(n281), .Y(n1781) );
  AOI22XL U497 ( .A0(N852), .A1(n240), .B0(n60), .B1(n280), .Y(n1784) );
  AOI22XL U498 ( .A0(N856), .A1(n239), .B0(n176), .B1(n347), .Y(n1780) );
  AOI22XL U499 ( .A0(N854), .A1(n231), .B0(n178), .B1(n284), .Y(n1782) );
  INVXL U500 ( .A(next_E[6]), .Y(n525) );
  NAND2XL U501 ( .A(N953), .B(n241), .Y(n524) );
  AOI21XL U502 ( .A0(n152), .A1(n208), .B0(n271), .Y(n523) );
  INVXL U503 ( .A(next_A[6]), .Y(n686) );
  AOI21XL U504 ( .A0(n210), .A1(n175), .B0(n269), .Y(n684) );
  AOI21XL U505 ( .A0(n176), .A1(n207), .B0(n271), .Y(n688) );
  AOI21XL U506 ( .A0(n179), .A1(n207), .B0(n272), .Y(n702) );
  INVXL U507 ( .A(next_A[1]), .Y(n708) );
  NAND2XL U508 ( .A(N820), .B(n713), .Y(n707) );
  AOI21XL U509 ( .A0(n60), .A1(n207), .B0(n267), .Y(n706) );
  INVXL U510 ( .A(next_A[4]), .Y(n695) );
  AOI2BB2XL U511 ( .B0(N918), .B1(n232), .A0N(n308), .A1N(n555), .Y(n550) );
  AOI2BB2XL U512 ( .B0(N916), .B1(n240), .A0N(n291), .A1N(n122), .Y(n552) );
  AOI2BB2XL U513 ( .B0(N873), .B1(n234), .A0N(n278), .A1N(n640), .Y(n572) );
  AOI2BB2XL U514 ( .B0(N853), .B1(n235), .A0N(n309), .A1N(n701), .Y(n574) );
  AOI21XL U515 ( .A0(N819), .A1(n236), .B0(n269), .Y(n711) );
  AOI22XL U516 ( .A0(next_A[0]), .A1(n287), .B0(n59), .B1(n207), .Y(n712) );
  INVX1 U517 ( .A(n368), .Y(n367) );
  INVXL U518 ( .A(next_A[3]), .Y(n700) );
  NAND2BXL U519 ( .AN(n710), .B(N1047), .Y(n383) );
  NAND2BXL U520 ( .AN(n710), .B(N1046), .Y(n386) );
  NAND2BXL U521 ( .AN(n710), .B(N1043), .Y(n390) );
  INVX1 U522 ( .A(n142), .Y(n264) );
  AOI222XL U523 ( .A0(n2353), .A1(n1396), .B0(n2262), .B1(n132), .C0(n2354), 
        .C1(n370), .Y(n2347) );
  AOI31XL U524 ( .A0(n777), .A1(n373), .A2(n2303), .B0(n1877), .Y(n2288) );
  AOI22XL U525 ( .A0(n2279), .A1(n130), .B0(n2215), .B1(n2225), .Y(n2281) );
  AOI211XL U526 ( .A0(n2419), .A1(n370), .B0(n2450), .C0(n2491), .Y(n2488) );
  AOI22XL U527 ( .A0(n137), .A1(n2329), .B0(n2440), .B1(n182), .Y(n2482) );
  AOI222XL U528 ( .A0(n2433), .A1(n370), .B0(n2264), .B1(n28), .C0(n2253), 
        .C1(n130), .Y(n2465) );
  AOI222XL U529 ( .A0(n2267), .A1(round[2]), .B0(n2262), .B1(n370), .C0(n2266), 
        .C1(n743), .Y(n2459) );
  AOI211XL U530 ( .A0(n2345), .A1(n137), .B0(n2360), .C0(n2425), .Y(n2421) );
  AOI222XL U531 ( .A0(n2298), .A1(n132), .B0(n2401), .B1(n131), .C0(n2392), 
        .C1(n28), .Y(n2394) );
  AOI222XL U532 ( .A0(n778), .A1(n182), .B0(n2392), .B1(n370), .C0(n2324), 
        .C1(n181), .Y(n2384) );
  AOI222XL U533 ( .A0(n2381), .A1(n367), .B0(n2364), .B1(n130), .C0(n2391), 
        .C1(n2345), .Y(n2385) );
  NOR2X1 U534 ( .A(n182), .B(n372), .Y(n130) );
  NOR2XL U535 ( .A(n367), .B(n365), .Y(n2212) );
  OAI32XL U536 ( .A0(n777), .A1(n372), .A2(n793), .B0(round[2]), .B1(n2321), 
        .Y(n2320) );
  AOI31XL U537 ( .A0(n791), .A1(n749), .A2(n758), .B0(n370), .Y(n2417) );
  AOI21XL U538 ( .A0(round[2]), .A1(n131), .B0(n2201), .Y(n2195) );
  AOI31XL U539 ( .A0(n181), .A1(round[2]), .A2(n131), .B0(n2481), .Y(n2480) );
  NOR2X1 U540 ( .A(n369), .B(n181), .Y(n132) );
  NOR2XL U541 ( .A(n365), .B(n793), .Y(n2264) );
  AOI21XL U542 ( .A0(n788), .A1(n2250), .B0(n367), .Y(n2380) );
  NAND2XL U543 ( .A(n137), .B(n181), .Y(n2223) );
  NOR2XL U544 ( .A(n367), .B(n181), .Y(n2345) );
  OAI2BB1X4 U545 ( .A0N(n375), .A1N(n374), .B0(n1433), .Y(n1848) );
  BUFX12 U546 ( .A(SHA256_result[108]), .Y(n148) );
  OAI211XL U547 ( .A0(n355), .A1(n963), .B0(n54), .C0(n1447), .Y(n2513) );
  NAND2XL U548 ( .A(H7[11]), .B(n257), .Y(n1447) );
  OAI211XL U549 ( .A0(n355), .A1(n962), .B0(n53), .C0(n1448), .Y(n2514) );
  NAND2XL U550 ( .A(H7[10]), .B(n256), .Y(n1448) );
  OAI211XL U551 ( .A0(n355), .A1(n960), .B0(n49), .C0(n1449), .Y(n2516) );
  NAND2XL U552 ( .A(H7[8]), .B(n257), .Y(n1449) );
  OAI211XL U553 ( .A0(n355), .A1(n956), .B0(n54), .C0(n1450), .Y(n2520) );
  NAND2XL U554 ( .A(H7[4]), .B(n257), .Y(n1450) );
  OAI211XL U555 ( .A0(n355), .A1(n955), .B0(n55), .C0(n1451), .Y(n2521) );
  NAND2XL U556 ( .A(H6[11]), .B(n255), .Y(n1534) );
  OAI211XL U557 ( .A0(n356), .A1(n927), .B0(n52), .C0(n1535), .Y(n2611) );
  NAND2XL U558 ( .A(H6[8]), .B(n255), .Y(n1535) );
  OAI211XL U559 ( .A0(n356), .A1(n926), .B0(n53), .C0(n1536), .Y(n2612) );
  NAND2XL U560 ( .A(H6[7]), .B(n254), .Y(n1536) );
  OAI211XL U561 ( .A0(n359), .A1(n905), .B0(n49), .C0(n1605), .Y(n2736) );
  NAND2XL U562 ( .A(H5[11]), .B(n257), .Y(n1605) );
  OAI211XL U563 ( .A0(n359), .A1(n901), .B0(n48), .C0(n1606), .Y(n2740) );
  NAND2XL U564 ( .A(H5[7]), .B(n255), .Y(n1606) );
  INVXL U565 ( .A(n148), .Y(n886) );
  OAI211XL U566 ( .A0(n358), .A1(n865), .B0(n51), .C0(n1574), .Y(n2673) );
  OAI211XL U567 ( .A0(n358), .A1(n863), .B0(n55), .C0(n1575), .Y(n2675) );
  OAI211XL U568 ( .A0(n358), .A1(n860), .B0(n53), .C0(n1576), .Y(n2678) );
  OAI211XL U569 ( .A0(n358), .A1(n859), .B0(n51), .C0(n1577), .Y(n2679) );
  OAI211XL U570 ( .A0(n358), .A1(n858), .B0(n53), .C0(n1578), .Y(n2680) );
  NAND2XL U571 ( .A(H3[3]), .B(n256), .Y(n1578) );
  NAND2XL U572 ( .A(H3[1]), .B(n254), .Y(n1579) );
  OAI211XL U573 ( .A0(n357), .A1(n831), .B0(n48), .C0(n1555), .Y(n2643) );
  OAI211XL U574 ( .A0(n357), .A1(n830), .B0(n49), .C0(n1556), .Y(n2644) );
  OAI211XL U575 ( .A0(n357), .A1(n828), .B0(n50), .C0(n1557), .Y(n2646) );
  OAI211XL U576 ( .A0(n357), .A1(n827), .B0(n51), .C0(n1558), .Y(n2647) );
  OAI211XL U577 ( .A0(n357), .A1(n826), .B0(n52), .C0(n1559), .Y(n2648) );
  NAND2XL U578 ( .A(H2[1]), .B(n252), .Y(n1560) );
  OAI211XL U579 ( .A0(n355), .A1(n806), .B0(n52), .C0(n1799), .Y(n2929) );
  NAND2XL U580 ( .A(H1[11]), .B(n249), .Y(n1799) );
  OAI211XL U581 ( .A0(n360), .A1(n805), .B0(n55), .C0(n1800), .Y(n2930) );
  OAI211XL U582 ( .A0(n355), .A1(n804), .B0(n55), .C0(n1801), .Y(n2931) );
  NAND2XL U583 ( .A(H1[9]), .B(n249), .Y(n1801) );
  OAI211XL U584 ( .A0(n355), .A1(n802), .B0(n56), .C0(n1802), .Y(n2933) );
  NAND2XL U585 ( .A(H1[7]), .B(n249), .Y(n1802) );
  OAI211XL U586 ( .A0(n355), .A1(n797), .B0(n56), .C0(n1803), .Y(n2938) );
  OAI211XL U587 ( .A0(n355), .A1(n976), .B0(n54), .C0(n1441), .Y(n2500) );
  NAND2XL U588 ( .A(H7[24]), .B(n258), .Y(n1441) );
  OAI211XL U589 ( .A0(n355), .A1(n975), .B0(n55), .C0(n1442), .Y(n2501) );
  NAND2XL U590 ( .A(H7[23]), .B(n258), .Y(n1442) );
  OAI211XL U591 ( .A0(n355), .A1(n974), .B0(n56), .C0(n1443), .Y(n2502) );
  NAND2XL U592 ( .A(H7[22]), .B(n258), .Y(n1443) );
  OAI211XL U593 ( .A0(n355), .A1(n973), .B0(n55), .C0(n1444), .Y(n2503) );
  NAND2XL U594 ( .A(H7[21]), .B(n258), .Y(n1444) );
  OAI211XL U595 ( .A0(n355), .A1(n436), .B0(n54), .C0(n1537), .Y(n2614) );
  AOI21XL U596 ( .A0(n208), .A1(SHA256_result[114]), .B0(n267), .Y(n482) );
  AOI21XL U597 ( .A0(SHA256_result[124]), .A1(n208), .B0(n267), .Y(n454) );
  BUFX8 U598 ( .A(SHA256_result[227]), .Y(n178) );
  NAND2XL U599 ( .A(H2[2]), .B(n256), .Y(n558) );
  NAND2XL U600 ( .A(H2[0]), .B(n256), .Y(n565) );
  INVXL U601 ( .A(n177), .Y(n692) );
  INVXL U602 ( .A(n178), .Y(n697) );
  NAND2XL U603 ( .A(H5[4]), .B(n253), .Y(n419) );
  NAND2XL U604 ( .A(H5[1]), .B(n254), .Y(n426) );
  INVXL U605 ( .A(n149), .Y(n504) );
  INVXL U606 ( .A(n151), .Y(n514) );
  NAND2XL U607 ( .A(H2[3]), .B(n255), .Y(n554) );
  AOI22XL U608 ( .A0(N1008), .A1(n235), .B0(n14), .B1(n353), .Y(n1611) );
  NAND2XL U609 ( .A(H6[3]), .B(n254), .Y(n1538) );
  NAND2XL U610 ( .A(H6[1]), .B(n254), .Y(n1539) );
  OAI211XL U611 ( .A0(n361), .A1(n87), .B0(n52), .C0(n1540), .Y(n2619) );
  NAND2XL U612 ( .A(H6[0]), .B(n254), .Y(n1540) );
  NAND2XL U613 ( .A(H5[3]), .B(n256), .Y(n1607) );
  NAND2XL U614 ( .A(H5[2]), .B(n250), .Y(n1608) );
  OAI211XL U615 ( .A0(n361), .A1(n451), .B0(n53), .C0(n1581), .Y(n2687) );
  OAI211XL U616 ( .A0(n361), .A1(n526), .B0(n54), .C0(n1590), .Y(n2710) );
  OAI211XL U617 ( .A0(n361), .A1(n80), .B0(n44), .C0(n1591), .Y(n2711) );
  NAND3XL U618 ( .A(n133), .B(n53), .C(n1580), .Y(n2685) );
  OR2XL U619 ( .A(n355), .B(n434), .Y(n133) );
  NAND3BXL U620 ( .AN(n509), .B(n53), .C(n1588), .Y(n2706) );
  INVXL U621 ( .A(n150), .Y(n508) );
  NAND3XL U622 ( .A(n134), .B(n52), .C(n1589), .Y(n2709) );
  OR2XL U623 ( .A(n355), .B(n522), .Y(n134) );
  NAND3XL U624 ( .A(n135), .B(n56), .C(n1872), .Y(n2999) );
  OR2XL U625 ( .A(n355), .B(n687), .Y(n135) );
  NAND3BXL U626 ( .AN(n705), .B(n54), .C(n1874), .Y(n3003) );
  OAI2BB2XL U627 ( .B0(n364), .B1(n961), .A0N(H7[9]), .A1N(n260), .Y(n2515) );
  OAI2BB2XL U628 ( .B0(n364), .B1(n959), .A0N(H7[7]), .A1N(n260), .Y(n2517) );
  OAI2BB2XL U629 ( .B0(n364), .B1(n958), .A0N(H7[6]), .A1N(n260), .Y(n2518) );
  OAI2BB2XL U630 ( .B0(n364), .B1(n957), .A0N(H7[5]), .A1N(n260), .Y(n2519) );
  OAI2BB2XL U631 ( .B0(n364), .B1(n929), .A0N(H6[10]), .A1N(n261), .Y(n2609)
         );
  OAI2BB2XL U632 ( .B0(n364), .B1(n928), .A0N(H6[9]), .A1N(n261), .Y(n2610) );
  OAI2BB2XL U633 ( .B0(n364), .B1(n925), .A0N(H6[6]), .A1N(n253), .Y(n2613) );
  OAI2BB2XL U634 ( .B0(n364), .B1(n904), .A0N(H5[10]), .A1N(n259), .Y(n2737)
         );
  OAI2BB2XL U635 ( .B0(n364), .B1(n903), .A0N(H5[9]), .A1N(n259), .Y(n2738) );
  OAI2BB2XL U636 ( .B0(n364), .B1(n902), .A0N(H5[8]), .A1N(n259), .Y(n2739) );
  OAI2BB2XL U637 ( .B0(n364), .B1(n900), .A0N(H5[6]), .A1N(n248), .Y(n2741) );
  INVXL U638 ( .A(n147), .Y(n889) );
  OAI2BB2XL U639 ( .B0(n364), .B1(n866), .A0N(H3[11]), .A1N(n259), .Y(n2672)
         );
  OAI2BB2XL U640 ( .B0(n364), .B1(n864), .A0N(H3[9]), .A1N(n261), .Y(n2674) );
  OAI2BB2XL U641 ( .B0(n364), .B1(n862), .A0N(H3[7]), .A1N(n261), .Y(n2676) );
  OAI2BB2XL U642 ( .B0(n364), .B1(n833), .A0N(H2[11]), .A1N(n259), .Y(n2641)
         );
  OAI2BB2XL U643 ( .B0(n364), .B1(n832), .A0N(H2[10]), .A1N(n261), .Y(n2642)
         );
  OAI2BB2XL U644 ( .B0(n364), .B1(n829), .A0N(H2[7]), .A1N(n260), .Y(n2645) );
  OAI2BB2XL U645 ( .B0(n364), .B1(n803), .A0N(H1[8]), .A1N(n249), .Y(n2932) );
  OAI2BB2XL U646 ( .B0(n364), .B1(n801), .A0N(H1[6]), .A1N(n257), .Y(n2934) );
  OAI2BB2XL U647 ( .B0(n364), .B1(n799), .A0N(H1[4]), .A1N(n251), .Y(n2936) );
  OAI2BB2XL U648 ( .B0(n364), .B1(n726), .A0N(H0[17]), .A1N(n255), .Y(n2987)
         );
  OAI2BB2XL U649 ( .B0(n364), .B1(n720), .A0N(H0[11]), .A1N(n254), .Y(n2993)
         );
  OAI2BB2XL U650 ( .B0(n364), .B1(n717), .A0N(H0[8]), .A1N(n251), .Y(n2996) );
  INVXL U651 ( .A(next_E[16]), .Y(n487) );
  AOI21XL U652 ( .A0(n208), .A1(SHA256_result[120]), .B0(n272), .Y(n469) );
  AOI2BB2XL U653 ( .B0(n189), .B1(SHA256_result[109]), .A0N(n316), .A1N(n494), 
        .Y(n495) );
  CLKBUFX8 U654 ( .A(SHA256_result[249]), .Y(n157) );
  CLKBUFX8 U655 ( .A(SHA256_result[240]), .Y(n165) );
  CLKBUFX8 U656 ( .A(SHA256_result[239]), .Y(n166) );
  CLKBUFX8 U657 ( .A(SHA256_result[251]), .Y(n155) );
  CLKBUFX8 U658 ( .A(SHA256_result[253]), .Y(n154) );
  NAND2XL U659 ( .A(H6[4]), .B(n253), .Y(n394) );
  NAND2XL U660 ( .A(H5[5]), .B(n253), .Y(n416) );
  NAND2XL U661 ( .A(H6[2]), .B(n253), .Y(n399) );
  AOI21XL U662 ( .A0(n210), .A1(SHA256_result[91]), .B0(n266), .Y(n409) );
  AOI22XL U663 ( .A0(N1020), .A1(n231), .B0(SHA256_result[73]), .B1(n285), .Y(
        n1514) );
  AOI22XL U664 ( .A0(N1001), .A1(n235), .B0(SHA256_result[118]), .B1(n349), 
        .Y(n1618) );
  AOI22XL U665 ( .A0(N894), .A1(n713), .B0(SHA256_result[203]), .B1(n348), .Y(
        n1742) );
  AOI22XL U666 ( .A0(N893), .A1(n713), .B0(SHA256_result[202]), .B1(n288), .Y(
        n1743) );
  AOI22XL U667 ( .A0(N890), .A1(n236), .B0(SHA256_result[199]), .B1(n343), .Y(
        n1746) );
  AOI22XL U668 ( .A0(N926), .A1(n243), .B0(SHA256_result[171]), .B1(n285), .Y(
        n1710) );
  AOI22XL U669 ( .A0(N922), .A1(n242), .B0(SHA256_result[167]), .B1(n344), .Y(
        n1714) );
  AOI22XL U670 ( .A0(N915), .A1(n240), .B0(n72), .B1(n347), .Y(n1721) );
  AOI22XL U671 ( .A0(N899), .A1(n11), .B0(SHA256_result[208]), .B1(n352), .Y(
        n1737) );
  AOI22XL U672 ( .A0(N924), .A1(n240), .B0(SHA256_result[169]), .B1(n350), .Y(
        n1712) );
  AOI22XL U673 ( .A0(N921), .A1(n241), .B0(SHA256_result[166]), .B1(n286), .Y(
        n1715) );
  AOI22XL U674 ( .A0(N1002), .A1(n713), .B0(SHA256_result[119]), .B1(n290), 
        .Y(n1617) );
  AOI22XL U675 ( .A0(N1033), .A1(n233), .B0(SHA256_result[86]), .B1(n346), .Y(
        n1501) );
  AOI22XL U676 ( .A0(N1030), .A1(n239), .B0(SHA256_result[83]), .B1(n289), .Y(
        n1504) );
  AOI22XL U677 ( .A0(N1029), .A1(n242), .B0(SHA256_result[82]), .B1(n281), .Y(
        n1505) );
  AOI22XL U678 ( .A0(N1024), .A1(n234), .B0(SHA256_result[77]), .B1(n346), .Y(
        n1510) );
  AOI21XL U679 ( .A0(n85), .A1(n208), .B0(n266), .Y(n402) );
  AOI22XL U680 ( .A0(N1045), .A1(n243), .B0(SHA256_result[34]), .B1(n288), .Y(
        n1486) );
  AOI22XL U681 ( .A0(N1044), .A1(n235), .B0(n85), .B1(n284), .Y(n1487) );
  AOI22XL U682 ( .A0(N1048), .A1(n236), .B0(SHA256_result[37]), .B1(n352), .Y(
        n1483) );
  AOI22XL U683 ( .A0(N1060), .A1(n235), .B0(SHA256_result[49]), .B1(n349), .Y(
        n1471) );
  AOI22XL U684 ( .A0(N1059), .A1(n242), .B0(SHA256_result[48]), .B1(n353), .Y(
        n1472) );
  AOI22XL U685 ( .A0(N1050), .A1(n238), .B0(SHA256_result[39]), .B1(n284), .Y(
        n1481) );
  AOI22XL U686 ( .A0(N1063), .A1(n239), .B0(SHA256_result[52]), .B1(n352), .Y(
        n1468) );
  AOI22XL U687 ( .A0(N1056), .A1(n713), .B0(n12), .B1(n283), .Y(n1475) );
  AOI22XL U688 ( .A0(N1055), .A1(n234), .B0(SHA256_result[44]), .B1(n347), .Y(
        n1476) );
  AOI22XL U689 ( .A0(N1062), .A1(n236), .B0(SHA256_result[51]), .B1(n348), .Y(
        n1469) );
  AOI22XL U690 ( .A0(N1061), .A1(n231), .B0(SHA256_result[50]), .B1(n345), .Y(
        n1470) );
  AOI22XL U691 ( .A0(N1049), .A1(n241), .B0(SHA256_result[38]), .B1(n352), .Y(
        n1482) );
  AOI22XL U692 ( .A0(N1052), .A1(n238), .B0(SHA256_result[41]), .B1(n342), .Y(
        n1479) );
  NAND2XL U693 ( .A(n86), .B(n191), .Y(n431) );
  AOI21XL U694 ( .A0(SHA256_result[37]), .A1(n208), .B0(n266), .Y(n392) );
  INVXL U695 ( .A(next_E[7]), .Y(n521) );
  INVXL U696 ( .A(next_E[3]), .Y(n536) );
  INVXL U697 ( .A(next_E[2]), .Y(n539) );
  INVXL U698 ( .A(next_E[1]), .Y(n542) );
  INVXL U699 ( .A(next_E[5]), .Y(n529) );
  AOI21XL U700 ( .A0(SHA256_result[101]), .A1(n207), .B0(n272), .Y(n527) );
  INVXL U701 ( .A(next_E[4]), .Y(n532) );
  AOI21XL U702 ( .A0(n43), .A1(n207), .B0(n272), .Y(n530) );
  AOI21XL U703 ( .A0(n15), .A1(n207), .B0(n267), .Y(n543) );
  AOI21XL U704 ( .A0(SHA256_result[35]), .A1(n207), .B0(n266), .Y(n397) );
  OAI211XL U705 ( .A0(n296), .A1(n443), .B0(n405), .C0(n404), .Y(n2620) );
  AOI21XL U706 ( .A0(n89), .A1(n208), .B0(n266), .Y(n404) );
  AOI21XL U707 ( .A0(SHA256_result[67]), .A1(n208), .B0(n266), .Y(n422) );
  AOI21XL U708 ( .A0(SHA256_result[66]), .A1(n208), .B0(n266), .Y(n424) );
  NAND2XL U709 ( .A(SHA256_result[69]), .B(n193), .Y(n418) );
  NAND2XL U710 ( .A(n66), .B(n191), .Y(n428) );
  NAND2XL U711 ( .A(n72), .B(n197), .Y(n564) );
  NAND2XL U712 ( .A(SHA256_result[36]), .B(n194), .Y(n396) );
  NAND2XL U713 ( .A(N1015), .B(n243), .Y(n395) );
  NAND2XL U714 ( .A(N884), .B(n233), .Y(n562) );
  AOI21XL U715 ( .A0(n121), .A1(n207), .B0(n267), .Y(n561) );
  NAND2XL U716 ( .A(N990), .B(n713), .Y(n413) );
  AOI21XL U717 ( .A0(n209), .A1(SHA256_result[75]), .B0(n266), .Y(n412) );
  NAND2XL U718 ( .A(N986), .B(n240), .Y(n415) );
  AOI21XL U719 ( .A0(n209), .A1(SHA256_result[71]), .B0(n266), .Y(n414) );
  NAND2XL U720 ( .A(SHA256_result[68]), .B(n192), .Y(n421) );
  NAND2XL U721 ( .A(N983), .B(n11), .Y(n420) );
  NAND2XL U722 ( .A(SHA256_result[163]), .B(n194), .Y(n557) );
  NAND2XL U723 ( .A(N886), .B(n235), .Y(n556) );
  NAND2XL U724 ( .A(n94), .B(n196), .Y(n560) );
  NAND2XL U725 ( .A(N885), .B(n240), .Y(n559) );
  AOI2BB2XL U726 ( .B0(N851), .B1(n235), .A0N(n298), .A1N(n98), .Y(n576) );
  NOR3XL U727 ( .A(output_enable), .B(round[6]), .C(n1848), .Y(n141) );
  AOI222XL U728 ( .A0(n2362), .A1(n367), .B0(n2363), .B1(n370), .C0(n2364), 
        .C1(n1396), .Y(n2355) );
  AOI31XL U729 ( .A0(n182), .A1(n1388), .A2(n2311), .B0(n2361), .Y(n2356) );
  AOI22XL U730 ( .A0(n2214), .A1(n367), .B0(n2336), .B1(n1370), .Y(n2330) );
  AOI221XL U731 ( .A0(n757), .A1(n1383), .B0(n2262), .B1(n181), .C0(n2263), 
        .Y(n2256) );
  AOI2BB2XL U732 ( .B0(n2254), .B1(round[2]), .A0N(n2243), .A1N(n1396), .Y(
        n2244) );
  AOI31XL U733 ( .A0(n2303), .A1(n370), .A2(n2215), .B0(n2267), .Y(n2476) );
  NOR3XL U734 ( .A(n2450), .B(n2225), .C(n2267), .Y(n2442) );
  AOI211XL U735 ( .A0(n2379), .A1(n370), .B0(n2416), .C0(n2417), .Y(n2415) );
  AND3X1 U736 ( .A(n1433), .B(n380), .C(inner_busy), .Y(n142) );
  NAND2XL U737 ( .A(output_enable), .B(n1433), .Y(n136) );
  NOR3XL U738 ( .A(n1370), .B(round[2]), .C(n139), .Y(n2400) );
  NOR3XL U739 ( .A(n777), .B(n1383), .C(n367), .Y(n2311) );
  NOR3XL U740 ( .A(n1383), .B(n181), .C(n752), .Y(n2217) );
  INVX1 U741 ( .A(n366), .Y(n365) );
  OAI22XL U742 ( .A0(round[3]), .A1(n2258), .B0(n2472), .B1(n1370), .Y(n2471)
         );
  NOR2XL U743 ( .A(n1388), .B(round[3]), .Y(n2216) );
  NOR2XL U744 ( .A(n1370), .B(round[3]), .Y(n2283) );
  AOI222XL U745 ( .A0(n2427), .A1(n1383), .B0(n2379), .B1(n1370), .C0(n2383), 
        .C1(n181), .Y(n2467) );
  AOI22XL U746 ( .A0(n29), .A1(SHA256_result[0]), .B0(n2022), .B1(
        SHA256_result[8]), .Y(n2189) );
  AOI22XL U747 ( .A0(n29), .A1(SHA256_result[1]), .B0(n2022), .B1(
        SHA256_result[9]), .Y(n2154) );
  AOI22XL U748 ( .A0(n29), .A1(SHA256_result[2]), .B0(n2022), .B1(
        SHA256_result[10]), .Y(n2133) );
  AOI22XL U749 ( .A0(n29), .A1(SHA256_result[3]), .B0(n2022), .B1(
        SHA256_result[11]), .Y(n2112) );
  AOI22XL U750 ( .A0(n29), .A1(SHA256_result[4]), .B0(n2022), .B1(
        SHA256_result[12]), .Y(n2091) );
  AOI22XL U751 ( .A0(n29), .A1(SHA256_result[5]), .B0(n2022), .B1(
        SHA256_result[13]), .Y(n2070) );
  AOI22XL U752 ( .A0(n29), .A1(SHA256_result[6]), .B0(n2022), .B1(
        SHA256_result[14]), .Y(n2049) );
  AOI22XL U753 ( .A0(n29), .A1(SHA256_result[7]), .B0(n2022), .B1(
        SHA256_result[15]), .Y(n2021) );
  AOI22XL U754 ( .A0(n2002), .A1(n94), .B0(n2003), .B1(SHA256_result[170]), 
        .Y(n2123) );
  AOI22XL U755 ( .A0(n1986), .A1(SHA256_result[199]), .B0(n1987), .B1(
        SHA256_result[207]), .Y(n1985) );
  AOI22XL U756 ( .A0(n1986), .A1(SHA256_result[194]), .B0(n1987), .B1(
        SHA256_result[202]), .Y(n2121) );
  AOI22XL U757 ( .A0(n1986), .A1(SHA256_result[195]), .B0(n1987), .B1(
        SHA256_result[203]), .Y(n2100) );
  AOI22XL U758 ( .A0(n2025), .A1(SHA256_result[39]), .B0(n2026), .B1(
        SHA256_result[47]), .Y(n2019) );
  AOI22XL U759 ( .A0(n2027), .A1(SHA256_result[48]), .B0(n2028), .B1(
        SHA256_result[56]), .Y(n2186) );
  AOI22XL U760 ( .A0(n2027), .A1(SHA256_result[49]), .B0(n2028), .B1(
        SHA256_result[57]), .Y(n2151) );
  AOI22XL U761 ( .A0(n2027), .A1(SHA256_result[50]), .B0(n2028), .B1(
        SHA256_result[58]), .Y(n2130) );
  AOI22XL U762 ( .A0(n2027), .A1(SHA256_result[51]), .B0(n2028), .B1(
        SHA256_result[59]), .Y(n2109) );
  AOI22XL U763 ( .A0(n2027), .A1(SHA256_result[52]), .B0(n2028), .B1(
        SHA256_result[60]), .Y(n2088) );
  AOI22XL U764 ( .A0(n2002), .A1(n121), .B0(n2003), .B1(SHA256_result[169]), 
        .Y(n2144) );
  AOI22XL U765 ( .A0(n2025), .A1(SHA256_result[38]), .B0(n2026), .B1(
        SHA256_result[46]), .Y(n2047) );
  AOI22XL U766 ( .A0(n2002), .A1(SHA256_result[166]), .B0(n2003), .B1(
        SHA256_result[174]), .Y(n2039) );
  AOI22XL U767 ( .A0(n2002), .A1(SHA256_result[167]), .B0(n2003), .B1(
        SHA256_result[175]), .Y(n1995) );
  AOI22XL U768 ( .A0(n2027), .A1(SHA256_result[53]), .B0(n2028), .B1(
        SHA256_result[61]), .Y(n2067) );
  AOI22XL U769 ( .A0(n2002), .A1(SHA256_result[163]), .B0(n2003), .B1(
        SHA256_result[171]), .Y(n2102) );
  AOI22XL U770 ( .A0(n2004), .A1(SHA256_result[177]), .B0(n2005), .B1(
        SHA256_result[185]), .Y(n2143) );
  AOI22XL U771 ( .A0(n2004), .A1(SHA256_result[179]), .B0(n2005), .B1(
        SHA256_result[187]), .Y(n2101) );
  AOI22XL U772 ( .A0(n2027), .A1(SHA256_result[55]), .B0(n2028), .B1(
        SHA256_result[63]), .Y(n2018) );
  AOI22XL U773 ( .A0(n2010), .A1(SHA256_result[71]), .B0(n2011), .B1(
        SHA256_result[79]), .Y(n2009) );
  AOI22XL U774 ( .A0(n2025), .A1(n85), .B0(n2026), .B1(SHA256_result[41]), .Y(
        n2152) );
  AOI22XL U775 ( .A0(n2025), .A1(SHA256_result[36]), .B0(n2026), .B1(
        SHA256_result[44]), .Y(n2089) );
  AOI22XL U776 ( .A0(n2025), .A1(SHA256_result[37]), .B0(n2026), .B1(n12), .Y(
        n2068) );
  AOI22XL U777 ( .A0(n2010), .A1(SHA256_result[70]), .B0(n2011), .B1(
        SHA256_result[78]), .Y(n2045) );
  AOI22XL U778 ( .A0(n2010), .A1(SHA256_result[67]), .B0(n2011), .B1(
        SHA256_result[75]), .Y(n2108) );
  AOI22XL U779 ( .A0(n1986), .A1(SHA256_result[193]), .B0(n1987), .B1(
        SHA256_result[201]), .Y(n2142) );
  AOI22XL U780 ( .A0(n2010), .A1(n66), .B0(n2011), .B1(SHA256_result[73]), .Y(
        n2150) );
  AOI22XL U781 ( .A0(n2010), .A1(SHA256_result[66]), .B0(n2011), .B1(
        SHA256_result[74]), .Y(n2129) );
  AOI22XL U782 ( .A0(n1986), .A1(SHA256_result[196]), .B0(n1987), .B1(
        SHA256_result[204]), .Y(n2079) );
  AOI22XL U783 ( .A0(n1986), .A1(SHA256_result[197]), .B0(n1987), .B1(
        SHA256_result[205]), .Y(n2058) );
  AOI22XL U784 ( .A0(n2010), .A1(SHA256_result[69]), .B0(n2011), .B1(
        SHA256_result[77]), .Y(n2066) );
  AOI22XL U785 ( .A0(n1986), .A1(SHA256_result[198]), .B0(n1987), .B1(
        SHA256_result[206]), .Y(n2037) );
  AOI22XL U786 ( .A0(n2027), .A1(SHA256_result[54]), .B0(n2028), .B1(
        SHA256_result[62]), .Y(n2046) );
  AOI22XL U787 ( .A0(n2004), .A1(SHA256_result[176]), .B0(n2005), .B1(
        SHA256_result[184]), .Y(n2170) );
  AOI22XL U788 ( .A0(n2004), .A1(SHA256_result[178]), .B0(n2005), .B1(
        SHA256_result[186]), .Y(n2122) );
  AOI22XL U789 ( .A0(n1986), .A1(SHA256_result[192]), .B0(n1987), .B1(
        SHA256_result[200]), .Y(n2163) );
  AOI22XL U790 ( .A0(n2002), .A1(SHA256_result[164]), .B0(n2003), .B1(
        SHA256_result[172]), .Y(n2081) );
  AOI22XL U791 ( .A0(n2002), .A1(SHA256_result[165]), .B0(n2003), .B1(
        SHA256_result[173]), .Y(n2060) );
  AOI22XL U792 ( .A0(n2025), .A1(n89), .B0(n2026), .B1(SHA256_result[40]), .Y(
        n2187) );
  AOI22XL U793 ( .A0(n2025), .A1(SHA256_result[34]), .B0(n2026), .B1(
        SHA256_result[42]), .Y(n2131) );
  AOI22XL U794 ( .A0(n2025), .A1(SHA256_result[35]), .B0(n2026), .B1(
        SHA256_result[43]), .Y(n2110) );
  AOI22XL U795 ( .A0(n2002), .A1(n72), .B0(n2003), .B1(SHA256_result[168]), 
        .Y(n2171) );
  AOI22XL U796 ( .A0(n2023), .A1(SHA256_result[16]), .B0(n2024), .B1(
        SHA256_result[24]), .Y(n2188) );
  AOI22XL U797 ( .A0(n2023), .A1(SHA256_result[17]), .B0(n2024), .B1(
        SHA256_result[25]), .Y(n2153) );
  AOI22XL U798 ( .A0(n2023), .A1(SHA256_result[20]), .B0(n2024), .B1(
        SHA256_result[28]), .Y(n2090) );
  AOI22XL U799 ( .A0(n2023), .A1(SHA256_result[21]), .B0(n2024), .B1(
        SHA256_result[29]), .Y(n2069) );
  AOI22XL U800 ( .A0(n2023), .A1(SHA256_result[18]), .B0(n2024), .B1(
        SHA256_result[26]), .Y(n2132) );
  AOI22XL U801 ( .A0(n2023), .A1(SHA256_result[19]), .B0(n2024), .B1(
        SHA256_result[27]), .Y(n2111) );
  AOI22XL U802 ( .A0(n2023), .A1(SHA256_result[22]), .B0(n2024), .B1(
        SHA256_result[30]), .Y(n2048) );
  AOI22XL U803 ( .A0(n2023), .A1(SHA256_result[23]), .B0(n2024), .B1(
        SHA256_result[31]), .Y(n2020) );
  AOI22XL U804 ( .A0(n2010), .A1(SHA256_result[68]), .B0(n2011), .B1(
        SHA256_result[76]), .Y(n2087) );
  AOI22XL U805 ( .A0(n1998), .A1(SHA256_result[128]), .B0(n1999), .B1(
        SHA256_result[136]), .Y(n2173) );
  AOI22XL U806 ( .A0(n1998), .A1(SHA256_result[130]), .B0(n1999), .B1(
        SHA256_result[138]), .Y(n2125) );
  AOI22XL U807 ( .A0(n1998), .A1(SHA256_result[131]), .B0(n1999), .B1(
        SHA256_result[139]), .Y(n2104) );
  AOI22XL U808 ( .A0(n1998), .A1(SHA256_result[129]), .B0(n1999), .B1(
        SHA256_result[137]), .Y(n2146) );
  AOI22XL U809 ( .A0(n2010), .A1(n86), .B0(n2011), .B1(SHA256_result[72]), .Y(
        n2181) );
  AOI22XL U810 ( .A0(n1992), .A1(n161), .B0(n1993), .B1(n13), .Y(n2076) );
  AOI22XL U811 ( .A0(n1990), .A1(n177), .B0(n1991), .B1(n169), .Y(n2077) );
  AOI22XL U812 ( .A0(n2016), .A1(SHA256_result[119]), .B0(n2017), .B1(
        SHA256_result[127]), .Y(n2006) );
  AOI22XL U813 ( .A0(n2012), .A1(SHA256_result[87]), .B0(n2013), .B1(
        SHA256_result[95]), .Y(n2008) );
  AOI22XL U814 ( .A0(n2016), .A1(SHA256_result[114]), .B0(n2017), .B1(
        SHA256_result[122]), .Y(n2126) );
  AOI22XL U815 ( .A0(n2012), .A1(SHA256_result[82]), .B0(n2013), .B1(
        SHA256_result[90]), .Y(n2128) );
  AOI22XL U816 ( .A0(n2016), .A1(n145), .B0(n2017), .B1(SHA256_result[123]), 
        .Y(n2105) );
  AOI22XL U817 ( .A0(n2012), .A1(SHA256_result[83]), .B0(n2013), .B1(
        SHA256_result[91]), .Y(n2107) );
  AOI22XL U818 ( .A0(n2016), .A1(n146), .B0(n2017), .B1(SHA256_result[121]), 
        .Y(n2147) );
  AOI22XL U819 ( .A0(n2012), .A1(SHA256_result[81]), .B0(n2013), .B1(
        SHA256_result[89]), .Y(n2149) );
  AOI22XL U820 ( .A0(n2016), .A1(SHA256_result[118]), .B0(n2017), .B1(n143), 
        .Y(n2042) );
  AOI22XL U821 ( .A0(n2012), .A1(SHA256_result[86]), .B0(n2013), .B1(
        SHA256_result[94]), .Y(n2044) );
  AOI22XL U822 ( .A0(n2014), .A1(n152), .B0(n2015), .B1(SHA256_result[110]), 
        .Y(n2043) );
  AOI22XL U823 ( .A0(n2016), .A1(SHA256_result[112]), .B0(n2017), .B1(
        SHA256_result[120]), .Y(n2178) );
  AOI22XL U824 ( .A0(n2012), .A1(SHA256_result[80]), .B0(n2013), .B1(
        SHA256_result[88]), .Y(n2180) );
  AOI22XL U825 ( .A0(n2014), .A1(n15), .B0(n2015), .B1(n151), .Y(n2179) );
  AOI22XL U826 ( .A0(n2016), .A1(n144), .B0(n2017), .B1(n14), .Y(n2063) );
  AOI22XL U827 ( .A0(n2012), .A1(SHA256_result[85]), .B0(n2013), .B1(
        SHA256_result[93]), .Y(n2065) );
  AOI22XL U828 ( .A0(n2014), .A1(SHA256_result[101]), .B0(n2015), .B1(
        SHA256_result[109]), .Y(n2064) );
  AOI22XL U829 ( .A0(n2016), .A1(SHA256_result[116]), .B0(n2017), .B1(
        SHA256_result[124]), .Y(n2084) );
  AOI22XL U830 ( .A0(n2012), .A1(SHA256_result[84]), .B0(n2013), .B1(
        SHA256_result[92]), .Y(n2086) );
  AOI22XL U831 ( .A0(n2014), .A1(n43), .B0(n2015), .B1(n148), .Y(n2085) );
  AOI22XL U832 ( .A0(n1992), .A1(n163), .B0(n1993), .B1(n156), .Y(n2118) );
  AOI22XL U833 ( .A0(n1988), .A1(SHA256_result[210]), .B0(n1989), .B1(
        SHA256_result[218]), .Y(n2120) );
  AOI22XL U834 ( .A0(n1990), .A1(n179), .B0(n1991), .B1(n171), .Y(n2119) );
  AOI22XL U835 ( .A0(n1992), .A1(n162), .B0(n1993), .B1(n155), .Y(n2097) );
  AOI22XL U836 ( .A0(n1988), .A1(SHA256_result[211]), .B0(n1989), .B1(
        SHA256_result[219]), .Y(n2099) );
  AOI22XL U837 ( .A0(n1990), .A1(n178), .B0(n1991), .B1(n170), .Y(n2098) );
  AOI22XL U838 ( .A0(n1992), .A1(SHA256_result[246]), .B0(n1993), .B1(n153), 
        .Y(n2034) );
  AOI22XL U839 ( .A0(n1990), .A1(n175), .B0(n1991), .B1(n167), .Y(n2035) );
  AOI22XL U840 ( .A0(n1992), .A1(n159), .B0(n1993), .B1(SHA256_result[255]), 
        .Y(n1982) );
  AOI22XL U841 ( .A0(n1990), .A1(n174), .B0(n1991), .B1(n166), .Y(n1983) );
  AOI22XL U842 ( .A0(n1992), .A1(n165), .B0(n1993), .B1(n158), .Y(n2160) );
  AOI22XL U843 ( .A0(n1988), .A1(SHA256_result[208]), .B0(n1989), .B1(
        SHA256_result[216]), .Y(n2162) );
  AOI22XL U844 ( .A0(n1990), .A1(n59), .B0(n1991), .B1(n173), .Y(n2161) );
  AOI22XL U845 ( .A0(n1992), .A1(n164), .B0(n1993), .B1(n157), .Y(n2139) );
  AOI22XL U846 ( .A0(n1988), .A1(SHA256_result[209]), .B0(n1989), .B1(
        SHA256_result[217]), .Y(n2141) );
  AOI22XL U847 ( .A0(n1990), .A1(n60), .B0(n1991), .B1(n172), .Y(n2140) );
  AOI22XL U848 ( .A0(n1992), .A1(n160), .B0(n1993), .B1(n154), .Y(n2055) );
  AOI22XL U849 ( .A0(n1990), .A1(n176), .B0(n1991), .B1(n168), .Y(n2056) );
  INVXL U850 ( .A(n13), .Y(n732) );
  INVXL U851 ( .A(SHA256_result[255]), .Y(n735) );
  INVXL U852 ( .A(SHA256_result[123]), .Y(n456) );
  INVXL U853 ( .A(SHA256_result[246]), .Y(n640) );
  INVXL U854 ( .A(SHA256_result[118]), .Y(n896) );
  INVXL U855 ( .A(SHA256_result[121]), .Y(n464) );
  INVXL U856 ( .A(SHA256_result[127]), .Y(n547) );
  INVXL U857 ( .A(SHA256_result[193]), .Y(n796) );
  INVXL U858 ( .A(SHA256_result[210]), .Y(n813) );
  INVXL U859 ( .A(SHA256_result[209]), .Y(n812) );
  INVXL U860 ( .A(SHA256_result[207]), .Y(n810) );
  INVXL U861 ( .A(SHA256_result[205]), .Y(n808) );
  INVXL U862 ( .A(SHA256_result[201]), .Y(n804) );
  INVXL U863 ( .A(SHA256_result[211]), .Y(n814) );
  INVXL U864 ( .A(SHA256_result[198]), .Y(n801) );
  INVXL U865 ( .A(SHA256_result[197]), .Y(n800) );
  INVXL U866 ( .A(SHA256_result[196]), .Y(n799) );
  INVXL U867 ( .A(SHA256_result[206]), .Y(n809) );
  INVXL U868 ( .A(SHA256_result[204]), .Y(n807) );
  INVXL U869 ( .A(SHA256_result[200]), .Y(n803) );
  INVXL U870 ( .A(SHA256_result[55]), .Y(n942) );
  INVXL U871 ( .A(SHA256_result[80]), .Y(n910) );
  INVXL U872 ( .A(SHA256_result[47]), .Y(n934) );
  INVXL U873 ( .A(SHA256_result[46]), .Y(n933) );
  INVXL U874 ( .A(SHA256_result[43]), .Y(n930) );
  INVXL U875 ( .A(SHA256_result[40]), .Y(n927) );
  INVXL U876 ( .A(SHA256_result[179]), .Y(n841) );
  INVXL U877 ( .A(SHA256_result[178]), .Y(n840) );
  INVXL U878 ( .A(SHA256_result[177]), .Y(n839) );
  INVXL U879 ( .A(SHA256_result[165]), .Y(n827) );
  INVXL U880 ( .A(SHA256_result[164]), .Y(n826) );
  INVXL U881 ( .A(SHA256_result[78]), .Y(n908) );
  INVXL U882 ( .A(SHA256_result[175]), .Y(n837) );
  INVXL U883 ( .A(SHA256_result[174]), .Y(n836) );
  INVXL U884 ( .A(SHA256_result[173]), .Y(n835) );
  INVXL U885 ( .A(SHA256_result[172]), .Y(n834) );
  INVXL U886 ( .A(SHA256_result[168]), .Y(n830) );
  INVXL U887 ( .A(SHA256_result[54]), .Y(n941) );
  INVXL U888 ( .A(SHA256_result[53]), .Y(n940) );
  INVXL U889 ( .A(SHA256_result[87]), .Y(n917) );
  INVXL U890 ( .A(SHA256_result[81]), .Y(n911) );
  INVXL U891 ( .A(SHA256_result[42]), .Y(n929) );
  INVXL U892 ( .A(SHA256_result[176]), .Y(n838) );
  INVXL U893 ( .A(SHA256_result[79]), .Y(n909) );
  INVXL U894 ( .A(SHA256_result[76]), .Y(n906) );
  INVXL U895 ( .A(SHA256_result[72]), .Y(n902) );
  INVXL U896 ( .A(SHA256_result[170]), .Y(n832) );
  INVXL U897 ( .A(SHA256_result[119]), .Y(n897) );
  INVXL U898 ( .A(SHA256_result[120]), .Y(n898) );
  INVXL U899 ( .A(n14), .Y(n448) );
  INVXL U900 ( .A(SHA256_result[208]), .Y(n811) );
  INVXL U901 ( .A(SHA256_result[199]), .Y(n802) );
  INVXL U902 ( .A(SHA256_result[203]), .Y(n806) );
  INVXL U903 ( .A(SHA256_result[202]), .Y(n805) );
  INVXL U904 ( .A(SHA256_result[194]), .Y(n797) );
  INVXL U905 ( .A(SHA256_result[195]), .Y(n798) );
  INVXL U906 ( .A(SHA256_result[71]), .Y(n901) );
  INVXL U907 ( .A(SHA256_result[39]), .Y(n926) );
  INVXL U908 ( .A(SHA256_result[75]), .Y(n905) );
  INVXL U909 ( .A(SHA256_result[49]), .Y(n936) );
  INVXL U910 ( .A(SHA256_result[48]), .Y(n935) );
  INVXL U911 ( .A(SHA256_result[82]), .Y(n912) );
  INVXL U912 ( .A(SHA256_result[166]), .Y(n828) );
  INVXL U913 ( .A(SHA256_result[44]), .Y(n931) );
  INVXL U914 ( .A(SHA256_result[77]), .Y(n907) );
  INVXL U915 ( .A(SHA256_result[169]), .Y(n831) );
  INVXL U916 ( .A(SHA256_result[52]), .Y(n939) );
  INVXL U917 ( .A(SHA256_result[51]), .Y(n938) );
  INVXL U918 ( .A(SHA256_result[50]), .Y(n937) );
  INVXL U919 ( .A(SHA256_result[38]), .Y(n925) );
  INVXL U920 ( .A(SHA256_result[86]), .Y(n916) );
  INVXL U921 ( .A(SHA256_result[85]), .Y(n915) );
  INVXL U922 ( .A(SHA256_result[84]), .Y(n914) );
  INVXL U923 ( .A(SHA256_result[83]), .Y(n913) );
  INVXL U924 ( .A(SHA256_result[70]), .Y(n900) );
  INVXL U925 ( .A(SHA256_result[167]), .Y(n829) );
  INVXL U926 ( .A(n12), .Y(n932) );
  INVXL U927 ( .A(SHA256_result[41]), .Y(n928) );
  INVXL U928 ( .A(SHA256_result[74]), .Y(n904) );
  INVXL U929 ( .A(SHA256_result[73]), .Y(n903) );
  INVXL U930 ( .A(SHA256_result[171]), .Y(n833) );
  INVXL U931 ( .A(SHA256_result[2]), .Y(n954) );
  NOR2XL U932 ( .A(n182), .B(n1383), .Y(n2411) );
  INVXL U933 ( .A(SHA256_result[131]), .Y(n858) );
  INVXL U934 ( .A(SHA256_result[1]), .Y(n953) );
  INVXL U935 ( .A(SHA256_result[21]), .Y(n973) );
  INVXL U936 ( .A(SHA256_result[129]), .Y(n856) );
  INVXL U937 ( .A(SHA256_result[11]), .Y(n963) );
  INVXL U938 ( .A(SHA256_result[23]), .Y(n975) );
  INVXL U939 ( .A(SHA256_result[22]), .Y(n974) );
  INVXL U940 ( .A(SHA256_result[15]), .Y(n967) );
  INVXL U941 ( .A(SHA256_result[14]), .Y(n966) );
  INVXL U942 ( .A(SHA256_result[10]), .Y(n962) );
  INVXL U943 ( .A(SHA256_result[8]), .Y(n960) );
  INVXL U944 ( .A(SHA256_result[5]), .Y(n957) );
  INVXL U945 ( .A(SHA256_result[20]), .Y(n972) );
  INVXL U946 ( .A(SHA256_result[17]), .Y(n969) );
  INVXL U947 ( .A(SHA256_result[16]), .Y(n968) );
  INVXL U948 ( .A(SHA256_result[7]), .Y(n959) );
  INVXL U949 ( .A(SHA256_result[13]), .Y(n965) );
  INVXL U950 ( .A(SHA256_result[12]), .Y(n964) );
  INVXL U951 ( .A(SHA256_result[19]), .Y(n971) );
  INVXL U952 ( .A(SHA256_result[18]), .Y(n970) );
  INVXL U953 ( .A(SHA256_result[6]), .Y(n958) );
  INVXL U954 ( .A(SHA256_result[130]), .Y(n857) );
  INVXL U955 ( .A(SHA256_result[128]), .Y(n855) );
  INVXL U956 ( .A(SHA256_result[9]), .Y(n961) );
  INVXL U957 ( .A(SHA256_result[0]), .Y(n952) );
  INVXL U958 ( .A(SHA256_result[3]), .Y(n955) );
  INVXL U959 ( .A(SHA256_result[4]), .Y(n956) );
  INVXL U960 ( .A(SHA256_result[163]), .Y(n555) );
  INVXL U961 ( .A(SHA256_result[122]), .Y(n460) );
  INVXL U962 ( .A(SHA256_result[101]), .Y(n526) );
  INVXL U963 ( .A(SHA256_result[124]), .Y(n451) );
  INVXL U964 ( .A(SHA256_result[110]), .Y(n888) );
  INVXL U965 ( .A(SHA256_result[112]), .Y(n890) );
  INVXL U966 ( .A(SHA256_result[109]), .Y(n887) );
  INVXL U967 ( .A(SHA256_result[107]), .Y(n500) );
  INVXL U968 ( .A(SHA256_result[192]), .Y(n795) );
  INVX1 U969 ( .A(n213), .Y(n207) );
  INVX1 U970 ( .A(n213), .Y(n208) );
  INVX1 U971 ( .A(n205), .Y(n210) );
  INVX1 U972 ( .A(n349), .Y(n306) );
  INVX1 U973 ( .A(n347), .Y(n305) );
  INVX1 U974 ( .A(n351), .Y(n304) );
  INVX1 U975 ( .A(n350), .Y(n303) );
  INVX1 U976 ( .A(n350), .Y(n302) );
  INVX1 U977 ( .A(n350), .Y(n301) );
  INVX1 U978 ( .A(n350), .Y(n300) );
  INVX1 U979 ( .A(n351), .Y(n297) );
  INVX1 U980 ( .A(n348), .Y(n313) );
  INVX1 U981 ( .A(n348), .Y(n314) );
  INVX1 U982 ( .A(n347), .Y(n318) );
  INVX1 U983 ( .A(n350), .Y(n319) );
  INVX1 U984 ( .A(n351), .Y(n320) );
  INVX1 U985 ( .A(n346), .Y(n322) );
  INVX1 U986 ( .A(n346), .Y(n321) );
  INVX1 U987 ( .A(n344), .Y(n327) );
  INVX1 U988 ( .A(n348), .Y(n312) );
  INVX1 U989 ( .A(n344), .Y(n328) );
  INVX1 U990 ( .A(n344), .Y(n329) );
  INVX1 U991 ( .A(n343), .Y(n330) );
  INVX1 U992 ( .A(n343), .Y(n331) );
  INVX1 U993 ( .A(n343), .Y(n332) );
  INVX1 U994 ( .A(n342), .Y(n333) );
  INVX1 U995 ( .A(n200), .Y(n212) );
  INVX1 U996 ( .A(n200), .Y(n213) );
  INVX1 U997 ( .A(n263), .Y(n250) );
  INVX1 U998 ( .A(n247), .Y(n251) );
  INVX1 U999 ( .A(n263), .Y(n254) );
  INVX1 U1000 ( .A(n247), .Y(n253) );
  INVX1 U1001 ( .A(n263), .Y(n252) );
  INVX1 U1002 ( .A(n247), .Y(n249) );
  INVX1 U1003 ( .A(n263), .Y(n255) );
  INVX1 U1004 ( .A(n263), .Y(n257) );
  INVX1 U1005 ( .A(n247), .Y(n248) );
  INVX1 U1006 ( .A(n263), .Y(n256) );
  INVX1 U1007 ( .A(n204), .Y(n229) );
  INVX1 U1008 ( .A(n203), .Y(n226) );
  INVX1 U1009 ( .A(n203), .Y(n227) );
  INVX1 U1010 ( .A(n204), .Y(n228) );
  INVX1 U1011 ( .A(n202), .Y(n221) );
  INVX1 U1012 ( .A(n202), .Y(n223) );
  INVX1 U1013 ( .A(n203), .Y(n224) );
  INVX1 U1014 ( .A(n201), .Y(n225) );
  INVX1 U1015 ( .A(n201), .Y(n216) );
  INVX1 U1016 ( .A(n201), .Y(n217) );
  INVX1 U1017 ( .A(n201), .Y(n218) );
  INVX1 U1018 ( .A(n202), .Y(n219) );
  INVX1 U1019 ( .A(n202), .Y(n220) );
  INVX1 U1020 ( .A(n202), .Y(n222) );
  INVX1 U1021 ( .A(n203), .Y(n214) );
  INVX1 U1022 ( .A(n201), .Y(n215) );
  INVX1 U1023 ( .A(n204), .Y(n211) );
  INVX1 U1024 ( .A(n362), .Y(n358) );
  INVX1 U1025 ( .A(n363), .Y(n356) );
  INVX1 U1026 ( .A(n362), .Y(n357) );
  INVX1 U1027 ( .A(n362), .Y(n359) );
  INVX1 U1028 ( .A(n138), .Y(n360) );
  INVX1 U1029 ( .A(n275), .Y(n346) );
  INVX1 U1030 ( .A(n275), .Y(n344) );
  INVX1 U1031 ( .A(n247), .Y(n260) );
  INVX1 U1032 ( .A(n247), .Y(n259) );
  INVX1 U1033 ( .A(n247), .Y(n261) );
  INVX1 U1034 ( .A(n204), .Y(n230) );
  INVX1 U1035 ( .A(n205), .Y(n203) );
  INVX1 U1036 ( .A(n205), .Y(n204) );
  INVX1 U1037 ( .A(n205), .Y(n201) );
  INVX1 U1038 ( .A(n205), .Y(n202) );
  INVX1 U1039 ( .A(n258), .Y(n263) );
  INVX1 U1040 ( .A(n714), .Y(n262) );
  INVX1 U1041 ( .A(n199), .Y(n187) );
  INVX1 U1042 ( .A(n198), .Y(n183) );
  INVX1 U1043 ( .A(n273), .Y(n268) );
  INVX1 U1044 ( .A(n273), .Y(n271) );
  INVX1 U1045 ( .A(n709), .Y(n206) );
  INVX1 U1046 ( .A(n713), .Y(n246) );
  INVX1 U1047 ( .A(n713), .Y(n245) );
  INVX1 U1048 ( .A(n709), .Y(n205) );
  INVX1 U1049 ( .A(n2336), .Y(n745) );
  INVX1 U1050 ( .A(n2402), .Y(n786) );
  INVX1 U1051 ( .A(n2286), .Y(n781) );
  INVX1 U1052 ( .A(n2354), .Y(n764) );
  NOR2X1 U1053 ( .A(n765), .B(n784), .Y(n2267) );
  INVX1 U1054 ( .A(n2326), .Y(n774) );
  NOR2X1 U1055 ( .A(n791), .B(n787), .Y(n2239) );
  INVX1 U1056 ( .A(n2211), .Y(n791) );
  INVX1 U1057 ( .A(n2360), .Y(n751) );
  NAND4X1 U1058 ( .A(n786), .B(n751), .C(n2276), .D(n762), .Y(n2319) );
  NAND2X1 U1059 ( .A(n2343), .B(n139), .Y(n2277) );
  INVX1 U1060 ( .A(n2353), .Y(n770) );
  AOI21X1 U1061 ( .A0(n787), .A1(n754), .B0(n793), .Y(n2439) );
  INVX1 U1062 ( .A(n2473), .Y(n743) );
  INVX1 U1063 ( .A(n2301), .Y(n767) );
  NAND2X1 U1064 ( .A(n760), .B(n752), .Y(n2328) );
  INVX1 U1065 ( .A(n2383), .Y(n748) );
  INVX1 U1066 ( .A(n2252), .Y(n742) );
  NAND2X1 U1067 ( .A(n768), .B(n764), .Y(n2315) );
  NAND2X1 U1068 ( .A(n761), .B(n791), .Y(n2352) );
  NOR2X1 U1069 ( .A(n187), .B(n636), .Y(n637) );
  AOI21XL U1070 ( .A0(next_A[24]), .A1(n341), .B0(n633), .Y(n634) );
  NOR2X1 U1071 ( .A(n187), .B(n632), .Y(n633) );
  INVX1 U1072 ( .A(n138), .Y(n354) );
  NAND2BX1 U1073 ( .AN(n381), .B(n1490), .Y(n1489) );
  INVX1 U1074 ( .A(n274), .Y(n266) );
  INVX1 U1075 ( .A(n184), .Y(n188) );
  INVX1 U1076 ( .A(n184), .Y(n190) );
  INVX1 U1077 ( .A(n184), .Y(n193) );
  INVX1 U1078 ( .A(n184), .Y(n191) );
  INVX1 U1079 ( .A(n184), .Y(n195) );
  INVX1 U1080 ( .A(n184), .Y(n194) );
  INVX1 U1081 ( .A(n184), .Y(n192) );
  INVX1 U1082 ( .A(n140), .Y(n273) );
  INVX1 U1083 ( .A(n184), .Y(n189) );
  INVX1 U1084 ( .A(n2455), .Y(n793) );
  INVX1 U1085 ( .A(n2225), .Y(n788) );
  NAND3X1 U1086 ( .A(n367), .B(n370), .C(n1877), .Y(n1858) );
  AOI31X1 U1087 ( .A0(n2375), .A1(n2376), .A2(n2377), .B0(n264), .Y(N2985) );
  NOR3X1 U1088 ( .A(n2380), .B(n2296), .C(n2370), .Y(n2376) );
  AOI211X1 U1089 ( .A0(n2326), .A1(n1396), .B0(n2378), .C0(n2359), .Y(n2377)
         );
  AOI31X1 U1090 ( .A0(n759), .A1(n783), .A2(n2191), .B0(n264), .Y(N3001) );
  INVX1 U1091 ( .A(n2193), .Y(n783) );
  INVX1 U1092 ( .A(n2194), .Y(n759) );
  AND4X2 U1093 ( .A(n785), .B(n755), .C(n774), .D(n775), .Y(n2191) );
  NOR2X1 U1094 ( .A(n784), .B(n790), .Y(n2286) );
  NOR2X1 U1095 ( .A(n792), .B(n787), .Y(n2402) );
  NOR2X1 U1096 ( .A(n746), .B(n369), .Y(n2336) );
  NOR2X1 U1097 ( .A(n765), .B(n790), .Y(n2354) );
  OAI21XL U1098 ( .A0(n372), .A1(n745), .B0(n2449), .Y(n2463) );
  NAND4X1 U1099 ( .A(n2340), .B(n741), .C(n774), .D(n755), .Y(n2397) );
  INVX1 U1100 ( .A(n2399), .Y(n755) );
  NAND3BX1 U1101 ( .AN(n2251), .B(n745), .C(n741), .Y(n2247) );
  INVX1 U1102 ( .A(n2419), .Y(n746) );
  AOI21X1 U1103 ( .A0(n745), .A1(n2223), .B0(n367), .Y(n2313) );
  INVX1 U1104 ( .A(n2212), .Y(n752) );
  NOR2X1 U1105 ( .A(n779), .B(n752), .Y(n2360) );
  NOR2X1 U1106 ( .A(n782), .B(n765), .Y(n2254) );
  INVX1 U1107 ( .A(n2382), .Y(n784) );
  NOR2X1 U1108 ( .A(n792), .B(n777), .Y(n2251) );
  NOR2X1 U1109 ( .A(n777), .B(n790), .Y(n2326) );
  OAI222XL U1110 ( .A0(n777), .A1(n760), .B0(n792), .B1(n742), .C0(n372), .C1(
        n2242), .Y(n2378) );
  NOR3X1 U1111 ( .A(n367), .B(n787), .C(n789), .Y(n2228) );
  NAND2X1 U1112 ( .A(n2475), .B(n372), .Y(n2243) );
  INVX1 U1113 ( .A(n2297), .Y(n760) );
  NOR2X1 U1114 ( .A(n139), .B(n369), .Y(n2252) );
  NOR2X1 U1115 ( .A(n784), .B(n372), .Y(n2427) );
  NOR2X1 U1116 ( .A(n789), .B(n752), .Y(n2260) );
  OAI22X1 U1117 ( .A0(n372), .A1(n792), .B0(n765), .B1(n789), .Y(n2433) );
  NOR2X1 U1118 ( .A(n761), .B(n790), .Y(n2324) );
  NOR2X1 U1119 ( .A(n2410), .B(n372), .Y(n2301) );
  NOR2X1 U1120 ( .A(n765), .B(n792), .Y(n2296) );
  NOR2X1 U1121 ( .A(n789), .B(n773), .Y(n2343) );
  NAND2X1 U1122 ( .A(n2326), .B(n372), .Y(n2276) );
  INVX1 U1123 ( .A(n2389), .Y(n785) );
  NOR2X1 U1124 ( .A(n773), .B(n790), .Y(n2238) );
  INVX1 U1125 ( .A(n132), .Y(n787) );
  INVX1 U1126 ( .A(n2449), .Y(n778) );
  NOR2X1 U1127 ( .A(n752), .B(n790), .Y(n2383) );
  NOR4BBX1 U1128 ( .AN(n2236), .BN(n2340), .C(n2302), .D(n2360), .Y(n2490) );
  AOI31X1 U1129 ( .A0(n769), .A1(n788), .A2(n2209), .B0(n372), .Y(n2208) );
  INVX1 U1130 ( .A(n2391), .Y(n768) );
  OAI22X1 U1131 ( .A0(n369), .A1(n2226), .B0(n792), .B1(n747), .Y(n2423) );
  INVX1 U1132 ( .A(n1877), .Y(n766) );
  INVX1 U1133 ( .A(n2329), .Y(n754) );
  NOR2X1 U1134 ( .A(n773), .B(n793), .Y(n2353) );
  NAND3X1 U1135 ( .A(n766), .B(n767), .C(n749), .Y(n2437) );
  INVX1 U1136 ( .A(n2325), .Y(n753) );
  NOR2X1 U1137 ( .A(n792), .B(n367), .Y(n2211) );
  AOI21X1 U1138 ( .A0(n2236), .A1(n770), .B0(n372), .Y(n2369) );
  INVX1 U1139 ( .A(n2371), .Y(n762) );
  INVX1 U1140 ( .A(n2335), .Y(n747) );
  NAND2X1 U1141 ( .A(n2272), .B(n2215), .Y(n2287) );
  NAND3X1 U1142 ( .A(n2276), .B(n762), .C(n2340), .Y(n2368) );
  NAND3X1 U1143 ( .A(n2261), .B(n749), .C(n748), .Y(n2453) );
  NAND3X1 U1144 ( .A(n2261), .B(n775), .C(n2209), .Y(n2259) );
  AOI21X1 U1145 ( .A0(n774), .A1(n786), .B0(n372), .Y(n2425) );
  AOI21X1 U1146 ( .A0(n2233), .A1(n786), .B0(n1396), .Y(n2274) );
  NAND2X1 U1147 ( .A(n372), .B(n1877), .Y(n2310) );
  NAND3X1 U1148 ( .A(n767), .B(n775), .C(n2310), .Y(n2307) );
  AOI21X1 U1149 ( .A0(n741), .A1(n766), .B0(n369), .Y(n2373) );
  OAI21XL U1150 ( .A0(n130), .A1(n773), .B0(n753), .Y(n2312) );
  OAI2BB1X1 U1151 ( .A0N(n131), .A1N(n2214), .B0(n2410), .Y(n2457) );
  NAND3X1 U1152 ( .A(n2261), .B(n2236), .C(n2226), .Y(n2284) );
  INVX1 U1153 ( .A(n2266), .Y(n772) );
  NAND2X1 U1154 ( .A(n2419), .B(n2382), .Y(n2237) );
  OAI2BB1X1 U1155 ( .A0N(n367), .A1N(n2343), .B0(n749), .Y(n2398) );
  INVX1 U1156 ( .A(n130), .Y(n761) );
  OAI222XL U1157 ( .A0(n784), .A1(n750), .B0(n752), .B1(n2223), .C0(n788), 
        .C1(n1396), .Y(n2350) );
  INVX1 U1158 ( .A(n2298), .Y(n750) );
  NOR2X1 U1159 ( .A(n369), .B(n793), .Y(n2381) );
  NOR3X1 U1160 ( .A(n777), .B(n793), .C(n367), .Y(n2229) );
  NAND2X1 U1161 ( .A(n2212), .B(n132), .Y(n2258) );
  INVX1 U1162 ( .A(n2300), .Y(n757) );
  NAND2X1 U1163 ( .A(n773), .B(n787), .Y(n2199) );
  INVX1 U1164 ( .A(n2264), .Y(n756) );
  AOI31X1 U1165 ( .A0(n375), .A1(n378), .A2(n376), .B0(n1848), .Y(n714) );
  OAI221XL U1166 ( .A0(n326), .A1(n947), .B0(n1456), .B1(n980), .C0(n1460), 
        .Y(n2528) );
  OAI221XL U1167 ( .A0(n306), .A1(n733), .B0(n222), .B1(n824), .C0(n1756), .Y(
        n2879) );
  AOI21X1 U1168 ( .A0(N880), .A1(n241), .B0(n272), .Y(n1756) );
  OAI221XL U1169 ( .A0(n326), .A1(n732), .B0(n220), .B1(n823), .C0(n1757), .Y(
        n2880) );
  AOI21X1 U1170 ( .A0(N879), .A1(n234), .B0(n272), .Y(n1757) );
  OAI221XL U1171 ( .A0(n334), .A1(n922), .B0(n229), .B1(n947), .C0(n1495), .Y(
        n2560) );
  OAI221XL U1172 ( .A0(n319), .A1(n823), .B0(n224), .B1(n850), .C0(n1725), .Y(
        n2847) );
  AOI21X1 U1173 ( .A0(N911), .A1(n232), .B0(n270), .Y(n1725) );
  OAI221XL U1174 ( .A0(n278), .A1(n851), .B0(n229), .B1(n884), .C0(n1692), .Y(
        n2814) );
  OAI211X1 U1175 ( .A0(n322), .A1(n659), .B0(n658), .C0(n657), .Y(n2957) );
  OAI211X1 U1176 ( .A0(n323), .A1(n656), .B0(n655), .C0(n654), .Y(n2956) );
  INVXL U1177 ( .A(next_A[16]), .Y(n656) );
  INVXL U1178 ( .A(next_A[19]), .Y(n649) );
  OAI211X1 U1179 ( .A0(n324), .A1(n662), .B0(n661), .C0(n660), .Y(n2958) );
  INVXL U1180 ( .A(next_A[14]), .Y(n662) );
  XOR3X2 U1181 ( .A(n176), .B(n165), .C(n157), .Y(f3_A_32[3]) );
  XOR3X2 U1182 ( .A(n177), .B(n166), .C(n158), .Y(f3_A_32[2]) );
  NAND3X1 U1183 ( .A(n630), .B(n629), .C(n628), .Y(n2947) );
  NAND2XL U1184 ( .A(next_E[30]), .B(n342), .Y(n445) );
  NOR2X1 U1185 ( .A(n897), .B(n185), .Y(n470) );
  NOR2X1 U1186 ( .A(n187), .B(n448), .Y(n449) );
  OAI2BB1X1 U1187 ( .A0N(N972), .A1N(n713), .B0(n466), .Y(n2786) );
  OAI2BB1X1 U1188 ( .A0N(N847), .A1N(n713), .B0(n619), .Y(n2944) );
  NOR2X1 U1189 ( .A(n732), .B(n187), .Y(n618) );
  INVXL U1190 ( .A(next_E[19]), .Y(n480) );
  OAI211X1 U1191 ( .A0(n325), .A1(n486), .B0(n485), .C0(n484), .Y(n2794) );
  INVXL U1192 ( .A(next_E[17]), .Y(n486) );
  AOI21XL U1193 ( .A0(next_E[27]), .A1(n283), .B0(n457), .Y(n458) );
  NOR2X1 U1194 ( .A(n187), .B(n456), .Y(n457) );
  OAI2BB1X1 U1195 ( .A0N(N837), .A1N(n713), .B0(n651), .Y(n2954) );
  AOI2BB2X1 U1196 ( .B0(n193), .B1(n163), .A0N(n336), .A1N(n650), .Y(n651) );
  INVXL U1197 ( .A(next_A[18]), .Y(n650) );
  OAI2BB1X1 U1198 ( .A0N(N968), .A1N(n239), .B0(n475), .Y(n2790) );
  AOI2BB2X1 U1199 ( .B0(n189), .B1(n144), .A0N(n334), .A1N(n474), .Y(n475) );
  INVXL U1200 ( .A(next_E[21]), .Y(n474) );
  OAI2BB1X1 U1201 ( .A0N(N840), .A1N(n231), .B0(n644), .Y(n2951) );
  AOI2BB2X1 U1202 ( .B0(n192), .B1(n160), .A0N(n279), .A1N(n643), .Y(n644) );
  INVXL U1203 ( .A(n33), .Y(n643) );
  OAI2BB1X1 U1204 ( .A0N(N841), .A1N(n243), .B0(n642), .Y(n2950) );
  AOI21XL U1205 ( .A0(next_A[22]), .A1(n289), .B0(n641), .Y(n642) );
  NOR2X1 U1206 ( .A(n735), .B(n184), .Y(n610) );
  NOR2X1 U1207 ( .A(n187), .B(n547), .Y(n548) );
  OAI2BB1X1 U1208 ( .A0N(N839), .A1N(n241), .B0(n646), .Y(n2952) );
  AOI2BB2X1 U1209 ( .B0(n191), .B1(n161), .A0N(n300), .A1N(n645), .Y(n646) );
  INVXL U1210 ( .A(next_A[20]), .Y(n645) );
  OAI2BB1X1 U1211 ( .A0N(N967), .A1N(n237), .B0(n477), .Y(n2791) );
  AOI2BB2X1 U1212 ( .B0(n195), .B1(SHA256_result[116]), .A0N(n310), .A1N(n476), 
        .Y(n477) );
  INVXL U1213 ( .A(n32), .Y(n476) );
  OAI2BB1X1 U1214 ( .A0N(N836), .A1N(n235), .B0(n653), .Y(n2955) );
  AOI2BB2X1 U1215 ( .B0(n194), .B1(n164), .A0N(n297), .A1N(n652), .Y(n653) );
  INVXL U1216 ( .A(next_A[17]), .Y(n652) );
  OAI2BB1X1 U1217 ( .A0N(N969), .A1N(n242), .B0(n473), .Y(n2789) );
  AOI21XL U1218 ( .A0(next_E[22]), .A1(n349), .B0(n472), .Y(n473) );
  NOR2X1 U1219 ( .A(n896), .B(n184), .Y(n472) );
  OAI221XL U1220 ( .A0(n333), .A1(n680), .B0(n710), .B1(n679), .C0(n678), .Y(
        n2964) );
  INVX1 U1221 ( .A(next_A[8]), .Y(n680) );
  INVX1 U1222 ( .A(N827), .Y(n679) );
  NAND2X1 U1223 ( .A(n190), .B(n173), .Y(n678) );
  OAI221XL U1224 ( .A0(n335), .A1(n683), .B0(n710), .B1(n682), .C0(n681), .Y(
        n2965) );
  INVX1 U1225 ( .A(next_A[7]), .Y(n683) );
  INVX1 U1226 ( .A(N826), .Y(n682) );
  NAND2X1 U1227 ( .A(n190), .B(n174), .Y(n681) );
  OAI221XL U1228 ( .A0(n295), .A1(n946), .B0(n1456), .B1(n979), .C0(n1461), 
        .Y(n2529) );
  OAI221XL U1229 ( .A0(n322), .A1(n944), .B0(n1456), .B1(n977), .C0(n1463), 
        .Y(n2531) );
  OAI221XL U1230 ( .A0(n1455), .A1(n943), .B0(n1456), .B1(n976), .C0(n1464), 
        .Y(n2532) );
  AOI21X1 U1231 ( .A0(N1067), .A1(n243), .B0(n496), .Y(n1464) );
  OAI221XL U1232 ( .A0(n325), .A1(n942), .B0(n1456), .B1(n975), .C0(n1465), 
        .Y(n2533) );
  OAI221XL U1233 ( .A0(n304), .A1(n941), .B0(n1456), .B1(n974), .C0(n1466), 
        .Y(n2534) );
  OAI221XL U1234 ( .A0(n320), .A1(n940), .B0(n1456), .B1(n973), .C0(n1467), 
        .Y(n2535) );
  OAI221XL U1235 ( .A0(n318), .A1(n934), .B0(n1456), .B1(n967), .C0(n1473), 
        .Y(n2541) );
  OAI221XL U1236 ( .A0(n305), .A1(n933), .B0(n1456), .B1(n966), .C0(n1474), 
        .Y(n2542) );
  OAI221XL U1237 ( .A0(n316), .A1(n930), .B0(n1456), .B1(n963), .C0(n1477), 
        .Y(n2545) );
  OAI221XL U1238 ( .A0(n335), .A1(n929), .B0(n1456), .B1(n962), .C0(n1478), 
        .Y(n2546) );
  OAI221XL U1239 ( .A0(n315), .A1(n927), .B0(n1456), .B1(n960), .C0(n1480), 
        .Y(n2548) );
  OAI221XL U1240 ( .A0(n306), .A1(n730), .B0(n222), .B1(n816), .C0(n1764), .Y(
        n2887) );
  OAI221XL U1241 ( .A0(n336), .A1(n727), .B0(n223), .B1(n813), .C0(n1767), .Y(
        n2890) );
  OAI221XL U1242 ( .A0(n307), .A1(n726), .B0(n221), .B1(n812), .C0(n1768), .Y(
        n2891) );
  OAI221XL U1243 ( .A0(n335), .A1(n731), .B0(n220), .B1(n822), .C0(n1758), .Y(
        n2881) );
  OAI221XL U1244 ( .A0(n313), .A1(n724), .B0(n215), .B1(n810), .C0(n1770), .Y(
        n2893) );
  OAI221XL U1245 ( .A0(n300), .A1(n722), .B0(n214), .B1(n808), .C0(n1772), .Y(
        n2895) );
  OAI221XL U1246 ( .A0(n298), .A1(n718), .B0(n215), .B1(n804), .C0(n1776), .Y(
        n2899) );
  AOI21X1 U1247 ( .A0(N860), .A1(n237), .B0(n270), .Y(n1776) );
  OAI221XL U1248 ( .A0(n324), .A1(n817), .B0(n225), .B1(n844), .C0(n1731), .Y(
        n2853) );
  OAI221XL U1249 ( .A0(n319), .A1(n814), .B0(n216), .B1(n841), .C0(n1734), .Y(
        n2856) );
  OAI221XL U1250 ( .A0(n292), .A1(n813), .B0(n216), .B1(n840), .C0(n1735), .Y(
        n2857) );
  OAI221XL U1251 ( .A0(n279), .A1(n812), .B0(n216), .B1(n839), .C0(n1736), .Y(
        n2858) );
  OAI221XL U1252 ( .A0(n301), .A1(n800), .B0(n219), .B1(n827), .C0(n1748), .Y(
        n2870) );
  OAI221XL U1253 ( .A0(n317), .A1(n799), .B0(n219), .B1(n826), .C0(n1749), .Y(
        n2871) );
  OAI221XL U1254 ( .A0(n300), .A1(n821), .B0(n224), .B1(n848), .C0(n1727), .Y(
        n2849) );
  AOI21X1 U1255 ( .A0(N909), .A1(n11), .B0(n270), .Y(n1727) );
  OAI221XL U1256 ( .A0(n291), .A1(n810), .B0(n217), .B1(n837), .C0(n1738), .Y(
        n2860) );
  OAI221XL U1257 ( .A0(n294), .A1(n809), .B0(n217), .B1(n836), .C0(n1739), .Y(
        n2861) );
  OAI221XL U1258 ( .A0(n338), .A1(n807), .B0(n218), .B1(n834), .C0(n1741), .Y(
        n2863) );
  OAI221XL U1259 ( .A0(n276), .A1(n803), .B0(n218), .B1(n830), .C0(n1745), .Y(
        n2867) );
  OAI221XL U1260 ( .A0(n320), .A1(n917), .B0(n230), .B1(n942), .C0(n1500), .Y(
        n2565) );
  OAI221XL U1261 ( .A0(n276), .A1(n921), .B0(n229), .B1(n946), .C0(n1496), .Y(
        n2561) );
  OAI221XL U1262 ( .A0(n279), .A1(n919), .B0(n230), .B1(n944), .C0(n1498), .Y(
        n2563) );
  OAI221XL U1263 ( .A0(n1455), .A1(n918), .B0(n230), .B1(n943), .C0(n1499), 
        .Y(n2564) );
  OAI221XL U1264 ( .A0(n308), .A1(n909), .B0(n225), .B1(n934), .C0(n1508), .Y(
        n2573) );
  OAI221XL U1265 ( .A0(n317), .A1(n908), .B0(n226), .B1(n933), .C0(n1509), .Y(
        n2574) );
  OAI221XL U1266 ( .A0(n309), .A1(n902), .B0(n227), .B1(n927), .C0(n1515), .Y(
        n2580) );
  OAI221XL U1267 ( .A0(n329), .A1(n898), .B0(n218), .B1(n918), .C0(n1616), .Y(
        n2755) );
  OAI221XL U1268 ( .A0(n297), .A1(n888), .B0(n227), .B1(n908), .C0(n1626), .Y(
        n2765) );
  OAI221XL U1269 ( .A0(n322), .A1(n848), .B0(n228), .B1(n881), .C0(n1695), .Y(
        n2817) );
  OAI221XL U1270 ( .A0(n314), .A1(n725), .B0(n214), .B1(n811), .C0(n1769), .Y(
        n2892) );
  OAI221XL U1271 ( .A0(n302), .A1(n716), .B0(n215), .B1(n802), .C0(n1778), .Y(
        n2901) );
  OAI221XL U1272 ( .A0(n301), .A1(n720), .B0(n214), .B1(n806), .C0(n1774), .Y(
        n2897) );
  OAI221XL U1273 ( .A0(n299), .A1(n719), .B0(n215), .B1(n805), .C0(n1775), .Y(
        n2898) );
  OAI221XL U1274 ( .A0(n96), .A1(n816), .B0(n215), .B1(n843), .C0(n1732), .Y(
        n2854) );
  OAI221XL U1275 ( .A0(n293), .A1(n801), .B0(n219), .B1(n828), .C0(n1747), .Y(
        n2869) );
  OAI221XL U1276 ( .A0(n318), .A1(n822), .B0(n224), .B1(n849), .C0(n1726), .Y(
        n2848) );
  AOI21X1 U1277 ( .A0(N910), .A1(n232), .B0(n270), .Y(n1726) );
  OAI221XL U1278 ( .A0(n277), .A1(n804), .B0(n218), .B1(n831), .C0(n1744), .Y(
        n2866) );
  OAI221XL U1279 ( .A0(n296), .A1(n837), .B0(n221), .B1(n870), .C0(n1706), .Y(
        n2828) );
  AOI21X1 U1280 ( .A0(N930), .A1(n231), .B0(n270), .Y(n1706) );
  OAI221XL U1281 ( .A0(n305), .A1(n911), .B0(n214), .B1(n936), .C0(n1506), .Y(
        n2571) );
  OAI221XL U1282 ( .A0(n1455), .A1(n910), .B0(n225), .B1(n935), .C0(n1507), 
        .Y(n2572) );
  OAI221XL U1283 ( .A0(n339), .A1(n901), .B0(n226), .B1(n926), .C0(n1516), .Y(
        n2581) );
  OAI221XL U1284 ( .A0(n321), .A1(n906), .B0(n226), .B1(n931), .C0(n1511), .Y(
        n2576) );
  OAI221XL U1285 ( .A0(n275), .A1(n892), .B0(n227), .B1(n912), .C0(n1622), .Y(
        n2761) );
  OAI221XL U1286 ( .A0(n316), .A1(n887), .B0(n228), .B1(n907), .C0(n1627), .Y(
        n2766) );
  OAI221XL U1287 ( .A0(n321), .A1(n846), .B0(n228), .B1(n879), .C0(n1697), .Y(
        n2819) );
  OAI221XL U1288 ( .A0(n339), .A1(n844), .B0(n228), .B1(n877), .C0(n1699), .Y(
        n2821) );
  OAI221XL U1289 ( .A0(n275), .A1(n839), .B0(n221), .B1(n872), .C0(n1704), .Y(
        n2826) );
  OAI221XL U1290 ( .A0(n295), .A1(n838), .B0(n221), .B1(n871), .C0(n1705), .Y(
        n2827) );
  OAI221XL U1291 ( .A0(n311), .A1(n827), .B0(n225), .B1(n860), .C0(n1716), .Y(
        n2838) );
  AOI21X1 U1292 ( .A0(N920), .A1(n239), .B0(n270), .Y(n1716) );
  OAI221XL U1293 ( .A0(n332), .A1(n826), .B0(n216), .B1(n859), .C0(n1717), .Y(
        n2839) );
  AOI21X1 U1294 ( .A0(N919), .A1(n240), .B0(n270), .Y(n1717) );
  OAI221XL U1295 ( .A0(n333), .A1(n836), .B0(n222), .B1(n869), .C0(n1707), .Y(
        n2829) );
  AOI21X1 U1296 ( .A0(N929), .A1(n239), .B0(n270), .Y(n1707) );
  OAI221XL U1297 ( .A0(n304), .A1(n834), .B0(n223), .B1(n867), .C0(n1709), .Y(
        n2831) );
  AOI21X1 U1298 ( .A0(N927), .A1(n241), .B0(n270), .Y(n1709) );
  OAI221XL U1299 ( .A0(n331), .A1(n832), .B0(n223), .B1(n865), .C0(n1711), .Y(
        n2833) );
  AOI21X1 U1300 ( .A0(N925), .A1(n242), .B0(n270), .Y(n1711) );
  OAI221XL U1301 ( .A0(n330), .A1(n830), .B0(n223), .B1(n863), .C0(n1713), .Y(
        n2835) );
  AOI21X1 U1302 ( .A0(N923), .A1(n234), .B0(n270), .Y(n1713) );
  OAI221XL U1303 ( .A0(n338), .A1(n841), .B0(n220), .B1(n874), .C0(n1702), .Y(
        n2824) );
  OAI221XL U1304 ( .A0(n277), .A1(n840), .B0(n220), .B1(n873), .C0(n1703), .Y(
        n2825) );
  OAI221XL U1305 ( .A0(n337), .A1(n835), .B0(n222), .B1(n868), .C0(n1708), .Y(
        n2830) );
  AOI21X1 U1306 ( .A0(N928), .A1(n235), .B0(n270), .Y(n1708) );
  NAND3BX1 U1307 ( .AN(n1848), .B(n380), .C(n379), .Y(n381) );
  INVX1 U1308 ( .A(n1858), .Y(n379) );
  OAI211X1 U1309 ( .A0(n278), .A1(n665), .B0(n664), .C0(n663), .Y(n2959) );
  OAI211X1 U1310 ( .A0(n303), .A1(n512), .B0(n511), .C0(n510), .Y(n2802) );
  OAI211X1 U1311 ( .A0(n302), .A1(n517), .B0(n516), .C0(n515), .Y(n2803) );
  NAND2X1 U1312 ( .A(n151), .B(n195), .Y(n516) );
  OAI211X1 U1313 ( .A0(n339), .A1(n525), .B0(n524), .C0(n523), .Y(n2805) );
  OAI211X1 U1314 ( .A0(n303), .A1(n668), .B0(n667), .C0(n666), .Y(n2960) );
  INVX1 U1315 ( .A(next_A[12]), .Y(n668) );
  OAI211X1 U1316 ( .A0(n326), .A1(n677), .B0(n676), .C0(n675), .Y(n2963) );
  INVX1 U1317 ( .A(next_A[9]), .Y(n677) );
  OAI211X1 U1318 ( .A0(n294), .A1(n686), .B0(n685), .C0(n684), .Y(n2966) );
  NAND2X1 U1319 ( .A(N825), .B(n238), .Y(n685) );
  OAI211X1 U1320 ( .A0(n277), .A1(n690), .B0(n689), .C0(n688), .Y(n2967) );
  INVX1 U1321 ( .A(next_A[5]), .Y(n690) );
  OAI211X1 U1322 ( .A0(n313), .A1(n695), .B0(n694), .C0(n693), .Y(n2968) );
  NAND2X1 U1323 ( .A(n177), .B(n197), .Y(n694) );
  OAI211X1 U1324 ( .A0(n301), .A1(n700), .B0(n699), .C0(n698), .Y(n2969) );
  NAND2X1 U1325 ( .A(n178), .B(n192), .Y(n699) );
  NAND2X1 U1326 ( .A(N822), .B(n231), .Y(n698) );
  OAI211X1 U1327 ( .A0(n338), .A1(n704), .B0(n703), .C0(n702), .Y(n2970) );
  INVX1 U1328 ( .A(next_A[2]), .Y(n704) );
  OAI211X1 U1329 ( .A0(n324), .A1(n708), .B0(n707), .C0(n706), .Y(n2971) );
  NAND2BX1 U1330 ( .AN(n575), .B(n574), .Y(n2906) );
  OAI21XL U1331 ( .A0(n797), .A1(n211), .B0(n671), .Y(n575) );
  XOR3X2 U1332 ( .A(n161), .B(n172), .C(n154), .Y(f3_A_32[7]) );
  XOR3X2 U1333 ( .A(n163), .B(n174), .C(n155), .Y(f3_A_32[5]) );
  XOR3X2 U1334 ( .A(n178), .B(n167), .C(n159), .Y(f3_A_32[1]) );
  XOR3X2 U1335 ( .A(n160), .B(n171), .C(n153), .Y(f3_A_32[8]) );
  XOR3X2 U1336 ( .A(n60), .B(n168), .C(n158), .Y(f3_A_32[11]) );
  XOR3X2 U1337 ( .A(n164), .B(n175), .C(n156), .Y(f3_A_32[4]) );
  XOR3X2 U1338 ( .A(n59), .B(n169), .C(n159), .Y(f3_A_32[10]) );
  XOR3X2 U1339 ( .A(n178), .B(n166), .C(n156), .Y(f3_A_32[13]) );
  OAI21XL U1340 ( .A0(n183), .A1(n796), .B0(n1784), .Y(n2907) );
  OAI21XL U1341 ( .A0(n186), .A1(n814), .B0(n1766), .Y(n2889) );
  OAI21XL U1342 ( .A0(n186), .A1(n801), .B0(n1779), .Y(n2902) );
  AOI22X1 U1343 ( .A0(N857), .A1(n232), .B0(n175), .B1(n344), .Y(n1779) );
  OAI21XL U1344 ( .A0(n186), .A1(n800), .B0(n1780), .Y(n2903) );
  OAI21XL U1345 ( .A0(n186), .A1(n799), .B0(n1781), .Y(n2904) );
  OAI21XL U1346 ( .A0(n187), .A1(n821), .B0(n1759), .Y(n2882) );
  AOI22X1 U1347 ( .A0(N877), .A1(n236), .B0(n156), .B1(n348), .Y(n1759) );
  OAI21XL U1348 ( .A0(n186), .A1(n809), .B0(n1771), .Y(n2894) );
  AOI22X1 U1349 ( .A0(N865), .A1(n11), .B0(n167), .B1(n340), .Y(n1771) );
  OAI21XL U1350 ( .A0(n186), .A1(n807), .B0(n1773), .Y(n2896) );
  AOI22X1 U1351 ( .A0(N863), .A1(n239), .B0(n169), .B1(n351), .Y(n1773) );
  OAI21XL U1352 ( .A0(n186), .A1(n803), .B0(n1777), .Y(n2900) );
  AOI22X1 U1353 ( .A0(N859), .A1(n235), .B0(n173), .B1(n351), .Y(n1777) );
  OAI21XL U1354 ( .A0(n183), .A1(n911), .B0(n1623), .Y(n2762) );
  AOI22X1 U1355 ( .A0(N996), .A1(n238), .B0(n146), .B1(n283), .Y(n1623) );
  OAI21XL U1358 ( .A0(n183), .A1(n909), .B0(n1625), .Y(n2764) );
  OAI21XL U1361 ( .A0(n183), .A1(n906), .B0(n1628), .Y(n2767) );
  OAI21XL U1364 ( .A0(n183), .A1(n902), .B0(n1632), .Y(n2771) );
  OAI21XL U1367 ( .A0(n187), .A1(n818), .B0(n1762), .Y(n2885) );
  OAI21XL U1368 ( .A0(n187), .A1(n815), .B0(n1765), .Y(n2888) );
  AOI22X1 U1371 ( .A0(N871), .A1(n233), .B0(n161), .B1(n286), .Y(n1765) );
  OAI21XL U1374 ( .A0(n186), .A1(n798), .B0(n1782), .Y(n2905) );
  OAI21XL U1377 ( .A0(n184), .A1(n915), .B0(n1619), .Y(n2758) );
  AOI22X1 U1382 ( .A0(N1000), .A1(n11), .B0(n144), .B1(n342), .Y(n1619) );
  OAI21XL U1383 ( .A0(n183), .A1(n914), .B0(n1620), .Y(n2759) );
  AOI22X1 U1387 ( .A0(N999), .A1(n243), .B0(SHA256_result[116]), .B1(n343), 
        .Y(n1620) );
  OAI21XL U1391 ( .A0(n183), .A1(n913), .B0(n1621), .Y(n2760) );
  OAI21XL U1396 ( .A0(n185), .A1(n900), .B0(n1634), .Y(n2773) );
  OAI21XL U1399 ( .A0(n183), .A1(n904), .B0(n1630), .Y(n2769) );
  OAI21XL U1400 ( .A0(n183), .A1(n903), .B0(n1631), .Y(n2770) );
  NAND3BX1 U1401 ( .AN(n568), .B(n567), .C(n566), .Y(n2883) );
  OAI21XL U1403 ( .A0(n820), .A1(n212), .B0(n671), .Y(n568) );
  NAND2BX1 U1404 ( .AN(n299), .B(n157), .Y(n567) );
  NAND2X1 U1405 ( .A(N876), .B(n241), .Y(n566) );
  NAND3BX1 U1408 ( .AN(n571), .B(n570), .C(n569), .Y(n2884) );
  OAI21XL U1409 ( .A0(n819), .A1(n211), .B0(n671), .Y(n571) );
  NAND2X1 U1410 ( .A(N875), .B(n234), .Y(n569) );
  NAND2BX1 U1414 ( .AN(n302), .B(n158), .Y(n570) );
  NAND3BX1 U1416 ( .AN(n384), .B(n383), .C(n382), .Y(n2552) );
  NAND2BX1 U1418 ( .AN(n956), .B(n388), .Y(n382) );
  OAI21XL U1420 ( .A0(n315), .A1(n438), .B0(n671), .Y(n384) );
  NAND3BX1 U1421 ( .AN(n387), .B(n386), .C(n385), .Y(n2553) );
  NAND2BX1 U1422 ( .AN(n955), .B(n388), .Y(n385) );
  OAI21XL U1423 ( .A0(n325), .A1(n440), .B0(n671), .Y(n387) );
  NAND3BX1 U1424 ( .AN(n391), .B(n390), .C(n389), .Y(n2556) );
  NAND2BX1 U1425 ( .AN(n952), .B(n388), .Y(n389) );
  OAI21XL U1426 ( .A0(n317), .A1(n87), .B0(n671), .Y(n391) );
  OAI211X1 U1427 ( .A0(n327), .A1(n507), .B0(n506), .C0(n505), .Y(n2801) );
  NAND2X1 U1428 ( .A(n149), .B(n195), .Y(n506) );
  NAND2X1 U1429 ( .A(n498), .B(n497), .Y(n2799) );
  INVX1 U1430 ( .A(n671), .Y(n496) );
  NAND2BX1 U1431 ( .AN(n551), .B(n550), .Y(n2840) );
  OAI21XL U1432 ( .A0(n858), .A1(n211), .B0(n671), .Y(n551) );
  NAND2BX1 U1433 ( .AN(n553), .B(n552), .Y(n2842) );
  OAI21XL U1434 ( .A0(n856), .A1(n230), .B0(n671), .Y(n553) );
  NAND2BX1 U1435 ( .AN(n573), .B(n572), .Y(n2886) );
  OAI21XL U1436 ( .A0(n817), .A1(n211), .B0(n671), .Y(n573) );
  OAI2BB1X1 U1437 ( .A0N(N830), .A1N(n236), .B0(n670), .Y(n2961) );
  AOI2BB2X1 U1438 ( .B0(n188), .B1(n170), .A0N(n309), .A1N(n669), .Y(n670) );
  INVXL U1439 ( .A(next_A[11]), .Y(n669) );
  NAND2X1 U1440 ( .A(n712), .B(n711), .Y(n2972) );
  NAND2X1 U1441 ( .A(n674), .B(n673), .Y(n2962) );
  AOI21X1 U1442 ( .A0(n210), .A1(n171), .B0(n672), .Y(n673) );
  AOI22XL U1443 ( .A0(next_A[10]), .A1(n289), .B0(N829), .B1(n236), .Y(n674)
         );
  INVXL U1444 ( .A(n671), .Y(n672) );
  XOR3X2 U1445 ( .A(n177), .B(n165), .C(n155), .Y(f3_A_32[14]) );
  XOR3X2 U1446 ( .A(n162), .B(n174), .C(n153), .Y(f3_A_32[17]) );
  XOR3X2 U1447 ( .A(n59), .B(n172), .C(n160), .Y(f3_A_32[19]) );
  XOR3X2 U1448 ( .A(n179), .B(n167), .C(n157), .Y(f3_A_32[12]) );
  NOR2X1 U1449 ( .A(round[2]), .B(round[3]), .Y(n2455) );
  AOI31X1 U1450 ( .A0(n2420), .A1(n2421), .A2(n2422), .B0(n264), .Y(N2980) );
  AOI2BB2X1 U1451 ( .B0(n2354), .B1(n369), .A0N(n793), .A1N(n2426), .Y(n2420)
         );
  AOI211X1 U1452 ( .A0(n2286), .A1(n365), .B0(n2423), .C0(n2424), .Y(n2422) );
  AOI31X1 U1453 ( .A0(n2404), .A1(n2405), .A2(n2406), .B0(n264), .Y(N2982) );
  NOR3BX1 U1454 ( .AN(n2410), .B(n2302), .C(n2308), .Y(n2405) );
  AOI211X1 U1455 ( .A0(n2411), .A1(n2389), .B0(n2412), .C0(n2229), .Y(n2404)
         );
  AOI211X1 U1456 ( .A0(n2286), .A1(n373), .B0(n2407), .C0(n2408), .Y(n2406) );
  AOI31X1 U1457 ( .A0(n2347), .A1(n2348), .A2(n2349), .B0(n265), .Y(N2988) );
  AOI211X1 U1458 ( .A0(n2286), .A1(n373), .B0(n2350), .C0(n2235), .Y(n2349) );
  AOI211X1 U1459 ( .A0(n21), .A1(n2352), .B0(n2201), .C0(n2275), .Y(n2348) );
  AOI31X1 U1460 ( .A0(n2464), .A1(n2465), .A2(n2466), .B0(n264), .Y(N2974) );
  AOI221X1 U1461 ( .A0(n2360), .A1(n180), .B0(n2311), .B1(n1396), .C0(n2457), 
        .Y(n2464) );
  NOR4BX1 U1462 ( .AN(n2467), .B(n2239), .C(n2324), .D(n2391), .Y(n2466) );
  AOI31X1 U1463 ( .A0(n2316), .A1(n744), .A2(n2317), .B0(n265), .Y(N2991) );
  AOI222X1 U1464 ( .A0(n2326), .A1(n1396), .B0(n28), .B1(n2328), .C0(n2216), 
        .C1(n2329), .Y(n2316) );
  INVX1 U1465 ( .A(n2322), .Y(n744) );
  AOI211X1 U1466 ( .A0(n2198), .A1(n132), .B0(n2319), .C0(n2320), .Y(n2317) );
  AOI31X1 U1467 ( .A0(n2393), .A1(n2394), .A2(n2395), .B0(n264), .Y(N2983) );
  AOI222X1 U1468 ( .A0(n2402), .A1(n1396), .B0(n2253), .B1(n182), .C0(n2382), 
        .C1(n2403), .Y(n2393) );
  AOI211X1 U1469 ( .A0(n181), .A1(n2396), .B0(n2397), .C0(n2398), .Y(n2395) );
  AOI31X1 U1470 ( .A0(n2482), .A1(n2483), .A2(n2484), .B0(n264), .Y(N2971) );
  NOR3X1 U1471 ( .A(n2213), .B(n2254), .C(n778), .Y(n2483) );
  AOI211X1 U1472 ( .A0(n2298), .A1(n28), .B0(n2485), .C0(n2408), .Y(n2484) );
  AOI31X1 U1473 ( .A0(n2202), .A1(n2203), .A2(n2204), .B0(n265), .Y(N3000) );
  AOI22X1 U1474 ( .A0(n2215), .A1(n2216), .B0(n2217), .B1(n369), .Y(n2202) );
  AOI222X1 U1475 ( .A0(n2211), .A1(n180), .B0(n2212), .B1(n2213), .C0(n2214), 
        .C1(n372), .Y(n2203) );
  AOI211X1 U1476 ( .A0(n2205), .A1(n130), .B0(n2207), .C0(n2208), .Y(n2204) );
  AOI31X1 U1477 ( .A0(n2337), .A1(n2338), .A2(n2339), .B0(n265), .Y(N2989) );
  AOI222X1 U1478 ( .A0(n132), .A1(n2328), .B0(n2344), .B1(n373), .C0(n2345), 
        .C1(n2303), .Y(n2338) );
  NOR4BX1 U1479 ( .AN(n2340), .B(n2251), .C(n2341), .D(n2217), .Y(n2339) );
  OR2X2 U1480 ( .A(n136), .B(n29), .Y(n1974) );
  INVX1 U1482 ( .A(output_enable), .Y(n375) );
  AOI31X1 U1483 ( .A0(n2458), .A1(n2459), .A2(n2460), .B0(n264), .Y(N2975) );
  NOR4BX1 U1484 ( .AN(n774), .B(n2286), .C(n2461), .D(n2254), .Y(n2460) );
  AOI221X1 U1485 ( .A0(n2402), .A1(n373), .B0(n2371), .B1(n372), .C0(n2463), 
        .Y(n2458) );
  AOI31X1 U1486 ( .A0(n2280), .A1(n2281), .A2(n2282), .B0(n265), .Y(N2994) );
  AOI2BB2X1 U1487 ( .B0(n372), .B1(n2286), .A0N(n2287), .A1N(n370), .Y(n2280)
         );
  AOI211X1 U1488 ( .A0(n2283), .A1(n1396), .B0(n2284), .C0(n2285), .Y(n2282)
         );
  AOI31X1 U1489 ( .A0(n2428), .A1(n2429), .A2(n2430), .B0(n264), .Y(N2979) );
  NOR4BX1 U1490 ( .AN(n2243), .B(n2391), .C(n2431), .D(n2432), .Y(n2430) );
  AOI22X1 U1491 ( .A0(n2251), .A1(n182), .B0(n28), .B1(n2433), .Y(n2429) );
  NOR2X1 U1492 ( .A(n2374), .B(n2424), .Y(n2428) );
  AOI31X1 U1493 ( .A0(n2288), .A1(n2289), .A2(n2290), .B0(n265), .Y(N2993) );
  NOR3X1 U1494 ( .A(n2301), .B(n2239), .C(n2302), .Y(n2289) );
  AOI31X1 U1495 ( .A0(n2384), .A1(n2385), .A2(n2386), .B0(n264), .Y(N2984) );
  NOR4BX1 U1496 ( .AN(n2387), .B(n2388), .C(n2389), .D(n2302), .Y(n2386) );
  AOI31X1 U1497 ( .A0(n2365), .A1(n2366), .A2(n2367), .B0(n265), .Y(N2986) );
  NOR4BX1 U1498 ( .AN(n2242), .B(n2368), .C(n2369), .D(n2370), .Y(n2367) );
  AOI211X1 U1499 ( .A0(n2238), .A1(n2215), .B0(n2372), .C0(n2373), .Y(n2366)
         );
  AOI21X1 U1500 ( .A0(n2275), .A1(n365), .B0(n2374), .Y(n2365) );
  AOI31X1 U1501 ( .A0(n2230), .A1(n2231), .A2(n2232), .B0(n265), .Y(N2998) );
  NOR3BX1 U1502 ( .AN(n2237), .B(n2238), .C(n2239), .Y(n2231) );
  NOR3BX1 U1503 ( .AN(n2233), .B(n2234), .C(n2235), .Y(n2232) );
  AOI31X1 U1504 ( .A0(n2487), .A1(n2488), .A2(n2489), .B0(n264), .Y(N2970) );
  AOI222X1 U1505 ( .A0(n28), .A1(n2297), .B0(n2427), .B1(n2216), .C0(n2252), 
        .C1(round[3]), .Y(n2487) );
  AND4X2 U1506 ( .A(n2490), .B(n764), .C(n2242), .D(n2209), .Y(n2489) );
  XOR3X2 U1507 ( .A(n163), .B(n175), .C(n154), .Y(f3_A_32[16]) );
  XOR3X2 U1508 ( .A(n177), .B(n168), .C(n157), .Y(f3_A_32[23]) );
  XOR3X2 U1509 ( .A(n179), .B(n170), .C(n159), .Y(f3_A_32[21]) );
  XOR3X2 U1510 ( .A(n178), .B(n169), .C(n158), .Y(f3_A_32[22]) );
  AOI21X1 U1511 ( .A0(n2451), .A1(n2452), .B0(n264), .Y(N2976) );
  AOI211X1 U1512 ( .A0(n2400), .A1(round[3]), .B0(n2456), .C0(n2457), .Y(n2451) );
  AOI211X1 U1513 ( .A0(n2440), .A1(n372), .B0(n2453), .C0(n2454), .Y(n2452) );
  OAI222XL U1514 ( .A0(n1396), .A1(n776), .B0(n180), .B1(n2226), .C0(n2215), 
        .C1(n787), .Y(n2456) );
  INVX1 U1515 ( .A(n142), .Y(n265) );
  NOR2X1 U1516 ( .A(n2155), .B(n136), .Y(N3189) );
  NOR4X1 U1517 ( .A(n2156), .B(n2157), .C(n2158), .D(n2159), .Y(n2155) );
  NAND4X1 U1518 ( .A(n2186), .B(n2187), .C(n2188), .D(n2189), .Y(n2156) );
  NAND4X1 U1519 ( .A(n2170), .B(n2171), .C(n2172), .D(n2173), .Y(n2158) );
  NOR2X1 U1520 ( .A(n2134), .B(n136), .Y(N3190) );
  NOR4X1 U1521 ( .A(n2135), .B(n2136), .C(n2137), .D(n2138), .Y(n2134) );
  NAND4X1 U1522 ( .A(n2151), .B(n2152), .C(n2153), .D(n2154), .Y(n2135) );
  NAND4X1 U1523 ( .A(n2143), .B(n2144), .C(n2145), .D(n2146), .Y(n2137) );
  NOR2X1 U1524 ( .A(n2113), .B(n136), .Y(N3191) );
  NOR4X1 U1525 ( .A(n2114), .B(n2115), .C(n2116), .D(n2117), .Y(n2113) );
  NAND4X1 U1526 ( .A(n2130), .B(n2131), .C(n2132), .D(n2133), .Y(n2114) );
  NAND4X1 U1527 ( .A(n2122), .B(n2123), .C(n2124), .D(n2125), .Y(n2116) );
  NOR2X1 U1528 ( .A(n2092), .B(n136), .Y(N3192) );
  NOR4X1 U1529 ( .A(n2093), .B(n2094), .C(n2095), .D(n2096), .Y(n2092) );
  NAND4X1 U1530 ( .A(n2109), .B(n2110), .C(n2111), .D(n2112), .Y(n2093) );
  NAND4X1 U1531 ( .A(n2101), .B(n2102), .C(n2103), .D(n2104), .Y(n2095) );
  NOR2X1 U1532 ( .A(n2071), .B(n136), .Y(N3193) );
  NOR4X1 U1533 ( .A(n2072), .B(n2073), .C(n2074), .D(n2075), .Y(n2071) );
  NAND4X1 U1534 ( .A(n2088), .B(n2089), .C(n2090), .D(n2091), .Y(n2072) );
  NAND4X1 U1535 ( .A(n2080), .B(n2081), .C(n2082), .D(n2083), .Y(n2074) );
  NOR2X1 U1536 ( .A(n2050), .B(n136), .Y(N3194) );
  NOR4X1 U1537 ( .A(n2051), .B(n2052), .C(n2053), .D(n2054), .Y(n2050) );
  NAND4X1 U1538 ( .A(n2067), .B(n2068), .C(n2069), .D(n2070), .Y(n2051) );
  NAND4X1 U1539 ( .A(n2059), .B(n2060), .C(n2061), .D(n2062), .Y(n2053) );
  NOR2X1 U1540 ( .A(n2029), .B(n136), .Y(N3195) );
  NOR4X1 U1541 ( .A(n2030), .B(n2031), .C(n2032), .D(n2033), .Y(n2029) );
  NAND4X1 U1542 ( .A(n2046), .B(n2047), .C(n2048), .D(n2049), .Y(n2030) );
  NAND4X1 U1543 ( .A(n2038), .B(n2039), .C(n2040), .D(n2041), .Y(n2032) );
  NOR2X1 U1544 ( .A(n1977), .B(n136), .Y(N3196) );
  NOR4X1 U1545 ( .A(n1978), .B(n1979), .C(n1980), .D(n1981), .Y(n1977) );
  NAND4X1 U1546 ( .A(n2018), .B(n2019), .C(n2020), .D(n2021), .Y(n1978) );
  NAND4X1 U1547 ( .A(n1994), .B(n1995), .C(n1996), .D(n1997), .Y(n1980) );
  OR2X2 U1548 ( .A(N3181), .B(n1974), .Y(N3199) );
  XOR3X2 U1549 ( .A(n176), .B(n167), .C(n156), .Y(f3_A_32[24]) );
  XOR3X2 U1550 ( .A(n164), .B(n173), .C(n154), .Y(f3_A_32[27]) );
  XOR3X2 U1551 ( .A(n166), .B(n175), .C(n155), .Y(f3_A_32[25]) );
  XOR3X2 U1552 ( .A(n163), .B(n172), .C(n153), .Y(f3_A_32[28]) );
  INVX1 U1553 ( .A(n371), .Y(n370) );
  INVX1 U1554 ( .A(n2217), .Y(n749) );
  OAI211X1 U1555 ( .A0(round[2]), .A1(n749), .B0(n2287), .C0(n2310), .Y(n2408)
         );
  NOR2X1 U1556 ( .A(n789), .B(n365), .Y(n2419) );
  INVX1 U1557 ( .A(n2392), .Y(n758) );
  NAND3X1 U1558 ( .A(n745), .B(n2210), .C(n2233), .Y(n2374) );
  NOR2X1 U1559 ( .A(n365), .B(n781), .Y(n2399) );
  XOR3X2 U1560 ( .A(n59), .B(n170), .C(n161), .Y(f3_A_32[30]) );
  OAI2BB1X1 U1561 ( .A0N(n181), .A1N(n2379), .B0(n755), .Y(n2359) );
  INVX1 U1562 ( .A(n2216), .Y(n792) );
  INVX1 U1563 ( .A(n2303), .Y(n790) );
  OAI2BB1X1 U1564 ( .A0N(n372), .A1N(n2381), .B0(n2480), .Y(n2479) );
  AOI31X1 U1565 ( .A0(n772), .A1(n786), .A2(n2351), .B0(n182), .Y(n2481) );
  NOR3X1 U1566 ( .A(n369), .B(n182), .C(n790), .Y(n2391) );
  NOR2X1 U1567 ( .A(n180), .B(n181), .Y(n2382) );
  OAI222XL U1568 ( .A0(n765), .A1(n779), .B0(n2390), .B1(n752), .C0(n21), .C1(
        n746), .Y(n2388) );
  NOR2X1 U1569 ( .A(n2213), .B(n2382), .Y(n2390) );
  OAI222XL U1570 ( .A0(n180), .A1(n751), .B0(n777), .B1(n756), .C0(n372), .C1(
        n2236), .Y(n2234) );
  NOR3X1 U1571 ( .A(n372), .B(round[2]), .C(n787), .Y(n2389) );
  OAI222XL U1572 ( .A0(n182), .A1(n2449), .B0(n761), .B1(n776), .C0(n372), 
        .C1(n768), .Y(n2445) );
  NOR2X1 U1573 ( .A(n2243), .B(round[2]), .Y(n2302) );
  OAI222XL U1574 ( .A0(n139), .A1(n2250), .B0(n2473), .B1(n780), .C0(n2486), 
        .C1(n761), .Y(n2485) );
  INVX1 U1575 ( .A(n2344), .Y(n780) );
  NOR3X1 U1576 ( .A(n2309), .B(n21), .C(n2401), .Y(n2486) );
  NOR2X1 U1577 ( .A(n2252), .B(n2254), .Y(n2321) );
  OAI31X1 U1578 ( .A0(n760), .A1(n181), .A2(round[3]), .B0(n2342), .Y(n2341)
         );
  AOI31X1 U1579 ( .A0(n761), .A1(n792), .A2(n28), .B0(n2343), .Y(n2342) );
  NOR2X1 U1580 ( .A(n777), .B(round[3]), .Y(n2253) );
  NOR3X1 U1581 ( .A(n182), .B(n180), .C(n789), .Y(n2370) );
  NAND2X1 U1582 ( .A(n2475), .B(n182), .Y(n2236) );
  NOR2X1 U1583 ( .A(n752), .B(round[2]), .Y(n2298) );
  NOR2X1 U1584 ( .A(n761), .B(round[2]), .Y(n2297) );
  NOR2X1 U1585 ( .A(n773), .B(round[2]), .Y(n2214) );
  OAI221XL U1586 ( .A0(n773), .A1(n2226), .B0(n761), .B1(n774), .C0(n2409), 
        .Y(n2407) );
  OAI21XL U1587 ( .A0(n2260), .A1(n2268), .B0(n370), .Y(n2409) );
  NOR2X1 U1588 ( .A(n773), .B(round[3]), .Y(n2266) );
  OAI211X1 U1589 ( .A0(n180), .A1(n760), .B0(n742), .C0(n754), .Y(n2278) );
  OAI22X1 U1590 ( .A0(n365), .A1(n785), .B0(n771), .B1(n139), .Y(n2424) );
  NOR3X1 U1591 ( .A(n365), .B(n180), .C(n792), .Y(n2450) );
  AOI221X1 U1592 ( .A0(n743), .A1(n180), .B0(n181), .B1(n372), .C0(n2427), .Y(
        n2426) );
  NAND2X1 U1593 ( .A(n130), .B(n2216), .Y(n2226) );
  INVX1 U1594 ( .A(n21), .Y(n777) );
  NOR2X1 U1595 ( .A(n784), .B(round[3]), .Y(n2475) );
  AOI211X1 U1596 ( .A0(n181), .A1(n2334), .B0(n2254), .C0(n2221), .Y(n2333) );
  OAI21XL U1597 ( .A0(n372), .A1(n790), .B0(n756), .Y(n2334) );
  NOR2X1 U1598 ( .A(n2351), .B(n765), .Y(n2308) );
  AOI31X1 U1599 ( .A0(n770), .A1(n776), .A2(n2250), .B0(n765), .Y(n2249) );
  INVX1 U1600 ( .A(n2213), .Y(n776) );
  NOR2X1 U1601 ( .A(n773), .B(n365), .Y(n2329) );
  NOR2X1 U1602 ( .A(n752), .B(n180), .Y(n2335) );
  OAI211X1 U1603 ( .A0(n180), .A1(round[2]), .B0(n772), .C0(n782), .Y(n2362)
         );
  INVX1 U1604 ( .A(n2205), .Y(n782) );
  NOR2X1 U1605 ( .A(n365), .B(n787), .Y(n2325) );
  NAND2X1 U1606 ( .A(n2325), .B(round[3]), .Y(n2242) );
  OAI211X1 U1607 ( .A0(n765), .A1(n771), .B0(n762), .C0(n2210), .Y(n2207) );
  NOR2X1 U1608 ( .A(n790), .B(n181), .Y(n2272) );
  OAI211X1 U1609 ( .A0(n2418), .A1(n1396), .B0(n2237), .C0(n766), .Y(n2416) );
  AOI21X1 U1610 ( .A0(n21), .A1(n789), .B0(n2344), .Y(n2418) );
  OAI2BB2X1 U1611 ( .B0(n372), .B1(n2351), .A0N(n1396), .A1N(n2221), .Y(n2235)
         );
  NOR2X1 U1612 ( .A(n792), .B(n182), .Y(n2363) );
  NOR2X1 U1613 ( .A(n792), .B(n181), .Y(n2309) );
  OAI21XL U1614 ( .A0(n182), .A1(n793), .B0(n760), .Y(n2403) );
  OAI21XL U1615 ( .A0(n180), .A1(n791), .B0(n2243), .Y(n2193) );
  INVX1 U1616 ( .A(n2400), .Y(n741) );
  NAND2BX1 U1617 ( .AN(n2250), .B(n130), .Y(n2340) );
  NOR3X1 U1618 ( .A(n789), .B(n182), .C(n777), .Y(n2263) );
  INVX1 U1619 ( .A(n2311), .Y(n775) );
  NAND2X1 U1620 ( .A(n2221), .B(n182), .Y(n2410) );
  NAND2X1 U1621 ( .A(n2303), .B(n132), .Y(n2209) );
  NAND2X1 U1622 ( .A(n2198), .B(n21), .Y(n2449) );
  NOR2X1 U1623 ( .A(n785), .B(round[3]), .Y(n2227) );
  NOR2X1 U1624 ( .A(n2236), .B(round[2]), .Y(n2371) );
  AOI21X1 U1625 ( .A0(n2210), .A1(n782), .B0(n1396), .Y(n2438) );
  NAND3BX1 U1626 ( .AN(n2227), .B(n781), .C(n2346), .Y(n2292) );
  NAND3X1 U1627 ( .A(round[3]), .B(n1396), .C(n21), .Y(n2346) );
  CLKINVX3 U1628 ( .A(n373), .Y(n372) );
  NAND3X1 U1629 ( .A(n748), .B(n2277), .C(n2462), .Y(n2461) );
  OAI21XL U1630 ( .A0(n2392), .A1(n2360), .B0(n180), .Y(n2462) );
  INVX1 U1631 ( .A(n2364), .Y(n771) );
  OAI221XL U1632 ( .A0(n372), .A1(n2223), .B0(round[2]), .B1(n753), .C0(n2224), 
        .Y(n2222) );
  OAI21XL U1633 ( .A0(n2225), .A1(n778), .B0(n182), .Y(n2224) );
  OAI21XL U1634 ( .A0(n2195), .A1(n180), .B0(n2196), .Y(n2194) );
  OAI21XL U1635 ( .A0(n137), .A1(n2198), .B0(n2199), .Y(n2196) );
  AOI2BB1X1 U1636 ( .A0N(n2221), .A1N(n2253), .B0(n765), .Y(n2432) );
  AOI21X1 U1637 ( .A0(n2243), .A1(n776), .B0(n182), .Y(n2240) );
  AOI21X1 U1638 ( .A0(n2276), .A1(n782), .B0(n365), .Y(n2412) );
  AOI21X1 U1639 ( .A0(n749), .A1(n747), .B0(round[2]), .Y(n2285) );
  INVX1 U1640 ( .A(n2279), .Y(n769) );
  INVX1 U1641 ( .A(n2283), .Y(n779) );
  NAND3BX1 U1642 ( .AN(n2275), .B(n2276), .C(n2277), .Y(n2273) );
  NAND3X1 U1643 ( .A(n2293), .B(n2294), .C(n2295), .Y(n2291) );
  OAI21XL U1644 ( .A0(n2298), .A1(n137), .B0(n21), .Y(n2293) );
  OAI21XL U1645 ( .A0(n2296), .A1(n2297), .B0(n181), .Y(n2295) );
  OAI21XL U1646 ( .A0(n2205), .A1(n2251), .B0(n2215), .Y(n2294) );
  AOI2BB1X1 U1647 ( .A0N(n2251), .A1N(n2238), .B0(n182), .Y(n2491) );
  AOI2BB1X1 U1648 ( .A0N(n2221), .A1N(n2401), .B0(n372), .Y(n2454) );
  XOR3X2 U1649 ( .A(n60), .B(n169), .C(n160), .Y(f3_A_32[31]) );
  OR2X2 U1650 ( .A(n365), .B(n372), .Y(n139) );
  INVX1 U1651 ( .A(n139), .Y(n2215) );
  INVX1 U1652 ( .A(n28), .Y(n773) );
  NOR3X1 U1653 ( .A(n761), .B(n180), .C(round[3]), .Y(n2431) );
  NAND2X1 U1654 ( .A(n132), .B(n365), .Y(n2300) );
  OAI21XL U1655 ( .A0(n180), .A1(n367), .B0(n2300), .Y(n2441) );
  NOR2X1 U1656 ( .A(n181), .B(n765), .Y(n2474) );
  INVX1 U1657 ( .A(n159), .Y(n636) );
  INVX1 U1658 ( .A(n156), .Y(n624) );
  INVX1 U1659 ( .A(n158), .Y(n632) );
  INVX1 U1660 ( .A(n170), .Y(n720) );
  INVX1 U1661 ( .A(n174), .Y(n716) );
  INVX1 U1662 ( .A(n164), .Y(n726) );
  INVX1 U1663 ( .A(n160), .Y(n730) );
  INVX1 U1664 ( .A(n163), .Y(n727) );
  INVX1 U1665 ( .A(n168), .Y(n722) );
  INVX1 U1666 ( .A(n171), .Y(n719) );
  INVX1 U1667 ( .A(n172), .Y(n718) );
  INVX1 U1668 ( .A(n165), .Y(n725) );
  INVX1 U1669 ( .A(n166), .Y(n724) );
  INVX1 U1670 ( .A(n154), .Y(n733) );
  INVX1 U1671 ( .A(n155), .Y(n731) );
  INVX1 U1672 ( .A(inner_busy), .Y(n374) );
  XOR3X2 U1673 ( .A(SHA256_result[103]), .B(SHA256_result[116]), .C(
        SHA256_result[121]), .Y(f4_E_32[14]) );
  OAI211X1 U1674 ( .A0(n355), .A1(n817), .B0(n52), .C0(n1792), .Y(n2918) );
  NAND2X1 U1675 ( .A(H1[22]), .B(n248), .Y(n1792) );
  OAI211X1 U1676 ( .A0(n355), .A1(n816), .B0(n44), .C0(n1793), .Y(n2919) );
  NAND2X1 U1677 ( .A(H1[21]), .B(n252), .Y(n1793) );
  OAI211X1 U1678 ( .A0(n355), .A1(n813), .B0(n55), .C0(n1794), .Y(n2922) );
  NAND2X1 U1679 ( .A(H1[18]), .B(n249), .Y(n1794) );
  OAI211X1 U1680 ( .A0(n355), .A1(n812), .B0(n50), .C0(n1795), .Y(n2923) );
  NAND2X1 U1681 ( .A(H1[17]), .B(n249), .Y(n1795) );
  OAI211X1 U1682 ( .A0(n359), .A1(n824), .B0(n55), .C0(n1787), .Y(n2911) );
  NAND2X1 U1683 ( .A(H1[29]), .B(n251), .Y(n1787) );
  OAI211X1 U1684 ( .A0(n359), .A1(n823), .B0(n55), .C0(n1788), .Y(n2912) );
  NAND2X1 U1685 ( .A(H1[28]), .B(n255), .Y(n1788) );
  OAI211X1 U1686 ( .A0(n359), .A1(n822), .B0(n44), .C0(n1789), .Y(n2913) );
  NAND2X1 U1687 ( .A(H1[27]), .B(n253), .Y(n1789) );
  OAI211X1 U1688 ( .A0(n355), .A1(n810), .B0(n50), .C0(n1797), .Y(n2925) );
  NAND2X1 U1689 ( .A(H1[15]), .B(n249), .Y(n1797) );
  OAI211X1 U1690 ( .A0(n355), .A1(n808), .B0(n51), .C0(n1798), .Y(n2927) );
  NAND2X1 U1691 ( .A(H1[13]), .B(n249), .Y(n1798) );
  OAI211X1 U1692 ( .A0(n356), .A1(n844), .B0(n54), .C0(n1546), .Y(n2630) );
  NAND2X1 U1693 ( .A(H2[22]), .B(n253), .Y(n1546) );
  OAI211X1 U1694 ( .A0(n356), .A1(n841), .B0(n50), .C0(n1548), .Y(n2633) );
  NAND2X1 U1695 ( .A(H2[19]), .B(n253), .Y(n1548) );
  OAI211X1 U1696 ( .A0(n356), .A1(n840), .B0(n51), .C0(n1549), .Y(n2634) );
  NAND2X1 U1697 ( .A(H2[18]), .B(n253), .Y(n1549) );
  OAI211X1 U1698 ( .A0(n356), .A1(n839), .B0(n52), .C0(n1550), .Y(n2635) );
  NAND2X1 U1699 ( .A(H2[17]), .B(n253), .Y(n1550) );
  NAND2X1 U1700 ( .A(H2[5]), .B(n252), .Y(n1558) );
  NAND2X1 U1701 ( .A(H2[4]), .B(n252), .Y(n1559) );
  OAI211X1 U1702 ( .A0(n356), .A1(n851), .B0(n53), .C0(n1542), .Y(n2623) );
  NAND2X1 U1703 ( .A(H2[29]), .B(n254), .Y(n1542) );
  OAI211X1 U1704 ( .A0(n356), .A1(n848), .B0(n44), .C0(n1545), .Y(n2626) );
  NAND2X1 U1705 ( .A(H2[26]), .B(n253), .Y(n1545) );
  OAI211X1 U1706 ( .A0(n356), .A1(n837), .B0(n54), .C0(n1551), .Y(n2637) );
  NAND2X1 U1707 ( .A(H2[15]), .B(n253), .Y(n1551) );
  OAI211X1 U1708 ( .A0(n356), .A1(n836), .B0(n48), .C0(n1552), .Y(n2638) );
  NAND2X1 U1709 ( .A(H2[14]), .B(n252), .Y(n1552) );
  OAI211X1 U1710 ( .A0(n356), .A1(n835), .B0(n50), .C0(n1553), .Y(n2639) );
  NAND2X1 U1711 ( .A(H2[13]), .B(n252), .Y(n1553) );
  OAI211X1 U1712 ( .A0(n357), .A1(n834), .B0(n44), .C0(n1554), .Y(n2640) );
  NAND2X1 U1713 ( .A(H2[12]), .B(n252), .Y(n1554) );
  NAND2X1 U1714 ( .A(H2[8]), .B(n252), .Y(n1556) );
  OAI211X1 U1715 ( .A0(n355), .A1(n942), .B0(n54), .C0(n1528), .Y(n2596) );
  NAND2X1 U1716 ( .A(H6[23]), .B(n256), .Y(n1528) );
  OAI211X1 U1717 ( .A0(n358), .A1(n947), .B0(n48), .C0(n1523), .Y(n2591) );
  NAND2X1 U1718 ( .A(H6[28]), .B(n257), .Y(n1523) );
  OAI211X1 U1719 ( .A0(n357), .A1(n946), .B0(n48), .C0(n1524), .Y(n2592) );
  NAND2X1 U1720 ( .A(H6[27]), .B(n256), .Y(n1524) );
  OAI211X1 U1721 ( .A0(n355), .A1(n944), .B0(n49), .C0(n1526), .Y(n2594) );
  NAND2X1 U1722 ( .A(H6[25]), .B(n256), .Y(n1526) );
  OAI211X1 U1723 ( .A0(n355), .A1(n943), .B0(n49), .C0(n1527), .Y(n2595) );
  NAND2X1 U1724 ( .A(H6[24]), .B(n253), .Y(n1527) );
  OAI211X1 U1725 ( .A0(n359), .A1(n934), .B0(n50), .C0(n1531), .Y(n2604) );
  NAND2X1 U1726 ( .A(H6[15]), .B(n255), .Y(n1531) );
  OAI211X1 U1727 ( .A0(n354), .A1(n933), .B0(n51), .C0(n1532), .Y(n2605) );
  NAND2X1 U1728 ( .A(H6[14]), .B(n255), .Y(n1532) );
  OAI211X1 U1729 ( .A0(n359), .A1(n910), .B0(n44), .C0(n1602), .Y(n2731) );
  NAND2X1 U1730 ( .A(H5[16]), .B(n250), .Y(n1602) );
  OAI211X1 U1731 ( .A0(n359), .A1(n918), .B0(n44), .C0(n1600), .Y(n2723) );
  NAND2X1 U1732 ( .A(H5[24]), .B(n250), .Y(n1600) );
  OAI211X1 U1733 ( .A0(n359), .A1(n908), .B0(n44), .C0(n1603), .Y(n2733) );
  NAND2X1 U1734 ( .A(H5[14]), .B(n250), .Y(n1603) );
  OAI211X1 U1735 ( .A0(n355), .A1(n795), .B0(n50), .C0(n1804), .Y(n2940) );
  NAND2X1 U1736 ( .A(n90), .B(n249), .Y(n1804) );
  OAI211X1 U1737 ( .A0(n360), .A1(n64), .B0(n56), .C0(n1595), .Y(n2715) );
  NAND2X1 U1738 ( .A(H4[0]), .B(n250), .Y(n1595) );
  OAI211X1 U1739 ( .A0(n358), .A1(n888), .B0(n51), .C0(n1586), .Y(n2701) );
  NAND2X1 U1740 ( .A(H4[14]), .B(n250), .Y(n1586) );
  NAND2X1 U1741 ( .A(H4[5]), .B(n252), .Y(n1590) );
  NAND2X1 U1742 ( .A(H4[4]), .B(n250), .Y(n1591) );
  OAI211X1 U1743 ( .A0(n359), .A1(n820), .B0(n55), .C0(n1790), .Y(n2915) );
  NAND2X1 U1744 ( .A(H1[25]), .B(n250), .Y(n1790) );
  OAI211X1 U1745 ( .A0(n355), .A1(n819), .B0(n44), .C0(n1791), .Y(n2916) );
  NAND2X1 U1746 ( .A(H1[24]), .B(n251), .Y(n1791) );
  OAI211X1 U1747 ( .A0(n360), .A1(n533), .B0(n44), .C0(n1592), .Y(n2712) );
  NAND2X1 U1748 ( .A(H4[3]), .B(n250), .Y(n1592) );
  NAND2X1 U1749 ( .A(H4[1]), .B(n250), .Y(n1594) );
  OAI211X1 U1750 ( .A0(n358), .A1(n892), .B0(n55), .C0(n1584), .Y(n2697) );
  NAND2X1 U1751 ( .A(H4[18]), .B(n253), .Y(n1584) );
  OAI211X1 U1752 ( .A0(n358), .A1(n898), .B0(n50), .C0(n1582), .Y(n2691) );
  NAND2X1 U1753 ( .A(H4[24]), .B(n256), .Y(n1582) );
  NAND2X1 U1754 ( .A(H1[2]), .B(n249), .Y(n1803) );
  OAI211X1 U1755 ( .A0(n361), .A1(n76), .B0(n44), .C0(n1593), .Y(n2713) );
  NAND2X1 U1756 ( .A(H4[2]), .B(n250), .Y(n1593) );
  OAI211X1 U1757 ( .A0(n328), .A1(n451), .B0(n407), .C0(n406), .Y(n2751) );
  AOI21X1 U1758 ( .A0(n210), .A1(SHA256_result[92]), .B0(n266), .Y(n407) );
  NAND2X1 U1759 ( .A(N1007), .B(n231), .Y(n406) );
  NAND2X1 U1760 ( .A(H4[28]), .B(n257), .Y(n1581) );
  NAND2X1 U1761 ( .A(H6[5]), .B(n254), .Y(n1537) );
  OAI211X1 U1762 ( .A0(n357), .A1(n881), .B0(n44), .C0(n1563), .Y(n2657) );
  NAND2X1 U1763 ( .A(H3[26]), .B(n252), .Y(n1563) );
  OAI211X1 U1764 ( .A0(n355), .A1(n811), .B0(n44), .C0(n1796), .Y(n2924) );
  NAND2X1 U1765 ( .A(H1[16]), .B(n249), .Y(n1796) );
  NAND2X1 U1766 ( .A(H1[10]), .B(n249), .Y(n1800) );
  OAI211X1 U1767 ( .A0(n359), .A1(n794), .B0(n56), .C0(n1786), .Y(n2909) );
  NAND2X1 U1768 ( .A(H1[31]), .B(n254), .Y(n1786) );
  OAI211X1 U1769 ( .A0(n356), .A1(n843), .B0(n55), .C0(n1547), .Y(n2631) );
  NAND2X1 U1770 ( .A(H2[21]), .B(n253), .Y(n1547) );
  NAND2X1 U1771 ( .A(H2[6]), .B(n252), .Y(n1557) );
  OAI211X1 U1772 ( .A0(n356), .A1(n850), .B0(n44), .C0(n1543), .Y(n2624) );
  NAND2X1 U1773 ( .A(H2[28]), .B(n254), .Y(n1543) );
  OAI211X1 U1774 ( .A0(n356), .A1(n849), .B0(n56), .C0(n1544), .Y(n2625) );
  NAND2X1 U1775 ( .A(H2[27]), .B(n253), .Y(n1544) );
  NAND2X1 U1776 ( .A(H2[9]), .B(n252), .Y(n1555) );
  OAI211X1 U1777 ( .A0(n357), .A1(n870), .B0(n54), .C0(n1570), .Y(n2668) );
  NAND2X1 U1778 ( .A(H3[15]), .B(n251), .Y(n1570) );
  OAI211X1 U1779 ( .A0(n361), .A1(n936), .B0(n52), .C0(n1529), .Y(n2602) );
  NAND2X1 U1780 ( .A(H6[17]), .B(n256), .Y(n1529) );
  OAI211X1 U1781 ( .A0(n361), .A1(n935), .B0(n45), .C0(n1530), .Y(n2603) );
  NAND2X1 U1782 ( .A(H6[16]), .B(n255), .Y(n1530) );
  OAI211X1 U1783 ( .A0(n354), .A1(n945), .B0(n53), .C0(n1525), .Y(n2593) );
  NAND2X1 U1784 ( .A(H6[26]), .B(n256), .Y(n1525) );
  OAI211X1 U1785 ( .A0(n356), .A1(n931), .B0(n51), .C0(n1533), .Y(n2607) );
  NAND2X1 U1786 ( .A(H6[12]), .B(n254), .Y(n1533) );
  OAI211X1 U1787 ( .A0(n359), .A1(n922), .B0(n48), .C0(n1597), .Y(n2719) );
  NAND2X1 U1788 ( .A(H5[28]), .B(n250), .Y(n1597) );
  OAI211X1 U1789 ( .A0(n359), .A1(n921), .B0(n50), .C0(n1598), .Y(n2720) );
  NAND2X1 U1790 ( .A(H5[27]), .B(n250), .Y(n1598) );
  OAI211X1 U1791 ( .A0(n359), .A1(n919), .B0(n49), .C0(n1599), .Y(n2722) );
  NAND2X1 U1792 ( .A(H5[25]), .B(n250), .Y(n1599) );
  OAI211X1 U1793 ( .A0(n359), .A1(n912), .B0(n53), .C0(n1601), .Y(n2729) );
  NAND2X1 U1794 ( .A(H5[18]), .B(n250), .Y(n1601) );
  OAI211X1 U1795 ( .A0(n359), .A1(n907), .B0(n51), .C0(n1604), .Y(n2734) );
  NAND2X1 U1796 ( .A(H5[13]), .B(n248), .Y(n1604) );
  OAI211X1 U1797 ( .A0(n357), .A1(n879), .B0(n48), .C0(n1564), .Y(n2659) );
  NAND2X1 U1798 ( .A(H3[24]), .B(n252), .Y(n1564) );
  OAI211X1 U1799 ( .A0(n360), .A1(n122), .B0(n53), .C0(n1560), .Y(n2651) );
  OAI211X1 U1800 ( .A0(n357), .A1(n877), .B0(n49), .C0(n1565), .Y(n2661) );
  NAND2X1 U1801 ( .A(H3[22]), .B(n251), .Y(n1565) );
  OAI211X1 U1802 ( .A0(n357), .A1(n872), .B0(n55), .C0(n1568), .Y(n2666) );
  NAND2X1 U1803 ( .A(H3[17]), .B(n251), .Y(n1568) );
  OAI211X1 U1804 ( .A0(n357), .A1(n871), .B0(n48), .C0(n1569), .Y(n2667) );
  NAND2X1 U1805 ( .A(H3[16]), .B(n251), .Y(n1569) );
  NAND2X1 U1806 ( .A(H3[5]), .B(n251), .Y(n1576) );
  NAND2X1 U1807 ( .A(H3[4]), .B(n251), .Y(n1577) );
  OAI211X1 U1808 ( .A0(n358), .A1(n982), .B0(n44), .C0(n1437), .Y(n2494) );
  NAND2X1 U1809 ( .A(H7[30]), .B(n257), .Y(n1437) );
  OAI211X1 U1810 ( .A0(n355), .A1(n980), .B0(n55), .C0(n1438), .Y(n2496) );
  NAND2X1 U1811 ( .A(H7[28]), .B(n255), .Y(n1438) );
  OAI211X1 U1812 ( .A0(n355), .A1(n979), .B0(n56), .C0(n1439), .Y(n2497) );
  NAND2X1 U1813 ( .A(H7[27]), .B(n257), .Y(n1439) );
  OAI211X1 U1814 ( .A0(n355), .A1(n977), .B0(n45), .C0(n1440), .Y(n2499) );
  NAND2X1 U1815 ( .A(H7[25]), .B(n257), .Y(n1440) );
  OAI211X1 U1816 ( .A0(n355), .A1(n967), .B0(n45), .C0(n1445), .Y(n2509) );
  NAND2X1 U1817 ( .A(H7[15]), .B(n257), .Y(n1445) );
  OAI211X1 U1818 ( .A0(n361), .A1(n966), .B0(n50), .C0(n1446), .Y(n2510) );
  NAND2X1 U1819 ( .A(H7[14]), .B(n257), .Y(n1446) );
  OAI211X1 U1820 ( .A0(n357), .A1(n884), .B0(n49), .C0(n1562), .Y(n2654) );
  NAND2X1 U1821 ( .A(H3[29]), .B(n252), .Y(n1562) );
  OAI211X1 U1822 ( .A0(n358), .A1(n869), .B0(n50), .C0(n1571), .Y(n2669) );
  NAND2X1 U1823 ( .A(H3[14]), .B(n251), .Y(n1571) );
  OAI211X1 U1824 ( .A0(n358), .A1(n867), .B0(n52), .C0(n1573), .Y(n2671) );
  NAND2X1 U1825 ( .A(H3[12]), .B(n251), .Y(n1573) );
  NAND2X1 U1826 ( .A(H3[10]), .B(n251), .Y(n1574) );
  NAND2X1 U1827 ( .A(H3[8]), .B(n251), .Y(n1575) );
  OAI211X1 U1828 ( .A0(n357), .A1(n854), .B0(n55), .C0(n1561), .Y(n2652) );
  NAND2X1 U1829 ( .A(H3[31]), .B(n252), .Y(n1561) );
  OAI211X1 U1830 ( .A0(n357), .A1(n874), .B0(n52), .C0(n1566), .Y(n2664) );
  NAND2X1 U1831 ( .A(H3[19]), .B(n251), .Y(n1566) );
  OAI211X1 U1832 ( .A0(n357), .A1(n873), .B0(n44), .C0(n1567), .Y(n2665) );
  NAND2X1 U1833 ( .A(H3[18]), .B(n251), .Y(n1567) );
  OAI211X1 U1834 ( .A0(n358), .A1(n868), .B0(n53), .C0(n1572), .Y(n2670) );
  NAND2X1 U1835 ( .A(H3[13]), .B(n251), .Y(n1572) );
  NAND2X1 U1836 ( .A(H7[3]), .B(n256), .Y(n1451) );
  OAI211X1 U1837 ( .A0(n359), .A1(n899), .B0(n49), .C0(n1596), .Y(n2716) );
  INVX1 U1838 ( .A(SHA256_result[95]), .Y(n899) );
  NAND2X1 U1839 ( .A(H5[31]), .B(n250), .Y(n1596) );
  OAI211X1 U1840 ( .A0(n358), .A1(n893), .B0(n55), .C0(n1583), .Y(n2696) );
  INVX1 U1841 ( .A(n145), .Y(n893) );
  NAND2X1 U1842 ( .A(H4[19]), .B(n252), .Y(n1583) );
  OAI211X1 U1843 ( .A0(n358), .A1(n891), .B0(n56), .C0(n1585), .Y(n2698) );
  INVX1 U1844 ( .A(n146), .Y(n891) );
  NAND2X1 U1845 ( .A(H4[17]), .B(n255), .Y(n1585) );
  OAI211X1 U1846 ( .A0(n358), .A1(n886), .B0(n56), .C0(n1587), .Y(n2703) );
  NAND2X1 U1847 ( .A(H4[12]), .B(n257), .Y(n1587) );
  OAI211X1 U1848 ( .A0(n361), .A1(n734), .B0(n52), .C0(n1860), .Y(n2974) );
  INVX1 U1849 ( .A(n153), .Y(n734) );
  NAND2X1 U1850 ( .A(H0[30]), .B(n249), .Y(n1860) );
  OAI211X1 U1851 ( .A0(n355), .A1(n733), .B0(n44), .C0(n1861), .Y(n2975) );
  NAND2X1 U1852 ( .A(H0[29]), .B(n249), .Y(n1861) );
  OAI211X1 U1853 ( .A0(n360), .A1(n731), .B0(n44), .C0(n1862), .Y(n2977) );
  NAND2X1 U1854 ( .A(H0[27]), .B(n248), .Y(n1862) );
  OAI211X1 U1855 ( .A0(n360), .A1(n627), .B0(n56), .C0(n1863), .Y(n2979) );
  INVX1 U1856 ( .A(n157), .Y(n627) );
  NAND2X1 U1857 ( .A(H0[25]), .B(n248), .Y(n1863) );
  OAI211X1 U1858 ( .A0(n360), .A1(n728), .B0(n44), .C0(n1864), .Y(n2985) );
  INVX1 U1859 ( .A(n162), .Y(n728) );
  NAND2X1 U1860 ( .A(H0[19]), .B(n248), .Y(n1864) );
  OAI211X1 U1861 ( .A0(n360), .A1(n725), .B0(n44), .C0(n1865), .Y(n2988) );
  NAND2X1 U1862 ( .A(H0[16]), .B(n248), .Y(n1865) );
  OAI211X1 U1863 ( .A0(n360), .A1(n724), .B0(n54), .C0(n1866), .Y(n2989) );
  NAND2X1 U1864 ( .A(H0[15]), .B(n248), .Y(n1866) );
  OAI211X1 U1865 ( .A0(n360), .A1(n723), .B0(n55), .C0(n1867), .Y(n2990) );
  INVX1 U1866 ( .A(n167), .Y(n723) );
  NAND2X1 U1867 ( .A(H0[14]), .B(n248), .Y(n1867) );
  OAI211X1 U1868 ( .A0(n360), .A1(n722), .B0(n54), .C0(n1868), .Y(n2991) );
  NAND2X1 U1869 ( .A(H0[13]), .B(n248), .Y(n1868) );
  OAI211X1 U1870 ( .A0(n360), .A1(n719), .B0(n44), .C0(n1869), .Y(n2994) );
  NAND2X1 U1871 ( .A(H0[10]), .B(n248), .Y(n1869) );
  OAI211X1 U1872 ( .A0(n360), .A1(n718), .B0(n56), .C0(n1870), .Y(n2995) );
  NAND2X1 U1873 ( .A(H0[9]), .B(n248), .Y(n1870) );
  OAI211X1 U1874 ( .A0(n360), .A1(n715), .B0(n50), .C0(n1871), .Y(n2998) );
  INVX1 U1875 ( .A(n175), .Y(n715) );
  NAND2X1 U1876 ( .A(H0[6]), .B(n248), .Y(n1871) );
  OAI211X1 U1877 ( .A0(n360), .A1(n701), .B0(n51), .C0(n1873), .Y(n3002) );
  NAND2X1 U1878 ( .A(H0[2]), .B(n248), .Y(n1873) );
  OAI211X1 U1879 ( .A0(n360), .A1(n98), .B0(n49), .C0(n1875), .Y(n3004) );
  NAND2X1 U1880 ( .A(H0[0]), .B(n256), .Y(n1875) );
  XOR3X2 U1881 ( .A(SHA256_result[101]), .B(SHA256_result[114]), .C(
        SHA256_result[119]), .Y(f4_E_32[12]) );
  OAI21XL U1882 ( .A0(n740), .A1(n981), .B0(n1459), .Y(n2527) );
  AOI22X1 U1883 ( .A0(N1072), .A1(n242), .B0(SHA256_result[61]), .B1(n286), 
        .Y(n1459) );
  XOR3X2 U1884 ( .A(n149), .B(n147), .C(n14), .Y(f4_E_32[4]) );
  XOR3X2 U1885 ( .A(SHA256_result[99]), .B(SHA256_result[112]), .C(n144), .Y(
        f4_E_32[10]) );
  XOR3X2 U1886 ( .A(n61), .B(SHA256_result[110]), .C(n145), .Y(f4_E_32[8]) );
  MX2X1 U1887 ( .A(SHA256_result[46]), .B(SHA256_result[78]), .S0(
        SHA256_result[110]), .Y(f1_EFG_32[14]) );
  MX2X1 U1888 ( .A(SHA256_result[43]), .B(SHA256_result[75]), .S0(
        SHA256_result[107]), .Y(f1_EFG_32[11]) );
  XOR3X2 U1889 ( .A(SHA256_result[98]), .B(n147), .C(SHA256_result[116]), .Y(
        f4_E_32[9]) );
  OAI2BB2X1 U1890 ( .B0(n364), .B1(n735), .A0N(H0[31]), .A1N(n258), .Y(n2973)
         );
  OAI2BB2X1 U1891 ( .B0(n364), .B1(n732), .A0N(H0[28]), .A1N(n258), .Y(n2976)
         );
  OAI2BB2X1 U1892 ( .B0(n364), .B1(n796), .A0N(H1[1]), .A1N(n258), .Y(n2939)
         );
  OAI2BB2X1 U1893 ( .B0(n364), .B1(n814), .A0N(H1[19]), .A1N(n253), .Y(n2921)
         );
  OAI2BB2X1 U1894 ( .B0(n364), .B1(n800), .A0N(H1[5]), .A1N(n258), .Y(n2935)
         );
  OAI2BB2X1 U1895 ( .B0(n364), .B1(n821), .A0N(H1[26]), .A1N(n249), .Y(n2914)
         );
  OAI2BB2X1 U1896 ( .B0(n364), .B1(n809), .A0N(H1[14]), .A1N(n258), .Y(n2926)
         );
  OAI2BB2X1 U1897 ( .B0(n364), .B1(n807), .A0N(H1[12]), .A1N(n252), .Y(n2928)
         );
  OAI2BB2X1 U1898 ( .B0(n364), .B1(n838), .A0N(H2[16]), .A1N(n259), .Y(n2636)
         );
  OAI2BB2X1 U1899 ( .B0(n364), .B1(n853), .A0N(H2[31]), .A1N(n261), .Y(n2621)
         );
  OAI2BB2X1 U1900 ( .B0(n364), .B1(n846), .A0N(H2[24]), .A1N(n248), .Y(n2628)
         );
  OAI2BB2X1 U1901 ( .B0(n364), .B1(n941), .A0N(H6[22]), .A1N(n261), .Y(n2597)
         );
  OAI2BB2X1 U1902 ( .B0(n364), .B1(n940), .A0N(H6[21]), .A1N(n261), .Y(n2598)
         );
  OAI2BB2X1 U1903 ( .B0(n364), .B1(n949), .A0N(H6[30]), .A1N(n260), .Y(n2589)
         );
  OAI2BB2X1 U1904 ( .B0(n364), .B1(n917), .A0N(H5[23]), .A1N(n259), .Y(n2724)
         );
  OAI2BB2X1 U1905 ( .B0(n364), .B1(n911), .A0N(H5[17]), .A1N(n259), .Y(n2730)
         );
  OAI2BB2X1 U1906 ( .B0(n364), .B1(n920), .A0N(H5[26]), .A1N(n260), .Y(n2721)
         );
  OAI2BB2X1 U1907 ( .B0(n364), .B1(n909), .A0N(H5[15]), .A1N(n259), .Y(n2732)
         );
  OAI2BB2X1 U1908 ( .B0(n364), .B1(n906), .A0N(H5[12]), .A1N(n259), .Y(n2735)
         );
  OAI2BB2X1 U1909 ( .B0(n364), .B1(n897), .A0N(H4[23]), .A1N(n261), .Y(n2692)
         );
  OAI2BB2X1 U1910 ( .B0(n364), .B1(n896), .A0N(H4[22]), .A1N(n260), .Y(n2693)
         );
  OAI2BB2X1 U1911 ( .B0(n364), .B1(n890), .A0N(H4[16]), .A1N(n260), .Y(n2699)
         );
  OAI2BB2X1 U1912 ( .B0(n364), .B1(n887), .A0N(H4[13]), .A1N(n260), .Y(n2702)
         );
  OAI2BB2X1 U1913 ( .B0(n364), .B1(n818), .A0N(H1[23]), .A1N(n256), .Y(n2917)
         );
  OAI2BB2X1 U1914 ( .B0(n364), .B1(n815), .A0N(H1[20]), .A1N(n257), .Y(n2920)
         );
  OAI2BB2X1 U1915 ( .B0(n364), .B1(n825), .A0N(H1[30]), .A1N(n255), .Y(n2910)
         );
  OAI2BB2X1 U1916 ( .B0(n364), .B1(n798), .A0N(H1[3]), .A1N(n258), .Y(n2937)
         );
  OAI2BB2X1 U1917 ( .B0(n364), .B1(n882), .A0N(H3[27]), .A1N(n250), .Y(n2656)
         );
  OAI2BB2X1 U1918 ( .B0(n364), .B1(n883), .A0N(H3[28]), .A1N(n252), .Y(n2655)
         );
  OAI2BB2X1 U1919 ( .B0(n364), .B1(n845), .A0N(H2[23]), .A1N(n251), .Y(n2629)
         );
  OAI2BB2X1 U1920 ( .B0(n364), .B1(n842), .A0N(H2[20]), .A1N(n258), .Y(n2632)
         );
  OAI2BB2X1 U1921 ( .B0(n364), .B1(n852), .A0N(H2[30]), .A1N(n248), .Y(n2622)
         );
  OAI2BB2X1 U1922 ( .B0(n364), .B1(n847), .A0N(H2[25]), .A1N(n260), .Y(n2627)
         );
  OAI2BB2X1 U1923 ( .B0(n364), .B1(n875), .A0N(H3[20]), .A1N(n261), .Y(n2663)
         );
  OAI2BB2X1 U1924 ( .B0(n364), .B1(n939), .A0N(H6[20]), .A1N(n261), .Y(n2599)
         );
  OAI2BB2X1 U1925 ( .B0(n364), .B1(n938), .A0N(H6[19]), .A1N(n261), .Y(n2600)
         );
  OAI2BB2X1 U1926 ( .B0(n364), .B1(n937), .A0N(H6[18]), .A1N(n261), .Y(n2601)
         );
  OAI2BB2X1 U1927 ( .B0(n364), .B1(n950), .A0N(H6[31]), .A1N(n260), .Y(n2588)
         );
  OAI2BB2X1 U1928 ( .B0(n364), .B1(n948), .A0N(H6[29]), .A1N(n260), .Y(n2590)
         );
  OAI2BB2X1 U1929 ( .B0(n364), .B1(n932), .A0N(H6[13]), .A1N(n261), .Y(n2606)
         );
  OAI2BB2X1 U1930 ( .B0(n364), .B1(n916), .A0N(H5[22]), .A1N(n259), .Y(n2725)
         );
  OAI2BB2X1 U1931 ( .B0(n364), .B1(n915), .A0N(H5[21]), .A1N(n259), .Y(n2726)
         );
  OAI2BB2X1 U1932 ( .B0(n364), .B1(n914), .A0N(H5[20]), .A1N(n259), .Y(n2727)
         );
  OAI2BB2X1 U1933 ( .B0(n364), .B1(n913), .A0N(H5[19]), .A1N(n259), .Y(n2728)
         );
  OAI2BB2X1 U1934 ( .B0(n364), .B1(n924), .A0N(H5[30]), .A1N(n260), .Y(n2717)
         );
  OAI2BB2X1 U1935 ( .B0(n364), .B1(n923), .A0N(H5[29]), .A1N(n260), .Y(n2718)
         );
  OAI2BB2X1 U1936 ( .B0(n364), .B1(n876), .A0N(H3[21]), .A1N(n261), .Y(n2662)
         );
  OAI2BB2X1 U1937 ( .B0(n364), .B1(n972), .A0N(H7[20]), .A1N(n254), .Y(n2504)
         );
  OAI2BB2X1 U1938 ( .B0(n364), .B1(n971), .A0N(H7[19]), .A1N(n259), .Y(n2505)
         );
  OAI2BB2X1 U1939 ( .B0(n364), .B1(n970), .A0N(H7[18]), .A1N(n259), .Y(n2506)
         );
  OAI2BB2X1 U1940 ( .B0(n364), .B1(n969), .A0N(H7[17]), .A1N(n259), .Y(n2507)
         );
  OAI2BB2X1 U1941 ( .B0(n364), .B1(n968), .A0N(H7[16]), .A1N(n259), .Y(n2508)
         );
  OAI2BB2X1 U1942 ( .B0(n364), .B1(n954), .A0N(n91), .A1N(n260), .Y(n2522) );
  OAI2BB2X1 U1943 ( .B0(n364), .B1(n953), .A0N(n92), .A1N(n260), .Y(n2523) );
  OAI2BB2X1 U1944 ( .B0(n364), .B1(n878), .A0N(H3[23]), .A1N(n261), .Y(n2660)
         );
  OAI2BB2X1 U1945 ( .B0(n364), .B1(n857), .A0N(H3[2]), .A1N(n261), .Y(n2681)
         );
  OAI2BB2X1 U1946 ( .B0(n364), .B1(n981), .A0N(H7[29]), .A1N(n256), .Y(n2495)
         );
  OAI2BB2X1 U1947 ( .B0(n364), .B1(n978), .A0N(H7[26]), .A1N(n249), .Y(n2498)
         );
  OAI2BB2X1 U1948 ( .B0(n364), .B1(n965), .A0N(H7[13]), .A1N(n259), .Y(n2511)
         );
  OAI2BB2X1 U1949 ( .B0(n364), .B1(n964), .A0N(H7[12]), .A1N(n259), .Y(n2512)
         );
  OAI2BB2X1 U1950 ( .B0(n364), .B1(n885), .A0N(H3[30]), .A1N(n250), .Y(n2653)
         );
  OAI2BB2X1 U1951 ( .B0(n364), .B1(n951), .A0N(H7[31]), .A1N(n258), .Y(n2493)
         );
  OAI2BB2X1 U1952 ( .B0(n364), .B1(n880), .A0N(H3[25]), .A1N(n261), .Y(n2658)
         );
  OAI21XL U1953 ( .A0(n364), .A1(n640), .B0(n639), .Y(n2982) );
  NAND2X1 U1954 ( .A(H0[22]), .B(n255), .Y(n639) );
  OAI2BB2X1 U1955 ( .B0(n364), .B1(n716), .A0N(H0[7]), .A1N(n258), .Y(n2997)
         );
  OAI2BB2X1 U1956 ( .B0(n364), .B1(n730), .A0N(H0[21]), .A1N(n258), .Y(n2983)
         );
  OAI2BB2X1 U1957 ( .B0(n364), .B1(n727), .A0N(H0[18]), .A1N(n258), .Y(n2986)
         );
  OAI21XL U1958 ( .A0(n364), .A1(n456), .B0(n455), .Y(n2688) );
  NAND2X1 U1959 ( .A(H4[27]), .B(n255), .Y(n455) );
  OAI21XL U1960 ( .A0(n364), .A1(n464), .B0(n463), .Y(n2690) );
  NAND2X1 U1961 ( .A(H4[25]), .B(n255), .Y(n463) );
  OAI2BB2X1 U1962 ( .B0(n364), .B1(n895), .A0N(H4[21]), .A1N(n260), .Y(n2694)
         );
  INVX1 U1963 ( .A(n144), .Y(n895) );
  OAI2BB2X1 U1964 ( .B0(n364), .B1(n894), .A0N(H4[20]), .A1N(n260), .Y(n2695)
         );
  INVX1 U1965 ( .A(SHA256_result[116]), .Y(n894) );
  OAI2BB2X1 U1966 ( .B0(n364), .B1(n889), .A0N(H4[15]), .A1N(n260), .Y(n2700)
         );
  OAI2BB2X1 U1967 ( .B0(n364), .B1(n729), .A0N(H0[20]), .A1N(n258), .Y(n2984)
         );
  INVX1 U1968 ( .A(n161), .Y(n729) );
  OAI21XL U1969 ( .A0(n364), .A1(n547), .B0(n546), .Y(n2684) );
  NAND2X1 U1970 ( .A(H4[31]), .B(n256), .Y(n546) );
  OAI2BB2X1 U1971 ( .B0(n364), .B1(n721), .A0N(H0[12]), .A1N(n258), .Y(n2992)
         );
  INVX1 U1972 ( .A(n169), .Y(n721) );
  INVX1 U1973 ( .A(n173), .Y(n717) );
  OAI21XL U1974 ( .A0(n364), .A1(n438), .B0(n394), .Y(n2615) );
  OAI21XL U1975 ( .A0(n364), .A1(n443), .B0(n429), .Y(n2747) );
  OAI21XL U1976 ( .A0(n364), .A1(n437), .B0(n419), .Y(n2743) );
  OAI21XL U1977 ( .A0(n364), .A1(n67), .B0(n426), .Y(n2746) );
  OAI21XL U1978 ( .A0(n364), .A1(n448), .B0(n447), .Y(n2686) );
  NAND2X1 U1979 ( .A(H4[29]), .B(n254), .Y(n447) );
  OAI21XL U1980 ( .A0(n364), .A1(n460), .B0(n459), .Y(n2689) );
  NAND2X1 U1981 ( .A(H4[26]), .B(n254), .Y(n459) );
  XOR3X2 U1982 ( .A(n43), .B(n146), .C(SHA256_result[118]), .Y(f4_E_32[11]) );
  OAI21XL U1983 ( .A0(n185), .A1(n883), .B0(n1693), .Y(n2815) );
  AOI22X1 U1984 ( .A0(N943), .A1(n713), .B0(SHA256_result[188]), .B1(n280), 
        .Y(n1693) );
  OAI21XL U1985 ( .A0(n364), .A1(n500), .B0(n499), .Y(n2704) );
  NAND2X1 U1986 ( .A(H4[11]), .B(n255), .Y(n499) );
  OAI21XL U1987 ( .A0(n364), .A1(n39), .B0(n518), .Y(n2708) );
  NAND2X1 U1988 ( .A(H4[7]), .B(n255), .Y(n518) );
  OAI21XL U1989 ( .A0(n183), .A1(n948), .B0(n1494), .Y(n2559) );
  AOI22X1 U1990 ( .A0(N1040), .A1(n236), .B0(SHA256_result[93]), .B1(n288), 
        .Y(n1494) );
  OAI21XL U1991 ( .A0(n364), .A1(n442), .B0(n399), .Y(n2617) );
  OAI21XL U1992 ( .A0(n364), .A1(n555), .B0(n554), .Y(n2649) );
  OAI21XL U1993 ( .A0(n364), .A1(n624), .B0(n623), .Y(n2978) );
  NAND2X1 U1994 ( .A(H0[26]), .B(n256), .Y(n623) );
  OAI21XL U1995 ( .A0(n364), .A1(n636), .B0(n635), .Y(n2981) );
  NAND2X1 U1996 ( .A(H0[23]), .B(n257), .Y(n635) );
  OAI21XL U1997 ( .A0(n364), .A1(n632), .B0(n631), .Y(n2980) );
  NAND2X1 U1998 ( .A(H0[24]), .B(n257), .Y(n631) );
  OAI21XL U1999 ( .A0(n364), .A1(n95), .B0(n558), .Y(n2650) );
  OAI21XL U2000 ( .A0(n364), .A1(n70), .B0(n565), .Y(n2876) );
  OAI21XL U2001 ( .A0(n364), .A1(n692), .B0(n691), .Y(n3000) );
  NAND2X1 U2002 ( .A(H0[4]), .B(n257), .Y(n691) );
  OAI21XL U2003 ( .A0(n364), .A1(n697), .B0(n696), .Y(n3001) );
  NAND2X1 U2004 ( .A(H0[3]), .B(n257), .Y(n696) );
  OAI21XL U2005 ( .A0(n364), .A1(n504), .B0(n503), .Y(n2705) );
  NAND2X1 U2006 ( .A(H4[10]), .B(n255), .Y(n503) );
  OAI21XL U2007 ( .A0(n364), .A1(n514), .B0(n513), .Y(n2707) );
  NAND2X1 U2008 ( .A(H4[8]), .B(n254), .Y(n513) );
  NAND2X1 U2009 ( .A(H4[9]), .B(n249), .Y(n1588) );
  NOR2X1 U2010 ( .A(n355), .B(n508), .Y(n509) );
  NAND2X1 U2011 ( .A(H4[6]), .B(n254), .Y(n1589) );
  INVX1 U2012 ( .A(n152), .Y(n522) );
  NAND2X1 U2013 ( .A(H0[5]), .B(n248), .Y(n1872) );
  INVX1 U2014 ( .A(n176), .Y(n687) );
  NAND2X1 U2015 ( .A(H0[1]), .B(n248), .Y(n1874) );
  NOR2X1 U2016 ( .A(n355), .B(n107), .Y(n705) );
  NAND2X1 U2017 ( .A(H4[30]), .B(n253), .Y(n1580) );
  INVX1 U2018 ( .A(n143), .Y(n434) );
  NAND3X1 U2019 ( .A(n469), .B(n468), .C(n467), .Y(n2787) );
  NAND2XL U2020 ( .A(next_E[24]), .B(n287), .Y(n468) );
  OAI211X1 U2021 ( .A0(n296), .A1(n483), .B0(n482), .C0(n481), .Y(n2793) );
  INVXL U2022 ( .A(next_E[18]), .Y(n483) );
  OAI211X1 U2023 ( .A0(n336), .A1(n493), .B0(n492), .C0(n491), .Y(n2797) );
  INVXL U2024 ( .A(next_E[14]), .Y(n493) );
  AOI2BB2X1 U2025 ( .B0(n188), .B1(SHA256_result[112]), .A0N(n275), .A1N(n487), 
        .Y(n488) );
  OAI21XL U2026 ( .A0(n59), .A1(SHA256_result[192]), .B0(n72), .Y(n609) );
  OAI211X1 U2027 ( .A0(n796), .A1(n320), .B0(n562), .C0(n561), .Y(n2874) );
  OAI211X1 U2028 ( .A0(n308), .A1(n456), .B0(n409), .C0(n408), .Y(n2752) );
  NAND2X1 U2029 ( .A(N1006), .B(n232), .Y(n408) );
  OAI211X1 U2030 ( .A0(n319), .A1(n464), .B0(n411), .C0(n410), .Y(n2754) );
  NAND2X1 U2031 ( .A(N1004), .B(n238), .Y(n410) );
  AOI21X1 U2032 ( .A0(n209), .A1(SHA256_result[89]), .B0(n266), .Y(n411) );
  NAND2X1 U2033 ( .A(N1011), .B(n239), .Y(n405) );
  NAND2X1 U2034 ( .A(N1016), .B(n234), .Y(n393) );
  OAI211XL U2035 ( .A0(n276), .A1(n67), .B0(n403), .C0(n402), .Y(n2587) );
  NAND2X1 U2036 ( .A(N1014), .B(n234), .Y(n398) );
  NAND2XL U2037 ( .A(SHA256_result[34]), .B(n193), .Y(n401) );
  NAND2X1 U2038 ( .A(N1013), .B(n243), .Y(n400) );
  OAI211X1 U2039 ( .A0(n306), .A1(n500), .B0(n413), .C0(n412), .Y(n2768) );
  OAI211X1 U2040 ( .A0(n332), .A1(n64), .B0(n431), .C0(n430), .Y(n2779) );
  NAND2X1 U2041 ( .A(N979), .B(n239), .Y(n430) );
  OAI211X1 U2042 ( .A0(n312), .A1(n526), .B0(n418), .C0(n417), .Y(n2774) );
  OAI211X1 U2043 ( .A0(n327), .A1(n80), .B0(n421), .C0(n420), .Y(n2775) );
  OAI211X1 U2044 ( .A0(n323), .A1(n533), .B0(n423), .C0(n422), .Y(n2776) );
  OAI211X1 U2045 ( .A0(n334), .A1(n76), .B0(n425), .C0(n424), .Y(n2777) );
  OAI211X1 U2046 ( .A0(n328), .A1(n521), .B0(n520), .C0(n519), .Y(n2804) );
  NAND2XL U2047 ( .A(SHA256_result[103]), .B(n196), .Y(n520) );
  NAND2X1 U2048 ( .A(N954), .B(n236), .Y(n519) );
  OAI211X1 U2049 ( .A0(n330), .A1(n529), .B0(n528), .C0(n527), .Y(n2806) );
  NAND2X1 U2050 ( .A(N952), .B(n242), .Y(n528) );
  OAI211X1 U2051 ( .A0(n331), .A1(n532), .B0(n531), .C0(n530), .Y(n2807) );
  NAND2X1 U2052 ( .A(N951), .B(n242), .Y(n531) );
  OAI211X1 U2053 ( .A0(n96), .A1(n536), .B0(n535), .C0(n534), .Y(n2808) );
  NAND2X1 U2054 ( .A(N950), .B(n238), .Y(n535) );
  AOI21XL U2055 ( .A0(SHA256_result[99]), .A1(n207), .B0(n267), .Y(n534) );
  OAI211X1 U2056 ( .A0(n329), .A1(n539), .B0(n538), .C0(n537), .Y(n2809) );
  NAND2X1 U2057 ( .A(N949), .B(n233), .Y(n538) );
  AOI21XL U2058 ( .A0(SHA256_result[98]), .A1(n207), .B0(n267), .Y(n537) );
  OAI211X1 U2059 ( .A0(n312), .A1(n542), .B0(n541), .C0(n540), .Y(n2810) );
  NAND2X1 U2060 ( .A(N948), .B(n242), .Y(n541) );
  AOI21XL U2061 ( .A0(n61), .A1(n207), .B0(n267), .Y(n540) );
  OAI211X1 U2062 ( .A0(n298), .A1(n545), .B0(n544), .C0(n543), .Y(n2811) );
  INVX1 U2063 ( .A(next_E[0]), .Y(n545) );
  OAI211X1 U2064 ( .A0(n321), .A1(n798), .B0(n557), .C0(n556), .Y(n2872) );
  OAI211X1 U2065 ( .A0(n333), .A1(n797), .B0(n560), .C0(n559), .Y(n2873) );
  OAI211X1 U2066 ( .A0(n299), .A1(n795), .B0(n564), .C0(n563), .Y(n2875) );
  NAND2X1 U2067 ( .A(N883), .B(n713), .Y(n563) );
  OAI21XL U2068 ( .A0(n740), .A1(n978), .B0(n1462), .Y(n2530) );
  AOI22X1 U2069 ( .A0(N1069), .A1(n241), .B0(SHA256_result[58]), .B1(n282), 
        .Y(n1462) );
  OAI21XL U2070 ( .A0(n740), .A1(n972), .B0(n1468), .Y(n2536) );
  OAI2BB1X1 U2071 ( .A0N(SHA256_result[199]), .A1N(n174), .B0(n602), .Y(
        f2_ABC_32[7]) );
  OAI21XL U2072 ( .A0(SHA256_result[199]), .A1(n174), .B0(SHA256_result[167]), 
        .Y(n602) );
  OAI2BB1X1 U2073 ( .A0N(SHA256_result[198]), .A1N(n175), .B0(n603), .Y(
        f2_ABC_32[6]) );
  OAI21XL U2074 ( .A0(SHA256_result[198]), .A1(n175), .B0(SHA256_result[166]), 
        .Y(n603) );
  OAI2BB1X1 U2075 ( .A0N(SHA256_result[201]), .A1N(n172), .B0(n600), .Y(
        f2_ABC_32[9]) );
  OAI2BB1X1 U2076 ( .A0N(SHA256_result[203]), .A1N(n170), .B0(n598), .Y(
        f2_ABC_32[11]) );
  OAI21XL U2077 ( .A0(SHA256_result[203]), .A1(n170), .B0(SHA256_result[171]), 
        .Y(n598) );
  OAI2BB1X1 U2079 ( .A0N(SHA256_result[197]), .A1N(n176), .B0(n604), .Y(
        f2_ABC_32[5]) );
  OAI21XL U2080 ( .A0(SHA256_result[197]), .A1(n176), .B0(SHA256_result[165]), 
        .Y(n604) );
  OAI2BB1X1 U2081 ( .A0N(SHA256_result[196]), .A1N(n177), .B0(n605), .Y(
        f2_ABC_32[4]) );
  OAI21XL U2082 ( .A0(SHA256_result[196]), .A1(n177), .B0(SHA256_result[164]), 
        .Y(n605) );
  OAI2BB1X1 U2083 ( .A0N(SHA256_result[200]), .A1N(n173), .B0(n601), .Y(
        f2_ABC_32[8]) );
  OAI21XL U2084 ( .A0(SHA256_result[200]), .A1(n173), .B0(SHA256_result[168]), 
        .Y(n601) );
  OAI2BB1X1 U2085 ( .A0N(SHA256_result[202]), .A1N(n171), .B0(n599), .Y(
        f2_ABC_32[10]) );
  OAI21XL U2086 ( .A0(SHA256_result[202]), .A1(n171), .B0(SHA256_result[170]), 
        .Y(n599) );
  XOR3X2 U2087 ( .A(n15), .B(SHA256_result[110]), .C(SHA256_result[123]), .Y(
        f4_E_32[21]) );
  XOR3X2 U2088 ( .A(n150), .B(SHA256_result[118]), .C(SHA256_result[123]), .Y(
        f4_E_32[16]) );
  XOR3X2 U2089 ( .A(n149), .B(SHA256_result[119]), .C(SHA256_result[124]), .Y(
        f4_E_32[17]) );
  XOR3X2 U2090 ( .A(SHA256_result[107]), .B(SHA256_result[120]), .C(n14), .Y(
        f4_E_32[18]) );
  MX2X1 U2091 ( .A(SHA256_result[48]), .B(SHA256_result[80]), .S0(
        SHA256_result[112]), .Y(f1_EFG_32[16]) );
  MX2X1 U2092 ( .A(SHA256_result[50]), .B(SHA256_result[82]), .S0(
        SHA256_result[114]), .Y(f1_EFG_32[18]) );
  XOR3X2 U2093 ( .A(n162), .B(n173), .C(n13), .Y(f3_A_32[6]) );
  XOR3X2 U2094 ( .A(SHA256_result[246]), .B(n170), .C(SHA256_result[255]), .Y(
        f3_A_32[9]) );
  XOR3X2 U2095 ( .A(SHA256_result[121]), .B(n148), .C(n143), .Y(f4_E_32[19])
         );
  XOR3X2 U2096 ( .A(n152), .B(n145), .C(SHA256_result[120]), .Y(f4_E_32[13])
         );
  XOR3X2 U2097 ( .A(n61), .B(n147), .C(SHA256_result[124]), .Y(f4_E_32[22]) );
  XOR3X2 U2098 ( .A(n151), .B(n144), .C(SHA256_result[122]), .Y(f4_E_32[15])
         );
  MX2X1 U2099 ( .A(SHA256_result[49]), .B(SHA256_result[81]), .S0(n146), .Y(
        f1_EFG_32[17]) );
  MX2X1 U2100 ( .A(SHA256_result[47]), .B(SHA256_result[79]), .S0(n147), .Y(
        f1_EFG_32[15]) );
  XOR3X2 U2101 ( .A(n149), .B(SHA256_result[101]), .C(SHA256_result[120]), .Y(
        f4_E_32[31]) );
  OAI21XL U2102 ( .A0(n185), .A1(n838), .B0(n1737), .Y(n2859) );
  OAI21XL U2103 ( .A0(n185), .A1(n846), .B0(n1729), .Y(n2851) );
  AOI22X1 U2104 ( .A0(N907), .A1(n237), .B0(SHA256_result[216]), .B1(n348), 
        .Y(n1729) );
  OAI21XL U2105 ( .A0(n185), .A1(n832), .B0(n1743), .Y(n2865) );
  OAI21XL U2106 ( .A0(n183), .A1(n941), .B0(n1501), .Y(n2566) );
  OAI21XL U2107 ( .A0(n183), .A1(n940), .B0(n1502), .Y(n2567) );
  AOI22X1 U2108 ( .A0(N1032), .A1(n234), .B0(SHA256_result[85]), .B1(n346), 
        .Y(n1502) );
  OAI21XL U2109 ( .A0(n183), .A1(n929), .B0(n1513), .Y(n2578) );
  OAI21XL U2110 ( .A0(n184), .A1(n917), .B0(n1617), .Y(n2756) );
  OAI21XL U2111 ( .A0(n184), .A1(n920), .B0(n1614), .Y(n2753) );
  AOI22X1 U2112 ( .A0(N1005), .A1(n231), .B0(SHA256_result[122]), .B1(n343), 
        .Y(n1614) );
  OAI21XL U2113 ( .A0(n185), .A1(n882), .B0(n1694), .Y(n2816) );
  AOI22X1 U2114 ( .A0(N942), .A1(n232), .B0(SHA256_result[187]), .B1(n283), 
        .Y(n1694) );
  OAI21XL U2115 ( .A0(n185), .A1(n845), .B0(n1730), .Y(n2852) );
  OAI21XL U2116 ( .A0(n185), .A1(n842), .B0(n1733), .Y(n2855) );
  AOI22X1 U2117 ( .A0(N903), .A1(n233), .B0(SHA256_result[212]), .B1(n290), 
        .Y(n1733) );
  OAI21XL U2118 ( .A0(n185), .A1(n829), .B0(n1746), .Y(n2868) );
  OAI21XL U2119 ( .A0(n185), .A1(n847), .B0(n1728), .Y(n2850) );
  AOI22X1 U2120 ( .A0(N908), .A1(n713), .B0(SHA256_result[217]), .B1(n350), 
        .Y(n1728) );
  OAI21XL U2121 ( .A0(n185), .A1(n833), .B0(n1742), .Y(n2864) );
  OAI21XL U2122 ( .A0(n184), .A1(n875), .B0(n1701), .Y(n2823) );
  AOI22X1 U2123 ( .A0(N935), .A1(n240), .B0(SHA256_result[180]), .B1(n282), 
        .Y(n1701) );
  OAI21XL U2124 ( .A0(n183), .A1(n939), .B0(n1503), .Y(n2568) );
  AOI22X1 U2125 ( .A0(N1031), .A1(n239), .B0(SHA256_result[84]), .B1(n340), 
        .Y(n1503) );
  OAI21XL U2126 ( .A0(n186), .A1(n938), .B0(n1504), .Y(n2569) );
  OAI21XL U2127 ( .A0(n183), .A1(n937), .B0(n1505), .Y(n2570) );
  OAI21XL U2128 ( .A0(n186), .A1(n925), .B0(n1517), .Y(n2582) );
  OAI21XL U2129 ( .A0(n186), .A1(n932), .B0(n1510), .Y(n2575) );
  OAI21XL U2130 ( .A0(n183), .A1(n928), .B0(n1514), .Y(n2579) );
  OAI21XL U2131 ( .A0(n184), .A1(n916), .B0(n1618), .Y(n2757) );
  OAI21XL U2132 ( .A0(n184), .A1(n876), .B0(n1700), .Y(n2822) );
  AOI22X1 U2133 ( .A0(N936), .A1(n239), .B0(SHA256_result[181]), .B1(n345), 
        .Y(n1700) );
  OAI21XL U2134 ( .A0(n740), .A1(n971), .B0(n1469), .Y(n2537) );
  OAI21XL U2135 ( .A0(n740), .A1(n970), .B0(n1470), .Y(n2538) );
  OAI21XL U2136 ( .A0(n740), .A1(n969), .B0(n1471), .Y(n2539) );
  OAI21XL U2137 ( .A0(n740), .A1(n968), .B0(n1472), .Y(n2540) );
  OAI21XL U2138 ( .A0(n740), .A1(n959), .B0(n1481), .Y(n2549) );
  OAI21XL U2139 ( .A0(n740), .A1(n958), .B0(n1482), .Y(n2550) );
  OAI21XL U2140 ( .A0(n740), .A1(n957), .B0(n1483), .Y(n2551) );
  OAI21XL U2141 ( .A0(n740), .A1(n954), .B0(n1486), .Y(n2554) );
  OAI21XL U2142 ( .A0(n740), .A1(n953), .B0(n1487), .Y(n2555) );
  OAI21XL U2143 ( .A0(n184), .A1(n878), .B0(n1698), .Y(n2820) );
  AOI22X1 U2144 ( .A0(N938), .A1(n236), .B0(SHA256_result[183]), .B1(n287), 
        .Y(n1698) );
  OAI21XL U2145 ( .A0(n184), .A1(n862), .B0(n1714), .Y(n2836) );
  OAI21XL U2146 ( .A0(n184), .A1(n861), .B0(n1715), .Y(n2837) );
  OAI21XL U2147 ( .A0(n186), .A1(n857), .B0(n1719), .Y(n2841) );
  AOI22XL U2148 ( .A0(N917), .A1(n237), .B0(n94), .B1(n284), .Y(n1719) );
  OAI21XL U2149 ( .A0(n186), .A1(n855), .B0(n1721), .Y(n2843) );
  OAI21XL U2150 ( .A0(n740), .A1(n965), .B0(n1475), .Y(n2543) );
  OAI21XL U2151 ( .A0(n740), .A1(n964), .B0(n1476), .Y(n2544) );
  OAI21XL U2152 ( .A0(n740), .A1(n961), .B0(n1479), .Y(n2547) );
  OAI21XL U2153 ( .A0(n184), .A1(n880), .B0(n1696), .Y(n2818) );
  AOI22X1 U2154 ( .A0(N940), .A1(n231), .B0(SHA256_result[185]), .B1(n341), 
        .Y(n1696) );
  OAI21XL U2155 ( .A0(n184), .A1(n866), .B0(n1710), .Y(n2832) );
  OAI21XL U2156 ( .A0(n184), .A1(n864), .B0(n1712), .Y(n2834) );
  OAI2BB1X1 U2157 ( .A0N(N958), .A1N(n233), .B0(n502), .Y(n2800) );
  AOI2BB2X1 U2158 ( .B0(SHA256_result[107]), .B1(n188), .A0N(n307), .A1N(n501), 
        .Y(n502) );
  INVXL U2159 ( .A(next_E[11]), .Y(n501) );
  OAI2BB1X1 U2160 ( .A0N(N960), .A1N(n239), .B0(n495), .Y(n2798) );
  INVXL U2161 ( .A(next_E[13]), .Y(n494) );
  NAND2BX1 U2162 ( .AN(n577), .B(n576), .Y(n2908) );
  OAI21XL U2163 ( .A0(n795), .A1(n230), .B0(n671), .Y(n577) );
  OAI2BB1X1 U2164 ( .A0N(SHA256_result[209]), .A1N(n164), .B0(n592), .Y(
        f2_ABC_32[17]) );
  OAI21XL U2165 ( .A0(SHA256_result[209]), .A1(n164), .B0(SHA256_result[177]), 
        .Y(n592) );
  OAI2BB1X1 U2166 ( .A0N(SHA256_result[206]), .A1N(n167), .B0(n595), .Y(
        f2_ABC_32[14]) );
  OAI21XL U2167 ( .A0(SHA256_result[206]), .A1(n167), .B0(SHA256_result[174]), 
        .Y(n595) );
  OAI2BB1X1 U2168 ( .A0N(SHA256_result[207]), .A1N(n166), .B0(n594), .Y(
        f2_ABC_32[15]) );
  OAI21XL U2169 ( .A0(SHA256_result[207]), .A1(n166), .B0(SHA256_result[175]), 
        .Y(n594) );
  OAI2BB1X1 U2170 ( .A0N(SHA256_result[204]), .A1N(n169), .B0(n597), .Y(
        f2_ABC_32[12]) );
  OAI21XL U2171 ( .A0(SHA256_result[204]), .A1(n169), .B0(SHA256_result[172]), 
        .Y(n597) );
  OAI2BB1X1 U2172 ( .A0N(SHA256_result[205]), .A1N(n168), .B0(n596), .Y(
        f2_ABC_32[13]) );
  OAI21XL U2173 ( .A0(SHA256_result[205]), .A1(n168), .B0(SHA256_result[173]), 
        .Y(n596) );
  XOR3X2 U2174 ( .A(SHA256_result[98]), .B(SHA256_result[112]), .C(n14), .Y(
        f4_E_32[23]) );
  XOR3X2 U2175 ( .A(SHA256_result[127]), .B(SHA256_result[109]), .C(
        SHA256_result[122]), .Y(f4_E_32[20]) );
  MX2X1 U2176 ( .A(SHA256_result[55]), .B(SHA256_result[87]), .S0(
        SHA256_result[119]), .Y(f1_EFG_32[23]) );
  MX2X1 U2177 ( .A(SHA256_result[54]), .B(SHA256_result[86]), .S0(
        SHA256_result[118]), .Y(f1_EFG_32[22]) );
  MX2X1 U2178 ( .A(SHA256_result[56]), .B(SHA256_result[88]), .S0(
        SHA256_result[120]), .Y(f1_EFG_32[24]) );
  XOR3X2 U2179 ( .A(n176), .B(n164), .C(n13), .Y(f3_A_32[15]) );
  XOR3X2 U2180 ( .A(n161), .B(n173), .C(SHA256_result[255]), .Y(f3_A_32[18])
         );
  XOR3X2 U2181 ( .A(SHA256_result[99]), .B(n146), .C(n143), .Y(f4_E_32[24]) );
  MX2X1 U2182 ( .A(SHA256_result[52]), .B(SHA256_result[84]), .S0(
        SHA256_result[116]), .Y(f1_EFG_32[20]) );
  MX2X1 U2183 ( .A(SHA256_result[53]), .B(SHA256_result[85]), .S0(n144), .Y(
        f1_EFG_32[21]) );
  INVX1 U2184 ( .A(n1488), .Y(n740) );
  OAI21XL U2185 ( .A0(first_block), .A1(n1489), .B0(n1490), .Y(n1488) );
  AOI31X1 U2186 ( .A0(n2476), .A1(n2477), .A2(n2478), .B0(n264), .Y(N2972) );
  AND3X2 U2187 ( .A(n2242), .B(n2210), .C(n781), .Y(n2477) );
  AOI211X1 U2188 ( .A0(n2325), .A1(n1388), .B0(n2479), .C0(n2193), .Y(n2478)
         );
  AOI31X1 U2189 ( .A0(n2442), .A1(n2443), .A2(n2444), .B0(n264), .Y(N2977) );
  NOR3X1 U2190 ( .A(n2301), .B(n2326), .C(n2268), .Y(n2443) );
  AOI211X1 U2191 ( .A0(n2345), .A1(n1388), .B0(n2445), .C0(n2446), .Y(n2444)
         );
  AOI31X1 U2192 ( .A0(n2355), .A1(n2356), .A2(n2357), .B0(n265), .Y(N2987) );
  AOI211X1 U2193 ( .A0(n2297), .A1(n1370), .B0(n2358), .C0(n2359), .Y(n2357)
         );
  AOI31X1 U2194 ( .A0(n2218), .A1(n2219), .A2(n2220), .B0(n265), .Y(N2999) );
  AOI31X1 U2195 ( .A0(n773), .A1(n1383), .A2(n2212), .B0(n2229), .Y(n2218) );
  NOR3BX1 U2196 ( .AN(n2226), .B(n2227), .C(n2228), .Y(n2219) );
  AOI211X1 U2197 ( .A0(n2221), .A1(n130), .B0(n2222), .C0(n763), .Y(n2220) );
  AOI31X1 U2198 ( .A0(n2413), .A1(n2414), .A2(n2415), .B0(n264), .Y(N2981) );
  AOI2BB2X1 U2199 ( .B0(n2214), .B1(n365), .A0N(n2223), .A1N(n765), .Y(n2413)
         );
  AOI22X1 U2200 ( .A0(n2335), .A1(n1383), .B0(n2266), .B1(n372), .Y(n2414) );
  AOI31X1 U2201 ( .A0(n2269), .A1(n2270), .A2(n2271), .B0(n265), .Y(N2995) );
  AOI2BB2X1 U2202 ( .B0(n2253), .B1(n131), .A0N(n2261), .A1N(n370), .Y(n2269)
         );
  AOI22X1 U2203 ( .A0(n2278), .A1(n1383), .B0(n2279), .B1(n2215), .Y(n2270) );
  AOI211X1 U2204 ( .A0(n2272), .A1(n1396), .B0(n2273), .C0(n2274), .Y(n2271)
         );
  AOI31X1 U2205 ( .A0(n2468), .A1(n2469), .A2(n2470), .B0(n264), .Y(N2973) );
  AOI32X1 U2206 ( .A0(n365), .A1(n1388), .A2(n2382), .B0(n130), .B1(n2475), 
        .Y(n2468) );
  AOI211X1 U2207 ( .A0(n2399), .A1(n373), .B0(n2471), .C0(n2463), .Y(n2470) );
  AOI31X1 U2208 ( .A0(n2255), .A1(n2256), .A2(n2257), .B0(n265), .Y(N2996) );
  NOR3BX1 U2209 ( .AN(n2258), .B(n2259), .C(n2260), .Y(n2257) );
  AOI21X1 U2210 ( .A0(n2264), .A1(n180), .B0(n763), .Y(n2255) );
  AOI31X1 U2211 ( .A0(n2434), .A1(n2435), .A2(n2436), .B0(n264), .Y(N2978) );
  AOI222X1 U2212 ( .A0(n2440), .A1(n2360), .B0(n2441), .B1(n1388), .C0(n2363), 
        .C1(n28), .Y(n2435) );
  NOR4BX1 U2213 ( .AN(n768), .B(n2437), .C(n2438), .D(n2439), .Y(n2436) );
  AOI31X1 U2214 ( .A0(n2244), .A1(n2245), .A2(n2246), .B0(n265), .Y(N2997) );
  AOI222X1 U2215 ( .A0(n2252), .A1(n1383), .B0(n2201), .B1(n1370), .C0(n2253), 
        .C1(n373), .Y(n2245) );
  NOR3X1 U2216 ( .A(n2247), .B(n2248), .C(n2249), .Y(n2246) );
  AOI31X1 U2217 ( .A0(n2304), .A1(n2305), .A2(n2306), .B0(n265), .Y(N2992) );
  AOI22X1 U2218 ( .A0(n2315), .A1(n1370), .B0(n2215), .B1(n2213), .Y(n2304) );
  NOR3X1 U2219 ( .A(n2307), .B(n2308), .C(n2248), .Y(n2306) );
  AOI211X1 U2220 ( .A0(n2216), .A1(n2312), .B0(n2313), .C0(n2314), .Y(n2305)
         );
  AOI31X1 U2221 ( .A0(n2330), .A1(n2331), .A2(n2332), .B0(n265), .Y(N2990) );
  AOI222X1 U2222 ( .A0(n2213), .A1(n752), .B0(n2309), .B1(n761), .C0(n2335), 
        .C1(n1383), .Y(n2331) );
  AND4X2 U2223 ( .A(n2333), .B(n785), .C(n2236), .D(n774), .Y(n2332) );
  OAI2BB1X1 U2224 ( .A0N(SHA256_result[214]), .A1N(SHA256_result[246]), .B0(
        n587), .Y(f2_ABC_32[22]) );
  OAI21XL U2225 ( .A0(SHA256_result[214]), .A1(SHA256_result[246]), .B0(
        SHA256_result[182]), .Y(n587) );
  OAI2BB1X1 U2226 ( .A0N(SHA256_result[212]), .A1N(n161), .B0(n589), .Y(
        f2_ABC_32[20]) );
  OAI21XL U2227 ( .A0(SHA256_result[212]), .A1(n161), .B0(SHA256_result[180]), 
        .Y(n589) );
  OAI2BB1X1 U2228 ( .A0N(SHA256_result[213]), .A1N(n160), .B0(n588), .Y(
        f2_ABC_32[21]) );
  OAI21XL U2229 ( .A0(SHA256_result[213]), .A1(n160), .B0(SHA256_result[181]), 
        .Y(n588) );
  OAI2BB1X1 U2230 ( .A0N(SHA256_result[211]), .A1N(n162), .B0(n590), .Y(
        f2_ABC_32[19]) );
  OAI21XL U2231 ( .A0(SHA256_result[211]), .A1(n162), .B0(SHA256_result[179]), 
        .Y(n590) );
  OAI2BB1X1 U2232 ( .A0N(SHA256_result[208]), .A1N(n165), .B0(n593), .Y(
        f2_ABC_32[16]) );
  OAI21XL U2233 ( .A0(SHA256_result[208]), .A1(n165), .B0(SHA256_result[176]), 
        .Y(n593) );
  OAI2BB1X1 U2234 ( .A0N(SHA256_result[210]), .A1N(n163), .B0(n591), .Y(
        f2_ABC_32[18]) );
  OAI21XL U2235 ( .A0(SHA256_result[210]), .A1(n163), .B0(SHA256_result[178]), 
        .Y(n591) );
  XOR3X2 U2236 ( .A(SHA256_result[127]), .B(n43), .C(SHA256_result[114]), .Y(
        f4_E_32[25]) );
  XOR3X2 U2237 ( .A(n15), .B(SHA256_result[101]), .C(n145), .Y(f4_E_32[26]) );
  XOR3X2 U2238 ( .A(n152), .B(n61), .C(SHA256_result[116]), .Y(f4_E_32[27]) );
  XOR3X2 U2239 ( .A(SHA256_result[98]), .B(SHA256_result[103]), .C(n144), .Y(
        f4_E_32[28]) );
  MX2X1 U2240 ( .A(SHA256_result[58]), .B(SHA256_result[90]), .S0(
        SHA256_result[122]), .Y(f1_EFG_32[26]) );
  MX2X1 U2241 ( .A(SHA256_result[60]), .B(SHA256_result[92]), .S0(
        SHA256_result[124]), .Y(f1_EFG_32[28]) );
  XOR3X2 U2242 ( .A(n60), .B(n171), .C(SHA256_result[246]), .Y(f3_A_32[20]) );
  MX2X1 U2243 ( .A(SHA256_result[59]), .B(SHA256_result[91]), .S0(
        SHA256_result[123]), .Y(f1_EFG_32[27]) );
  MX2X1 U2244 ( .A(SHA256_result[57]), .B(SHA256_result[89]), .S0(
        SHA256_result[121]), .Y(f1_EFG_32[25]) );
  OR2X2 U2245 ( .A(N3183), .B(n1974), .Y(N3201) );
  OR2X2 U2246 ( .A(N3182), .B(n1974), .Y(N3200) );
  OR2X2 U2247 ( .A(N3180), .B(n1974), .Y(N3198) );
  OR2X2 U2248 ( .A(n983), .B(n1974), .Y(N3197) );
  OAI2BB1X1 U2249 ( .A0N(SHA256_result[215]), .A1N(n159), .B0(n586), .Y(
        f2_ABC_32[23]) );
  OAI21XL U2250 ( .A0(SHA256_result[215]), .A1(n159), .B0(SHA256_result[183]), 
        .Y(n586) );
  OAI2BB1X1 U2251 ( .A0N(SHA256_result[217]), .A1N(n157), .B0(n584), .Y(
        f2_ABC_32[25]) );
  OAI21XL U2252 ( .A0(SHA256_result[217]), .A1(n157), .B0(SHA256_result[185]), 
        .Y(n584) );
  OAI2BB1X1 U2253 ( .A0N(SHA256_result[216]), .A1N(n158), .B0(n585), .Y(
        f2_ABC_32[24]) );
  OAI21XL U2254 ( .A0(SHA256_result[216]), .A1(n158), .B0(SHA256_result[184]), 
        .Y(n585) );
  OAI2BB1X1 U2255 ( .A0N(SHA256_result[218]), .A1N(n156), .B0(n583), .Y(
        f2_ABC_32[26]) );
  OAI21XL U2256 ( .A0(SHA256_result[218]), .A1(n156), .B0(SHA256_result[186]), 
        .Y(n583) );
  XOR3X2 U2257 ( .A(n150), .B(n43), .C(SHA256_result[119]), .Y(f4_E_32[30]) );
  XOR3X2 U2258 ( .A(n151), .B(SHA256_result[99]), .C(SHA256_result[118]), .Y(
        f4_E_32[29]) );
  MX2X1 U2259 ( .A(SHA256_result[61]), .B(SHA256_result[93]), .S0(n14), .Y(
        f1_EFG_32[29]) );
  XOR3X2 U2260 ( .A(n165), .B(n174), .C(n13), .Y(f3_A_32[26]) );
  MX2X1 U2261 ( .A(SHA256_result[62]), .B(SHA256_result[94]), .S0(n143), .Y(
        f1_EFG_32[30]) );
  NOR2X1 U2262 ( .A(n764), .B(n1370), .Y(n2268) );
  AOI211X1 U2263 ( .A0(n743), .A1(n1383), .B0(n2336), .C0(n2324), .Y(n2472) );
  OAI2BB1X1 U2264 ( .A0N(SHA256_result[220]), .A1N(n13), .B0(n581), .Y(
        f2_ABC_32[28]) );
  OAI21XL U2265 ( .A0(SHA256_result[220]), .A1(n13), .B0(SHA256_result[188]), 
        .Y(n581) );
  OAI2BB1X1 U2266 ( .A0N(SHA256_result[219]), .A1N(n155), .B0(n582), .Y(
        f2_ABC_32[27]) );
  OAI21XL U2267 ( .A0(SHA256_result[219]), .A1(n155), .B0(SHA256_result[187]), 
        .Y(n582) );
  OAI2BB1X1 U2268 ( .A0N(SHA256_result[222]), .A1N(n153), .B0(n579), .Y(
        f2_ABC_32[30]) );
  OAI21XL U2269 ( .A0(SHA256_result[222]), .A1(n153), .B0(SHA256_result[190]), 
        .Y(n579) );
  OAI2BB1X1 U2270 ( .A0N(SHA256_result[221]), .A1N(n154), .B0(n580), .Y(
        f2_ABC_32[29]) );
  OAI21XL U2271 ( .A0(SHA256_result[221]), .A1(n154), .B0(SHA256_result[189]), 
        .Y(n580) );
  INVX1 U2272 ( .A(n2265), .Y(n763) );
  AOI221X1 U2273 ( .A0(n367), .A1(n2266), .B0(n1388), .B1(n2267), .C0(n2268), 
        .Y(n2265) );
  XOR3X2 U2274 ( .A(n162), .B(n171), .C(SHA256_result[255]), .Y(f3_A_32[29])
         );
  MX2X1 U2275 ( .A(SHA256_result[63]), .B(SHA256_result[95]), .S0(
        SHA256_result[127]), .Y(f1_EFG_32[31]) );
  NOR2X1 U2276 ( .A(n777), .B(n1388), .Y(n2213) );
  NOR2X1 U2277 ( .A(n784), .B(n1388), .Y(n2221) );
  OAI222XL U2278 ( .A0(n753), .A1(n1388), .B0(n2323), .B1(n181), .C0(n770), 
        .C1(n373), .Y(n2322) );
  AOI211X1 U2279 ( .A0(n1383), .A1(n2215), .B0(n2296), .C0(n2324), .Y(n2323)
         );
  OAI222XL U2280 ( .A0(n793), .A1(n139), .B0(n373), .B1(n769), .C0(n1388), 
        .C1(n751), .Y(n2358) );
  NOR2X1 U2281 ( .A(read_counter[4]), .B(read_counter[0]), .Y(n2183) );
  NOR2X1 U2282 ( .A(n983), .B(read_counter[4]), .Y(n2182) );
  OAI221XL U2283 ( .A0(n790), .A1(n367), .B0(n1388), .B1(n752), .C0(n2261), 
        .Y(n2396) );
  NOR2X1 U2284 ( .A(n761), .B(n1388), .Y(n2392) );
  NOR3X1 U2285 ( .A(read_counter[2]), .B(read_counter[3]), .C(read_counter[1]), 
        .Y(n2174) );
  NOR2X1 U2286 ( .A(n1383), .B(n372), .Y(n2198) );
  NOR2X1 U2287 ( .A(n773), .B(n1388), .Y(n2279) );
  OAI31X1 U2288 ( .A0(n765), .A1(n787), .A2(n1383), .B0(n2287), .Y(n2361) );
  NOR2X1 U2289 ( .A(n784), .B(n1383), .Y(n2205) );
  NOR2X1 U2290 ( .A(n1383), .B(n369), .Y(n2401) );
  NAND2X1 U2291 ( .A(n778), .B(n1388), .Y(n2210) );
  NAND2X1 U2292 ( .A(n132), .B(n1383), .Y(n2250) );
  NOR2X1 U2293 ( .A(n760), .B(n1383), .Y(n2201) );
  NOR2X1 U2294 ( .A(n2243), .B(n1388), .Y(n2275) );
  NOR2X1 U2295 ( .A(n773), .B(n1383), .Y(n2364) );
  NOR2X1 U2296 ( .A(n139), .B(n1388), .Y(n2262) );
  NAND2X1 U2297 ( .A(n21), .B(n1388), .Y(n2351) );
  NOR2X1 U2298 ( .A(n792), .B(n1370), .Y(n2344) );
  NOR2X1 U2299 ( .A(n761), .B(n1383), .Y(n2379) );
  AOI31X1 U2300 ( .A0(n1388), .A1(n1370), .A2(n2215), .B0(n2308), .Y(n2387) );
  AOI22X1 U2301 ( .A0(n1998), .A1(SHA256_result[132]), .B0(n1999), .B1(
        SHA256_result[140]), .Y(n2083) );
  AOI22X1 U2302 ( .A0(n1998), .A1(SHA256_result[133]), .B0(n1999), .B1(
        SHA256_result[141]), .Y(n2062) );
  AOI22X1 U2303 ( .A0(n1998), .A1(SHA256_result[134]), .B0(n1999), .B1(
        SHA256_result[142]), .Y(n2041) );
  AOI22X1 U2304 ( .A0(n1998), .A1(SHA256_result[135]), .B0(n1999), .B1(
        SHA256_result[143]), .Y(n1997) );
  AOI22X1 U2305 ( .A0(n2000), .A1(SHA256_result[144]), .B0(n2001), .B1(
        SHA256_result[152]), .Y(n2172) );
  AOI22X1 U2306 ( .A0(n2000), .A1(SHA256_result[145]), .B0(n2001), .B1(
        SHA256_result[153]), .Y(n2145) );
  AOI22X1 U2307 ( .A0(n2000), .A1(SHA256_result[146]), .B0(n2001), .B1(
        SHA256_result[154]), .Y(n2124) );
  AOI22X1 U2308 ( .A0(n2000), .A1(SHA256_result[147]), .B0(n2001), .B1(
        SHA256_result[155]), .Y(n2103) );
  AOI22X1 U2309 ( .A0(n2000), .A1(SHA256_result[148]), .B0(n2001), .B1(
        SHA256_result[156]), .Y(n2082) );
  AOI22X1 U2310 ( .A0(n2000), .A1(SHA256_result[149]), .B0(n2001), .B1(
        SHA256_result[157]), .Y(n2061) );
  AOI22X1 U2311 ( .A0(n2000), .A1(SHA256_result[150]), .B0(n2001), .B1(
        SHA256_result[158]), .Y(n2040) );
  AOI22X1 U2312 ( .A0(n2000), .A1(SHA256_result[151]), .B0(n2001), .B1(
        SHA256_result[159]), .Y(n1996) );
  AOI22X1 U2313 ( .A0(n2004), .A1(SHA256_result[180]), .B0(n2005), .B1(
        SHA256_result[188]), .Y(n2080) );
  AOI22X1 U2314 ( .A0(n2004), .A1(SHA256_result[181]), .B0(n2005), .B1(
        SHA256_result[189]), .Y(n2059) );
  AOI22X1 U2315 ( .A0(n2004), .A1(SHA256_result[182]), .B0(n2005), .B1(
        SHA256_result[190]), .Y(n2038) );
  AOI22X1 U2316 ( .A0(n2004), .A1(SHA256_result[183]), .B0(n2005), .B1(
        SHA256_result[191]), .Y(n1994) );
  AOI21X1 U2317 ( .A0(n2242), .A1(n754), .B0(n1388), .Y(n2241) );
  AOI21X1 U2318 ( .A0(n749), .A1(n2258), .B0(n1388), .Y(n2372) );
  NAND4X1 U2319 ( .A(n2160), .B(n2161), .C(n2162), .D(n2163), .Y(n2159) );
  NAND4X1 U2320 ( .A(n2139), .B(n2140), .C(n2141), .D(n2142), .Y(n2138) );
  NAND4X1 U2321 ( .A(n2118), .B(n2119), .C(n2120), .D(n2121), .Y(n2117) );
  NAND4X1 U2322 ( .A(n2097), .B(n2098), .C(n2099), .D(n2100), .Y(n2096) );
  NAND4X1 U2323 ( .A(n2076), .B(n2077), .C(n2078), .D(n2079), .Y(n2075) );
  AOI22X1 U2324 ( .A0(n1988), .A1(SHA256_result[212]), .B0(n1989), .B1(
        SHA256_result[220]), .Y(n2078) );
  NAND4X1 U2325 ( .A(n2055), .B(n2056), .C(n2057), .D(n2058), .Y(n2054) );
  AOI22X1 U2326 ( .A0(n1988), .A1(SHA256_result[213]), .B0(n1989), .B1(
        SHA256_result[221]), .Y(n2057) );
  NAND4X1 U2327 ( .A(n2034), .B(n2035), .C(n2036), .D(n2037), .Y(n2033) );
  AOI22X1 U2328 ( .A0(n1988), .A1(SHA256_result[214]), .B0(n1989), .B1(
        SHA256_result[222]), .Y(n2036) );
  NAND4X1 U2329 ( .A(n1982), .B(n1983), .C(n1984), .D(n1985), .Y(n1981) );
  AOI22X1 U2330 ( .A0(n1988), .A1(SHA256_result[215]), .B0(n1989), .B1(
        SHA256_result[223]), .Y(n1984) );
  NAND4X1 U2331 ( .A(n2178), .B(n2179), .C(n2180), .D(n2181), .Y(n2157) );
  NAND4X1 U2332 ( .A(n2147), .B(n2148), .C(n2149), .D(n2150), .Y(n2136) );
  AOI22XL U2333 ( .A0(n2014), .A1(n61), .B0(n2015), .B1(n150), .Y(n2148) );
  NAND4X1 U2334 ( .A(n2126), .B(n2127), .C(n2128), .D(n2129), .Y(n2115) );
  AOI22XL U2335 ( .A0(n2014), .A1(SHA256_result[98]), .B0(n2015), .B1(n149), 
        .Y(n2127) );
  NAND4X1 U2336 ( .A(n2105), .B(n2106), .C(n2107), .D(n2108), .Y(n2094) );
  AOI22XL U2337 ( .A0(n2014), .A1(SHA256_result[99]), .B0(n2015), .B1(
        SHA256_result[107]), .Y(n2106) );
  NAND4X1 U2338 ( .A(n2084), .B(n2085), .C(n2086), .D(n2087), .Y(n2073) );
  NAND4X1 U2339 ( .A(n2063), .B(n2064), .C(n2065), .D(n2066), .Y(n2052) );
  NAND4X1 U2340 ( .A(n2042), .B(n2043), .C(n2044), .D(n2045), .Y(n2031) );
  NAND4X1 U2341 ( .A(n2006), .B(n2007), .C(n2008), .D(n2009), .Y(n1979) );
  AOI22XL U2342 ( .A0(n2014), .A1(SHA256_result[103]), .B0(n2015), .B1(n147), 
        .Y(n2007) );
  NOR2BX1 U2343 ( .AN(n2185), .B(read_counter[3]), .Y(n2175) );
  OAI21XL U2344 ( .A0(round[3]), .A1(n2447), .B0(n2448), .Y(n2446) );
  AOI22X1 U2345 ( .A0(n761), .A1(n1370), .B0(n2212), .B1(n180), .Y(n2447) );
  OAI21XL U2346 ( .A0(n2260), .A1(n2403), .B0(n369), .Y(n2448) );
  INVX1 U2347 ( .A(read_counter[1]), .Y(n984) );
  BUFX3 U2348 ( .A(n371), .Y(n180) );
  NOR2X1 U2349 ( .A(n984), .B(read_counter[2]), .Y(n2185) );
  OAI2BB1X1 U2350 ( .A0N(SHA256_result[223]), .A1N(SHA256_result[255]), .B0(
        n578), .Y(f2_ABC_32[31]) );
  OAI21XL U2351 ( .A0(SHA256_result[223]), .A1(SHA256_result[255]), .B0(
        SHA256_result[191]), .Y(n578) );
  AND3X2 U2352 ( .A(read_counter[2]), .B(read_counter[1]), .C(read_counter[3]), 
        .Y(n2169) );
  NOR2X1 U2353 ( .A(n985), .B(read_counter[3]), .Y(n2190) );
  INVX1 U2354 ( .A(read_counter[2]), .Y(n985) );
  INVX1 U2355 ( .A(read_counter[0]), .Y(n983) );
  NOR2X1 U2356 ( .A(n1388), .B(n369), .Y(n2440) );
  NOR3X1 U2357 ( .A(n752), .B(n1383), .C(n1370), .Y(n2314) );
  INVX1 U2358 ( .A(SHA256_result[218]), .Y(n821) );
  INVX1 U2359 ( .A(SHA256_result[191]), .Y(n853) );
  INVX1 U2360 ( .A(SHA256_result[184]), .Y(n846) );
  INVX1 U2361 ( .A(SHA256_result[62]), .Y(n949) );
  INVX1 U2362 ( .A(SHA256_result[90]), .Y(n920) );
  INVX1 U2363 ( .A(SHA256_result[214]), .Y(n817) );
  INVX1 U2364 ( .A(SHA256_result[215]), .Y(n818) );
  INVX1 U2365 ( .A(SHA256_result[212]), .Y(n815) );
  INVX1 U2366 ( .A(SHA256_result[213]), .Y(n816) );
  INVX1 U2367 ( .A(SHA256_result[222]), .Y(n825) );
  INVX1 U2368 ( .A(SHA256_result[221]), .Y(n824) );
  INVX1 U2369 ( .A(SHA256_result[220]), .Y(n823) );
  INVX1 U2370 ( .A(SHA256_result[219]), .Y(n822) );
  INVX1 U2371 ( .A(SHA256_result[155]), .Y(n882) );
  INVX1 U2372 ( .A(SHA256_result[156]), .Y(n883) );
  INVX1 U2373 ( .A(SHA256_result[183]), .Y(n845) );
  INVX1 U2374 ( .A(SHA256_result[180]), .Y(n842) );
  INVX1 U2375 ( .A(SHA256_result[182]), .Y(n844) );
  INVX1 U2376 ( .A(SHA256_result[190]), .Y(n852) );
  INVX1 U2377 ( .A(SHA256_result[185]), .Y(n847) );
  INVX1 U2378 ( .A(SHA256_result[189]), .Y(n851) );
  INVX1 U2379 ( .A(SHA256_result[186]), .Y(n848) );
  INVX1 U2380 ( .A(SHA256_result[148]), .Y(n875) );
  INVX1 U2381 ( .A(SHA256_result[63]), .Y(n950) );
  INVX1 U2382 ( .A(SHA256_result[61]), .Y(n948) );
  INVX1 U2383 ( .A(SHA256_result[60]), .Y(n947) );
  INVX1 U2384 ( .A(SHA256_result[59]), .Y(n946) );
  INVX1 U2385 ( .A(SHA256_result[57]), .Y(n944) );
  INVX1 U2386 ( .A(SHA256_result[56]), .Y(n943) );
  INVX1 U2387 ( .A(SHA256_result[94]), .Y(n924) );
  INVX1 U2388 ( .A(SHA256_result[93]), .Y(n923) );
  INVX1 U2389 ( .A(SHA256_result[88]), .Y(n918) );
  INVX1 U2390 ( .A(SHA256_result[149]), .Y(n876) );
  INVX1 U2391 ( .A(SHA256_result[151]), .Y(n878) );
  INVX1 U2392 ( .A(SHA256_result[135]), .Y(n862) );
  INVX1 U2393 ( .A(SHA256_result[134]), .Y(n861) );
  INVX1 U2394 ( .A(SHA256_result[29]), .Y(n981) );
  INVX1 U2395 ( .A(SHA256_result[26]), .Y(n978) );
  INVX1 U2396 ( .A(SHA256_result[158]), .Y(n885) );
  INVX1 U2397 ( .A(SHA256_result[31]), .Y(n951) );
  INVX1 U2398 ( .A(SHA256_result[153]), .Y(n880) );
  INVX1 U2399 ( .A(SHA256_result[139]), .Y(n866) );
  INVX1 U2400 ( .A(SHA256_result[137]), .Y(n864) );
  INVX1 U2401 ( .A(SHA256_result[217]), .Y(n820) );
  INVX1 U2402 ( .A(SHA256_result[216]), .Y(n819) );
  INVXL U2403 ( .A(SHA256_result[99]), .Y(n533) );
  INVX1 U2404 ( .A(SHA256_result[154]), .Y(n881) );
  INVX1 U2405 ( .A(SHA256_result[223]), .Y(n794) );
  INVX1 U2406 ( .A(SHA256_result[181]), .Y(n843) );
  INVX1 U2407 ( .A(SHA256_result[188]), .Y(n850) );
  INVX1 U2408 ( .A(SHA256_result[187]), .Y(n849) );
  INVX1 U2409 ( .A(SHA256_result[143]), .Y(n870) );
  INVX1 U2410 ( .A(SHA256_result[92]), .Y(n922) );
  INVX1 U2411 ( .A(SHA256_result[91]), .Y(n921) );
  INVX1 U2412 ( .A(SHA256_result[89]), .Y(n919) );
  INVX1 U2413 ( .A(SHA256_result[58]), .Y(n945) );
  INVX1 U2414 ( .A(SHA256_result[152]), .Y(n879) );
  INVX1 U2415 ( .A(SHA256_result[150]), .Y(n877) );
  INVX1 U2416 ( .A(SHA256_result[145]), .Y(n872) );
  INVX1 U2417 ( .A(SHA256_result[144]), .Y(n871) );
  INVX1 U2418 ( .A(SHA256_result[133]), .Y(n860) );
  INVX1 U2419 ( .A(SHA256_result[132]), .Y(n859) );
  INVX1 U2420 ( .A(SHA256_result[30]), .Y(n982) );
  INVX1 U2421 ( .A(SHA256_result[28]), .Y(n980) );
  INVX1 U2422 ( .A(SHA256_result[27]), .Y(n979) );
  INVX1 U2423 ( .A(SHA256_result[25]), .Y(n977) );
  INVX1 U2424 ( .A(SHA256_result[24]), .Y(n976) );
  INVX1 U2425 ( .A(SHA256_result[157]), .Y(n884) );
  INVX1 U2426 ( .A(SHA256_result[142]), .Y(n869) );
  INVX1 U2427 ( .A(SHA256_result[140]), .Y(n867) );
  INVX1 U2428 ( .A(SHA256_result[138]), .Y(n865) );
  INVX1 U2429 ( .A(SHA256_result[136]), .Y(n863) );
  INVX1 U2430 ( .A(SHA256_result[159]), .Y(n854) );
  INVX1 U2431 ( .A(SHA256_result[147]), .Y(n874) );
  INVX1 U2432 ( .A(SHA256_result[146]), .Y(n873) );
  INVX1 U2433 ( .A(SHA256_result[141]), .Y(n868) );
  AOI21XL U2434 ( .A0(next_A[28]), .A1(n353), .B0(n618), .Y(n619) );
  AOI21XL U2435 ( .A0(next_E[25]), .A1(n281), .B0(n465), .Y(n466) );
  NAND2XL U2436 ( .A(next_E[28]), .B(n281), .Y(n453) );
  AOI21XL U2437 ( .A0(next_E[23]), .A1(n280), .B0(n470), .Y(n471) );
  AOI21XL U2438 ( .A0(next_E[29]), .A1(n289), .B0(n449), .Y(n450) );
  NAND2XL U2439 ( .A(next_A[29]), .B(n280), .Y(n616) );
  AOI21XL U2440 ( .A0(next_A[23]), .A1(n290), .B0(n637), .Y(n638) );
  AOI2BB2XL U2441 ( .B0(n189), .B1(n147), .A0N(n292), .A1N(n489), .Y(n490) );
  OAI2BB1X1 U2442 ( .A0N(N962), .A1N(n241), .B0(n490), .Y(n2796) );
  INVXL U2443 ( .A(next_A[13]), .Y(n665) );
  INVXL U2444 ( .A(next_E[15]), .Y(n489) );
  INVXL U2445 ( .A(next_A[15]), .Y(n659) );
  AOI21XL U2446 ( .A0(next_E[26]), .A1(n285), .B0(n461), .Y(n462) );
  NAND2XL U2447 ( .A(next_A[27]), .B(n341), .Y(n621) );
  AOI21XL U2448 ( .A0(next_A[26]), .A1(n288), .B0(n625), .Y(n626) );
  NAND2XL U2449 ( .A(next_A[25]), .B(n282), .Y(n629) );
  XOR3X4 U2450 ( .A(n150), .B(SHA256_result[110]), .C(SHA256_result[124]), .Y(
        f4_E_32[3]) );
  NOR2X1 U2451 ( .A(read_counter[1]), .B(read_counter[0]), .Y(n737) );
  AOI21X1 U2452 ( .A0(read_counter[0]), .A1(read_counter[1]), .B0(n737), .Y(
        n736) );
  INVX1 U2453 ( .A(n736), .Y(N3180) );
  NAND2X1 U2454 ( .A(n737), .B(n985), .Y(n738) );
  OAI21XL U2455 ( .A0(n737), .A1(n985), .B0(n738), .Y(N3181) );
  XNOR2X1 U2456 ( .A(read_counter[3]), .B(n738), .Y(N3182) );
  NOR2X1 U2457 ( .A(read_counter[3]), .B(n738), .Y(n739) );
  XOR2X1 U2458 ( .A(read_counter[4]), .B(n739), .Y(N3183) );
endmodule


module controller_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module controller ( clk, reset, first_block, last_block, output_enable, busy, 
        inner_busy );
  input clk, reset, first_block, last_block;
  output output_enable, busy, inner_busy;
  wire   N10, N11, N24, N25, N26, N27, N28, N29, N30, N45, N46, N47, N48, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n1, n13, n14, n15, n16;
  wire   [1:0] state;
  wire   [6:0] counter1;
  wire   [4:0] counter2;
  wire   [4:2] add_93_carry;

  AND2X2 U10 ( .A(counter2[1]), .B(counter2[0]), .Y(n23) );
  controller_DW01_inc_1 add_82 ( .A(counter1), .SUM({N30, N29, N28, N27, N26, 
        N25, N24}) );
  DFFTRX1 counter2_reg_4_ ( .D(N48), .RN(n15), .CK(clk), .Q(counter2[4]) );
  DFFTRX1 counter2_reg_3_ ( .D(N47), .RN(n15), .CK(clk), .Q(counter2[3]) );
  DFFTRX1 counter2_reg_2_ ( .D(N46), .RN(n15), .CK(clk), .Q(counter2[2]) );
  DFFTRX1 counter1_reg_6_ ( .D(N30), .RN(n19), .CK(clk), .Q(counter1[6]) );
  DFFTRX1 counter2_reg_1_ ( .D(N45), .RN(n15), .CK(clk), .Q(counter2[1]) );
  DFFTRX1 counter2_reg_0_ ( .D(n1), .RN(n15), .CK(clk), .Q(counter2[0]), .QN(
        n1) );
  DFFTRX1 counter1_reg_5_ ( .D(N29), .RN(n19), .CK(clk), .Q(counter1[5]) );
  DFFTRX1 counter1_reg_4_ ( .D(N28), .RN(n19), .CK(clk), .Q(counter1[4]) );
  DFFTRX1 counter1_reg_3_ ( .D(N27), .RN(n19), .CK(clk), .Q(counter1[3]) );
  DFFTRX1 counter1_reg_2_ ( .D(N26), .RN(n19), .CK(clk), .Q(counter1[2]) );
  DFFTRX1 counter1_reg_1_ ( .D(N25), .RN(n19), .CK(clk), .Q(counter1[1]) );
  DFFTRX1 counter1_reg_0_ ( .D(N24), .RN(n19), .CK(clk), .Q(counter1[0]) );
  DFFHQX1 state_reg_0_ ( .D(N10), .CK(clk), .Q(state[0]) );
  DFFHQX1 state_reg_1_ ( .D(N11), .CK(clk), .Q(state[1]) );
  NOR2BX2 U3 ( .AN(state[1]), .B(state[0]), .Y(output_enable) );
  NOR2BX1 U4 ( .AN(state[0]), .B(state[1]), .Y(inner_busy) );
  NOR2XL U5 ( .A(state[1]), .B(state[0]), .Y(n17) );
  AOI22XL U6 ( .A0(first_block), .A1(n17), .B0(inner_busy), .B1(n21), .Y(n24)
         );
  INVXL U7 ( .A(inner_busy), .Y(n14) );
  NAND2BXL U8 ( .AN(reset), .B(output_enable), .Y(n18) );
  INVX1 U9 ( .A(n17), .Y(busy) );
  INVX1 U11 ( .A(n18), .Y(n15) );
  AOI211X1 U12 ( .A0(n16), .A1(n20), .B0(n13), .C0(reset), .Y(n19) );
  INVX1 U13 ( .A(n21), .Y(n13) );
  INVX1 U14 ( .A(last_block), .Y(n16) );
  NOR2X1 U15 ( .A(reset), .B(n24), .Y(N10) );
  OAI32X1 U16 ( .A0(n14), .A1(reset), .A2(n21), .B0(n22), .B1(n18), .Y(N11) );
  AND4X2 U17 ( .A(counter2[4]), .B(counter2[3]), .C(n23), .D(counter2[2]), .Y(
        n22) );
  NAND2X1 U18 ( .A(counter1[6]), .B(n20), .Y(n21) );
  ADDHXL U19 ( .A(counter2[1]), .B(counter2[0]), .CO(add_93_carry[2]), .S(N45)
         );
  ADDHXL U20 ( .A(counter2[2]), .B(add_93_carry[2]), .CO(add_93_carry[3]), .S(
        N46) );
  ADDHXL U21 ( .A(counter2[3]), .B(add_93_carry[3]), .CO(add_93_carry[4]), .S(
        N47) );
  NOR4X1 U22 ( .A(counter1[2]), .B(counter1[1]), .C(counter1[0]), .D(n25), .Y(
        n20) );
  OR3XL U23 ( .A(counter1[5]), .B(counter1[4]), .C(counter1[3]), .Y(n25) );
  XOR2X1 U24 ( .A(add_93_carry[4]), .B(counter2[4]), .Y(N48) );
endmodule


module top ( clk, reset, data, write_enable, last_block, first_block, busy, 
        digest, output_enable );
  input [31:0] data;
  output [7:0] digest;
  input clk, reset, write_enable, last_block, first_block;
  output busy, output_enable;
  wire   inner_busy;
  wire   [31:0] Wt;

  message_schedule our_message_schedule ( .clk(clk), .reset(reset), .data(data), .write_enable(write_enable), .inner_busy(inner_busy), .Wt(Wt) );
  hash_core our_hash_core ( .clk(clk), .reset(reset), .Wt(Wt), .inner_busy(
        inner_busy), .first_block(first_block), .output_enable(output_enable), 
        .digest(digest) );
  controller our_controller ( .clk(clk), .reset(reset), .first_block(
        first_block), .last_block(last_block), .output_enable(output_enable), 
        .busy(busy), .inner_busy(inner_busy) );
endmodule


module sha256_chip ( clk, reset, data, write_enable, last_block, first_block, 
        busy, digest, output_enable );
  input [31:0] data;
  output [7:0] digest;
  input clk, reset, write_enable, last_block, first_block;
  output busy, output_enable;
  wire   net_clk, net_reset, net_write_enable, net_last_block, net_first_block,
         net_busy, net_output_enable;
  wire   [31:0] net_data;
  wire   [7:0] net_digest;

  PIW PIW_clk ( .PAD(clk), .C(net_clk) );
  PIW PIW_reset ( .PAD(reset), .C(net_reset) );
  PIW PIW_data0 ( .PAD(data[0]), .C(net_data[0]) );
  PIW PIW_data1 ( .PAD(data[1]), .C(net_data[1]) );
  PIW PIW_data2 ( .PAD(data[2]), .C(net_data[2]) );
  PIW PIW_data3 ( .PAD(data[3]), .C(net_data[3]) );
  PIW PIW_data4 ( .PAD(data[4]), .C(net_data[4]) );
  PIW PIW_data5 ( .PAD(data[5]), .C(net_data[5]) );
  PIW PIW_data6 ( .PAD(data[6]), .C(net_data[6]) );
  PIW PIW_data7 ( .PAD(data[7]), .C(net_data[7]) );
  PIW PIW_data8 ( .PAD(data[8]), .C(net_data[8]) );
  PIW PIW_data9 ( .PAD(data[9]), .C(net_data[9]) );
  PIW PIW_data10 ( .PAD(data[10]), .C(net_data[10]) );
  PIW PIW_data11 ( .PAD(data[11]), .C(net_data[11]) );
  PIW PIW_data12 ( .PAD(data[12]), .C(net_data[12]) );
  PIW PIW_data13 ( .PAD(data[13]), .C(net_data[13]) );
  PIW PIW_data14 ( .PAD(data[14]), .C(net_data[14]) );
  PIW PIW_data15 ( .PAD(data[15]), .C(net_data[15]) );
  PIW PIW_data16 ( .PAD(data[16]), .C(net_data[16]) );
  PIW PIW_data17 ( .PAD(data[17]), .C(net_data[17]) );
  PIW PIW_data18 ( .PAD(data[18]), .C(net_data[18]) );
  PIW PIW_data19 ( .PAD(data[19]), .C(net_data[19]) );
  PIW PIW_data20 ( .PAD(data[20]), .C(net_data[20]) );
  PIW PIW_data21 ( .PAD(data[21]), .C(net_data[21]) );
  PIW PIW_data22 ( .PAD(data[22]), .C(net_data[22]) );
  PIW PIW_data23 ( .PAD(data[23]), .C(net_data[23]) );
  PIW PIW_data24 ( .PAD(data[24]), .C(net_data[24]) );
  PIW PIW_data25 ( .PAD(data[25]), .C(net_data[25]) );
  PIW PIW_data26 ( .PAD(data[26]), .C(net_data[26]) );
  PIW PIW_data27 ( .PAD(data[27]), .C(net_data[27]) );
  PIW PIW_data28 ( .PAD(data[28]), .C(net_data[28]) );
  PIW PIW_data29 ( .PAD(data[29]), .C(net_data[29]) );
  PIW PIW_data30 ( .PAD(data[30]), .C(net_data[30]) );
  PIW PIW_data31 ( .PAD(data[31]), .C(net_data[31]) );
  PIW PIW_write_enable ( .PAD(write_enable), .C(net_write_enable) );
  PIW PIW_last_block ( .PAD(last_block), .C(net_last_block) );
  PIW PIW_first_block ( .PAD(first_block), .C(net_first_block) );
  PO8W PO8W_busy ( .I(net_busy), .PAD(busy) );
  PO8W PO8W_digest0 ( .I(net_digest[0]), .PAD(digest[0]) );
  PO8W PO8W_digest1 ( .I(net_digest[1]), .PAD(digest[1]) );
  PO8W PO8W_digest2 ( .I(net_digest[2]), .PAD(digest[2]) );
  PO8W PO8W_digest3 ( .I(net_digest[3]), .PAD(digest[3]) );
  PO8W PO8W_digest4 ( .I(net_digest[4]), .PAD(digest[4]) );
  PO8W PO8W_digest5 ( .I(net_digest[5]), .PAD(digest[5]) );
  PO8W PO8W_digest6 ( .I(net_digest[6]), .PAD(digest[6]) );
  PO8W PO8W_digest7 ( .I(net_digest[7]), .PAD(digest[7]) );
  PO8W PO8W_output_enable ( .I(net_output_enable), .PAD(output_enable) );
  top inst_top ( .clk(net_clk), .reset(net_reset), .data(net_data), 
        .write_enable(net_write_enable), .last_block(net_last_block), 
        .first_block(net_first_block), .busy(net_busy), .digest(net_digest), 
        .output_enable(net_output_enable) );
endmodule


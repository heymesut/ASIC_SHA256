
module message_schedule_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module message_schedule_DW01_add_2 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1;
  wire   [31:1] carry;

  ADDFHX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX4 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX4 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX4 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX4 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX4 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFHX4 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX4 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX4 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  INVX4 U1 ( .A(n1), .Y(carry[1]) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND2X4 U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
endmodule


module message_schedule_DW01_add_6 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224;

  NOR2X2 U2 ( .A(n58), .B(n60), .Y(n219) );
  OR2X4 U3 ( .A(n193), .B(n170), .Y(n1) );
  NAND2X1 U4 ( .A(n1), .B(n171), .Y(n191) );
  NAND2XL U5 ( .A(n208), .B(n3), .Y(n4) );
  NAND2X1 U6 ( .A(n2), .B(n209), .Y(n5) );
  NAND2X2 U7 ( .A(n4), .B(n5), .Y(SUM[10]) );
  INVXL U8 ( .A(n208), .Y(n2) );
  INVX1 U9 ( .A(n209), .Y(n3) );
  OAI21X4 U10 ( .A0(n17), .A1(n210), .B0(n29), .Y(n208) );
  NAND2X2 U11 ( .A(n205), .B(n7), .Y(n8) );
  NAND2X2 U12 ( .A(n6), .B(n206), .Y(n9) );
  NAND2X4 U13 ( .A(n8), .B(n9), .Y(SUM[11]) );
  INVX2 U14 ( .A(n205), .Y(n6) );
  INVXL U15 ( .A(n206), .Y(n7) );
  XOR2X2 U16 ( .A(n65), .B(n15), .Y(SUM[30]) );
  NAND2X1 U17 ( .A(n10), .B(n128), .Y(n107) );
  OAI21X2 U18 ( .A0(n169), .A1(n14), .B0(n158), .Y(n154) );
  INVX1 U19 ( .A(n159), .Y(n158) );
  OAI21XL U20 ( .A0(n160), .A1(n22), .B0(n161), .Y(n159) );
  OAI21XL U21 ( .A0(n18), .A1(n166), .B0(n167), .Y(n163) );
  OAI21XL U22 ( .A0(n213), .A1(n214), .B0(n35), .Y(n174) );
  INVX2 U23 ( .A(n30), .Y(n193) );
  NAND2X1 U24 ( .A(n103), .B(n104), .Y(n83) );
  OR2X2 U25 ( .A(A[5]), .B(B[5]), .Y(n45) );
  NAND2X1 U26 ( .A(B[4]), .B(A[4]), .Y(n48) );
  NOR2X1 U27 ( .A(A[9]), .B(B[9]), .Y(n17) );
  INVX1 U28 ( .A(n198), .Y(n203) );
  INVX1 U29 ( .A(n188), .Y(n187) );
  NAND2X1 U30 ( .A(n151), .B(n141), .Y(n149) );
  BUFX3 U31 ( .A(n127), .Y(n10) );
  OAI21XL U32 ( .A0(n131), .A1(n132), .B0(n133), .Y(n127) );
  NAND2X1 U33 ( .A(n124), .B(n119), .Y(n122) );
  NAND2X4 U34 ( .A(n154), .B(n155), .Y(n131) );
  OAI21X4 U35 ( .A0(n19), .A1(n193), .B0(n32), .Y(n27) );
  NOR2XL U36 ( .A(n49), .B(n54), .Y(n223) );
  NAND2XL U37 ( .A(B[9]), .B(A[9]), .Y(n29) );
  OR2XL U38 ( .A(A[4]), .B(B[4]), .Y(n46) );
  OR2X1 U39 ( .A(A[6]), .B(B[6]), .Y(n215) );
  XOR2X1 U40 ( .A(n76), .B(n68), .Y(SUM[29]) );
  OR2X1 U41 ( .A(A[1]), .B(B[1]), .Y(n73) );
  OAI21X1 U42 ( .A0(n67), .A1(n68), .B0(n69), .Y(n65) );
  NOR2BXL U43 ( .AN(n57), .B(n58), .Y(n56) );
  NAND2X1 U44 ( .A(B[1]), .B(A[1]), .Y(n74) );
  NAND2X1 U45 ( .A(B[6]), .B(A[6]), .Y(n39) );
  NAND2XL U46 ( .A(B[2]), .B(A[2]), .Y(n61) );
  OAI21XL U47 ( .A0(n148), .A1(n137), .B0(n136), .Y(n146) );
  OAI21XL U48 ( .A0(n59), .A1(n60), .B0(n61), .Y(n55) );
  NOR2XL U49 ( .A(n48), .B(n49), .Y(n42) );
  INVX1 U50 ( .A(n165), .Y(n164) );
  XOR2X1 U51 ( .A(n122), .B(n16), .Y(SUM[22]) );
  NOR2X1 U52 ( .A(A[13]), .B(B[13]), .Y(n18) );
  NAND2XL U53 ( .A(B[5]), .B(A[5]), .Y(n43) );
  NAND2X1 U54 ( .A(B[8]), .B(A[8]), .Y(n32) );
  OAI2BB1X2 U55 ( .A0N(n211), .A1N(n47), .B0(n212), .Y(n30) );
  CLKINVX3 U56 ( .A(n168), .Y(n211) );
  OAI21X2 U57 ( .A0(n21), .A1(n190), .B0(n166), .Y(n188) );
  INVX2 U58 ( .A(n191), .Y(n190) );
  INVX2 U59 ( .A(n27), .Y(n210) );
  OAI21X2 U60 ( .A0(n187), .A1(n18), .B0(n167), .Y(n185) );
  NAND2XL U61 ( .A(n215), .B(n216), .Y(n214) );
  NAND3BX2 U62 ( .AN(n179), .B(n57), .C(n177), .Y(n47) );
  NOR2BXL U63 ( .AN(n165), .B(n182), .Y(n186) );
  XOR2X2 U64 ( .A(n183), .B(n184), .Y(SUM[15]) );
  NOR2BXL U65 ( .AN(n161), .B(n22), .Y(n184) );
  INVXL U66 ( .A(n221), .Y(n58) );
  NOR2BX1 U67 ( .AN(n142), .B(n134), .Y(n133) );
  XNOR2X1 U68 ( .A(n98), .B(n11), .Y(SUM[26]) );
  NAND2X1 U69 ( .A(n91), .B(n86), .Y(n11) );
  NOR2BXL U70 ( .AN(n48), .B(n54), .Y(n53) );
  NOR2BXL U71 ( .AN(n39), .B(n38), .Y(n41) );
  NOR2BXL U72 ( .AN(n141), .B(n139), .Y(n153) );
  NOR2BXL U73 ( .AN(n32), .B(n19), .Y(n31) );
  INVXL U74 ( .A(n170), .Y(n175) );
  AOI21XL U75 ( .A0(n176), .A1(n177), .B0(n168), .Y(n173) );
  NOR2XL U76 ( .A(n178), .B(n179), .Y(n176) );
  NAND3XL U77 ( .A(n45), .B(n46), .C(n47), .Y(n44) );
  XNOR2X1 U78 ( .A(n103), .B(n12), .Y(SUM[24]) );
  NAND2X1 U79 ( .A(n94), .B(n104), .Y(n12) );
  XNOR2X1 U80 ( .A(n77), .B(n13), .Y(SUM[28]) );
  NAND2X1 U81 ( .A(n80), .B(n78), .Y(n13) );
  NAND2XL U82 ( .A(n61), .B(n75), .Y(n71) );
  NAND2XL U83 ( .A(n65), .B(n66), .Y(n64) );
  NAND2XL U84 ( .A(B[3]), .B(A[3]), .Y(n57) );
  NAND2XL U85 ( .A(B[7]), .B(A[7]), .Y(n35) );
  NAND2XL U86 ( .A(B[10]), .B(A[10]), .Y(n200) );
  NAND2XL U87 ( .A(B[11]), .B(A[11]), .Y(n197) );
  NOR2XL U88 ( .A(A[0]), .B(B[0]), .Y(n24) );
  AND2X1 U89 ( .A(B[0]), .B(A[0]), .Y(n25) );
  NOR2XL U90 ( .A(A[12]), .B(B[12]), .Y(n21) );
  NAND2XL U91 ( .A(B[0]), .B(A[0]), .Y(n26) );
  NAND2XL U92 ( .A(B[17]), .B(A[17]), .Y(n141) );
  NAND2XL U93 ( .A(B[13]), .B(A[13]), .Y(n167) );
  NAND2XL U94 ( .A(B[15]), .B(A[15]), .Y(n161) );
  NAND3XL U95 ( .A(A[0]), .B(B[0]), .C(n73), .Y(n72) );
  AND2X1 U96 ( .A(n74), .B(n72), .Y(n59) );
  AND2X2 U97 ( .A(n171), .B(n172), .Y(n14) );
  INVX1 U98 ( .A(n174), .Y(n212) );
  NAND2X1 U99 ( .A(n223), .B(n224), .Y(n168) );
  NOR2X1 U100 ( .A(n36), .B(n38), .Y(n224) );
  INVX1 U101 ( .A(n45), .Y(n49) );
  INVX1 U102 ( .A(n215), .Y(n38) );
  NAND3BX1 U103 ( .AN(n20), .B(n143), .C(n144), .Y(n132) );
  AOI21X1 U104 ( .A0(n194), .A1(n195), .B0(n196), .Y(n171) );
  INVX1 U105 ( .A(n197), .Y(n196) );
  OAI2BB1X1 U106 ( .A0N(n198), .A1N(n199), .B0(n200), .Y(n195) );
  OAI21XL U107 ( .A0(n17), .A1(n32), .B0(n29), .Y(n199) );
  NOR2X1 U108 ( .A(n217), .B(n218), .Y(n213) );
  NAND2X1 U109 ( .A(n39), .B(n43), .Y(n218) );
  INVX1 U110 ( .A(n46), .Y(n54) );
  INVX1 U111 ( .A(n75), .Y(n60) );
  INVX1 U112 ( .A(n216), .Y(n36) );
  NOR2BX1 U113 ( .AN(n200), .B(n203), .Y(n209) );
  XOR2X1 U114 ( .A(n27), .B(n28), .Y(SUM[9]) );
  NOR2BX1 U115 ( .AN(n29), .B(n17), .Y(n28) );
  XOR2X1 U116 ( .A(n188), .B(n189), .Y(SUM[13]) );
  NOR2BX1 U117 ( .AN(n167), .B(n18), .Y(n189) );
  XOR2X1 U118 ( .A(n185), .B(n186), .Y(SUM[14]) );
  XOR2X1 U119 ( .A(n33), .B(n34), .Y(SUM[7]) );
  NOR2BX1 U120 ( .AN(n35), .B(n36), .Y(n34) );
  OAI21XL U121 ( .A0(n37), .A1(n38), .B0(n39), .Y(n33) );
  INVX1 U122 ( .A(n40), .Y(n37) );
  NOR2BX1 U123 ( .AN(n197), .B(n204), .Y(n206) );
  OAI21XL U124 ( .A0(n207), .A1(n203), .B0(n200), .Y(n205) );
  INVX1 U125 ( .A(n208), .Y(n207) );
  XOR2X1 U126 ( .A(n146), .B(n147), .Y(SUM[19]) );
  NOR2BX1 U127 ( .AN(n142), .B(n20), .Y(n147) );
  INVX1 U128 ( .A(n149), .Y(n148) );
  OAI2BB1X1 U129 ( .A0N(n162), .A1N(n185), .B0(n165), .Y(n183) );
  NAND2X1 U130 ( .A(n83), .B(n94), .Y(n101) );
  NAND2X1 U131 ( .A(n131), .B(n140), .Y(n152) );
  OAI21XL U132 ( .A0(n173), .A1(n174), .B0(n175), .Y(n172) );
  NAND3BX1 U133 ( .AN(n42), .B(n43), .C(n44), .Y(n40) );
  NAND2X1 U134 ( .A(n100), .B(n95), .Y(n98) );
  NAND2X1 U135 ( .A(n84), .B(n101), .Y(n100) );
  NAND2X1 U136 ( .A(n105), .B(n106), .Y(n103) );
  AOI21X1 U137 ( .A0(n111), .A1(n109), .B0(n112), .Y(n105) );
  NAND4BXL U138 ( .AN(n107), .B(n108), .C(n109), .D(n110), .Y(n106) );
  INVX1 U139 ( .A(n113), .Y(n112) );
  NOR2X1 U140 ( .A(n49), .B(n48), .Y(n217) );
  NAND2X1 U141 ( .A(n201), .B(n202), .Y(n170) );
  NOR2X1 U142 ( .A(n203), .B(n204), .Y(n201) );
  NOR2X1 U143 ( .A(n19), .B(n17), .Y(n202) );
  INVX1 U144 ( .A(n222), .Y(n179) );
  NAND2BX1 U145 ( .AN(n61), .B(n221), .Y(n222) );
  NAND2X1 U146 ( .A(n144), .B(n152), .Y(n151) );
  AND2X2 U147 ( .A(n63), .B(n66), .Y(n15) );
  AOI21X1 U148 ( .A0(n77), .A1(n78), .B0(n79), .Y(n68) );
  INVX1 U149 ( .A(n80), .Y(n79) );
  INVX1 U150 ( .A(n70), .Y(n67) );
  INVX1 U151 ( .A(n143), .Y(n137) );
  XOR2X1 U152 ( .A(n101), .B(n102), .Y(SUM[25]) );
  NOR2BX1 U153 ( .AN(n95), .B(n93), .Y(n102) );
  NAND2X1 U154 ( .A(n69), .B(n70), .Y(n76) );
  XOR2X1 U155 ( .A(n50), .B(n51), .Y(SUM[5]) );
  NAND2X1 U156 ( .A(n45), .B(n43), .Y(n50) );
  AOI21X1 U157 ( .A0(n47), .A1(n46), .B0(n52), .Y(n51) );
  INVX1 U158 ( .A(n48), .Y(n52) );
  INVX1 U159 ( .A(n144), .Y(n139) );
  INVX1 U160 ( .A(n162), .Y(n182) );
  INVX1 U161 ( .A(n194), .Y(n204) );
  XOR2X1 U162 ( .A(n55), .B(n56), .Y(SUM[3]) );
  XOR2X1 U163 ( .A(n47), .B(n53), .Y(SUM[4]) );
  AOI21X1 U164 ( .A0(n135), .A1(n136), .B0(n20), .Y(n134) );
  NAND2BX1 U165 ( .AN(n137), .B(n138), .Y(n135) );
  OAI21XL U166 ( .A0(n139), .A1(n140), .B0(n141), .Y(n138) );
  XOR2X1 U167 ( .A(n10), .B(n129), .Y(SUM[20]) );
  NOR2BX1 U168 ( .AN(n118), .B(n130), .Y(n129) );
  INVX1 U169 ( .A(n128), .Y(n130) );
  XOR2X1 U170 ( .A(n191), .B(n192), .Y(SUM[12]) );
  NOR2BX1 U171 ( .AN(n166), .B(n21), .Y(n192) );
  XOR2X1 U172 ( .A(n40), .B(n41), .Y(SUM[6]) );
  XOR2X1 U173 ( .A(n152), .B(n153), .Y(SUM[17]) );
  XOR2X1 U174 ( .A(n125), .B(n126), .Y(SUM[21]) );
  NOR2BX1 U175 ( .AN(n119), .B(n117), .Y(n126) );
  XOR2X1 U176 ( .A(n71), .B(n59), .Y(SUM[2]) );
  XOR2X1 U177 ( .A(n120), .B(n121), .Y(SUM[23]) );
  NAND2X1 U178 ( .A(n113), .B(n109), .Y(n120) );
  AOI21X1 U179 ( .A0(n110), .A1(n122), .B0(n123), .Y(n121) );
  INVX1 U180 ( .A(n115), .Y(n123) );
  XOR2X1 U181 ( .A(n96), .B(n97), .Y(SUM[27]) );
  NAND2X1 U182 ( .A(n89), .B(n85), .Y(n96) );
  AOI21X1 U183 ( .A0(n86), .A1(n98), .B0(n99), .Y(n97) );
  INVX1 U184 ( .A(n91), .Y(n99) );
  XOR2X1 U185 ( .A(n30), .B(n31), .Y(SUM[8]) );
  XOR2X1 U186 ( .A(n149), .B(n150), .Y(SUM[18]) );
  NOR2BX1 U187 ( .AN(n136), .B(n137), .Y(n150) );
  XOR2X1 U188 ( .A(n154), .B(n156), .Y(SUM[16]) );
  NOR2BX1 U189 ( .AN(n140), .B(n157), .Y(n156) );
  INVX1 U190 ( .A(n155), .Y(n157) );
  AND2X2 U191 ( .A(n115), .B(n110), .Y(n16) );
  NAND2X1 U192 ( .A(n107), .B(n118), .Y(n125) );
  AOI21X1 U193 ( .A0(n162), .A1(n163), .B0(n164), .Y(n160) );
  NAND2X1 U194 ( .A(n108), .B(n125), .Y(n124) );
  NAND2X1 U195 ( .A(n81), .B(n82), .Y(n77) );
  AOI21X1 U196 ( .A0(n87), .A1(n85), .B0(n88), .Y(n81) );
  NAND4BXL U197 ( .AN(n83), .B(n84), .C(n85), .D(n86), .Y(n82) );
  INVX1 U198 ( .A(n89), .Y(n88) );
  INVX1 U199 ( .A(n57), .Y(n178) );
  NAND2X1 U200 ( .A(n74), .B(n73), .Y(n145) );
  NAND2X1 U201 ( .A(n180), .B(n181), .Y(n169) );
  NOR2X1 U202 ( .A(n22), .B(n182), .Y(n181) );
  NOR2X1 U203 ( .A(n18), .B(n21), .Y(n180) );
  INVX1 U204 ( .A(n108), .Y(n117) );
  NAND2X1 U205 ( .A(n114), .B(n115), .Y(n111) );
  NAND2X1 U206 ( .A(n110), .B(n116), .Y(n114) );
  OAI21XL U207 ( .A0(n117), .A1(n118), .B0(n119), .Y(n116) );
  INVX1 U208 ( .A(n84), .Y(n93) );
  NAND2X1 U209 ( .A(n90), .B(n91), .Y(n87) );
  NAND2X1 U210 ( .A(n86), .B(n92), .Y(n90) );
  OAI21XL U211 ( .A0(n93), .A1(n94), .B0(n95), .Y(n92) );
  NAND3X1 U212 ( .A(n219), .B(n73), .C(n220), .Y(n177) );
  OAI2BB1X1 U213 ( .A0N(B[0]), .A1N(A[0]), .B0(n74), .Y(n220) );
  OR2X2 U214 ( .A(A[3]), .B(B[3]), .Y(n221) );
  OR2X2 U215 ( .A(A[2]), .B(B[2]), .Y(n75) );
  OR2X2 U216 ( .A(A[7]), .B(B[7]), .Y(n216) );
  OR2X2 U217 ( .A(A[10]), .B(B[10]), .Y(n198) );
  NOR2X1 U218 ( .A(A[8]), .B(B[8]), .Y(n19) );
  NOR2X1 U219 ( .A(A[19]), .B(B[19]), .Y(n20) );
  NAND2X1 U220 ( .A(B[16]), .B(A[16]), .Y(n140) );
  NAND2X1 U221 ( .A(B[12]), .B(A[12]), .Y(n166) );
  NAND2X1 U222 ( .A(B[14]), .B(A[14]), .Y(n165) );
  OR2X2 U223 ( .A(A[17]), .B(B[17]), .Y(n144) );
  OR2X2 U224 ( .A(A[14]), .B(B[14]), .Y(n162) );
  OR2X2 U225 ( .A(A[11]), .B(B[11]), .Y(n194) );
  OR2X2 U226 ( .A(A[18]), .B(B[18]), .Y(n143) );
  XOR2X1 U227 ( .A(n26), .B(n145), .Y(SUM[1]) );
  NOR2X1 U228 ( .A(A[15]), .B(B[15]), .Y(n22) );
  OR2X2 U229 ( .A(A[22]), .B(B[22]), .Y(n110) );
  NAND2X1 U230 ( .A(B[20]), .B(A[20]), .Y(n118) );
  NAND2X1 U231 ( .A(B[18]), .B(A[18]), .Y(n136) );
  NAND2X1 U232 ( .A(B[22]), .B(A[22]), .Y(n115) );
  OR2X2 U233 ( .A(A[23]), .B(B[23]), .Y(n109) );
  NAND2X1 U234 ( .A(B[21]), .B(A[21]), .Y(n119) );
  OR2X2 U235 ( .A(A[21]), .B(B[21]), .Y(n108) );
  NOR2X1 U236 ( .A(n24), .B(n25), .Y(SUM[0]) );
  NAND2X1 U237 ( .A(B[23]), .B(A[23]), .Y(n113) );
  OR2X2 U238 ( .A(A[24]), .B(B[24]), .Y(n104) );
  NAND2X1 U239 ( .A(B[19]), .B(A[19]), .Y(n142) );
  OR2X2 U240 ( .A(A[16]), .B(B[16]), .Y(n155) );
  OR2X2 U241 ( .A(A[20]), .B(B[20]), .Y(n128) );
  OR2X2 U242 ( .A(A[26]), .B(B[26]), .Y(n86) );
  NAND2X1 U243 ( .A(B[24]), .B(A[24]), .Y(n94) );
  NAND2X1 U244 ( .A(B[26]), .B(A[26]), .Y(n91) );
  OR2X2 U245 ( .A(A[27]), .B(B[27]), .Y(n85) );
  NAND2X1 U246 ( .A(B[25]), .B(A[25]), .Y(n95) );
  OR2X2 U247 ( .A(A[25]), .B(B[25]), .Y(n84) );
  NAND2X1 U248 ( .A(B[27]), .B(A[27]), .Y(n89) );
  NAND2X1 U249 ( .A(B[30]), .B(A[30]), .Y(n63) );
  NAND2X1 U250 ( .A(B[29]), .B(A[29]), .Y(n69) );
  NAND2X1 U251 ( .A(B[28]), .B(A[28]), .Y(n80) );
  OR2X2 U252 ( .A(A[28]), .B(B[28]), .Y(n78) );
  OR2X2 U253 ( .A(A[30]), .B(B[30]), .Y(n66) );
  OR2X2 U254 ( .A(A[29]), .B(B[29]), .Y(n70) );
  XOR3X2 U255 ( .A(B[31]), .B(A[31]), .C(n62), .Y(SUM[31]) );
  NAND2X1 U256 ( .A(n63), .B(n64), .Y(n62) );
endmodule


module message_schedule_DW01_add_8 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221;

  CLKINVX3 U2 ( .A(n216), .Y(n28) );
  INVX2 U3 ( .A(n189), .Y(n188) );
  OR2X4 U4 ( .A(A[28]), .B(B[28]), .Y(n74) );
  OR2X4 U5 ( .A(A[10]), .B(B[10]), .Y(n205) );
  OR2X4 U6 ( .A(A[11]), .B(B[11]), .Y(n200) );
  NAND2X2 U7 ( .A(B[30]), .B(A[30]), .Y(n56) );
  OAI21X2 U8 ( .A0(n39), .A1(n179), .B0(n214), .Y(n21) );
  INVX2 U9 ( .A(n81), .Y(n80) );
  CLKINVX3 U10 ( .A(n79), .Y(n4) );
  OAI21XL U11 ( .A0(n175), .A1(n171), .B0(n176), .Y(n174) );
  INVX1 U12 ( .A(n210), .Y(n203) );
  INVX1 U13 ( .A(n181), .Y(n170) );
  INVX1 U14 ( .A(n74), .Y(n64) );
  NAND2X1 U15 ( .A(B[28]), .B(A[28]), .Y(n65) );
  OR2X2 U16 ( .A(A[27]), .B(B[27]), .Y(n88) );
  NOR2X2 U17 ( .A(n57), .B(n58), .Y(n51) );
  INVX1 U18 ( .A(n59), .Y(n57) );
  XNOR2X2 U19 ( .A(B[31]), .B(A[31]), .Y(n49) );
  INVX1 U20 ( .A(n178), .Y(n214) );
  OAI21XL U21 ( .A0(n188), .A1(n12), .B0(n167), .Y(n186) );
  OAI211X1 U22 ( .A0(n82), .A1(n83), .B0(n84), .C0(n85), .Y(n79) );
  OR2X2 U23 ( .A(A[25]), .B(B[25]), .Y(n96) );
  NOR2X1 U24 ( .A(A[25]), .B(B[25]), .Y(n82) );
  INVX4 U25 ( .A(n66), .Y(n3) );
  OR2X2 U26 ( .A(n2), .B(n86), .Y(n1) );
  NOR2X4 U27 ( .A(A[27]), .B(B[27]), .Y(n2) );
  XOR2X1 U28 ( .A(n72), .B(n73), .Y(SUM[29]) );
  NOR2X4 U29 ( .A(A[30]), .B(B[30]), .Y(n58) );
  NAND2X1 U30 ( .A(B[27]), .B(A[27]), .Y(n81) );
  XNOR2X2 U31 ( .A(B[30]), .B(A[30]), .Y(n60) );
  NAND2X2 U32 ( .A(n95), .B(n84), .Y(n93) );
  NAND2X2 U33 ( .A(n96), .B(n97), .Y(n95) );
  INVX1 U34 ( .A(n93), .Y(n91) );
  NAND4BBX1 U35 ( .AN(n14), .BN(n15), .C(n34), .D(n216), .Y(n179) );
  OR2X4 U36 ( .A(A[7]), .B(B[7]), .Y(n216) );
  NAND3BX1 U37 ( .AN(n82), .B(n87), .C(n88), .Y(n77) );
  INVX1 U38 ( .A(n63), .Y(n62) );
  NAND2X1 U39 ( .A(B[29]), .B(A[29]), .Y(n63) );
  OAI21X4 U40 ( .A0(n54), .A1(n55), .B0(n56), .Y(n53) );
  AND2X4 U41 ( .A(n59), .B(n52), .Y(n6) );
  OAI2BB1X2 U42 ( .A0N(n66), .A1N(n74), .B0(n65), .Y(n10) );
  XOR2X4 U43 ( .A(n49), .B(n50), .Y(SUM[31]) );
  AOI21X4 U44 ( .A0(n51), .A1(n52), .B0(n53), .Y(n50) );
  NOR2X4 U45 ( .A(n1), .B(n4), .Y(n5) );
  NOR2X4 U46 ( .A(n5), .B(n80), .Y(n78) );
  NOR2X4 U47 ( .A(n6), .B(n62), .Y(n61) );
  XOR2X4 U48 ( .A(n61), .B(n60), .Y(SUM[30]) );
  NAND2X2 U49 ( .A(n7), .B(n8), .Y(n9) );
  NAND2X4 U50 ( .A(n9), .B(n106), .Y(n100) );
  CLKINVX2 U51 ( .A(n104), .Y(n7) );
  INVX1 U52 ( .A(n105), .Y(n8) );
  NAND2X2 U53 ( .A(n127), .B(n128), .Y(n104) );
  AOI21X2 U54 ( .A0(n107), .A1(n108), .B0(n109), .Y(n106) );
  NAND2X4 U55 ( .A(n100), .B(n101), .Y(n76) );
  OAI21X4 U56 ( .A0(n64), .A1(n3), .B0(n65), .Y(n52) );
  NAND2X1 U57 ( .A(n76), .B(n99), .Y(n97) );
  NAND2X1 U58 ( .A(B[9]), .B(A[9]), .Y(n20) );
  OAI21X4 U59 ( .A0(n76), .A1(n77), .B0(n78), .Y(n66) );
  OAI21XL U60 ( .A0(n197), .A1(n198), .B0(n199), .Y(n196) );
  INVX2 U61 ( .A(n10), .Y(n73) );
  NAND2X1 U62 ( .A(B[25]), .B(A[25]), .Y(n84) );
  NAND2X1 U63 ( .A(B[13]), .B(A[13]), .Y(n167) );
  NAND2X1 U64 ( .A(B[14]), .B(A[14]), .Y(n168) );
  NOR2X1 U65 ( .A(A[13]), .B(B[13]), .Y(n12) );
  NAND2X2 U66 ( .A(n160), .B(n161), .Y(n134) );
  OAI2BB1XL U67 ( .A0N(n195), .A1N(n21), .B0(n176), .Y(n193) );
  NAND3BXL U68 ( .AN(n111), .B(n117), .C(n118), .Y(n105) );
  OAI21X1 U69 ( .A0(n91), .A1(n86), .B0(n92), .Y(n89) );
  NAND4BBXL U70 ( .AN(n24), .BN(n13), .C(n205), .D(n200), .Y(n171) );
  NAND2XL U71 ( .A(n134), .B(n137), .Y(n158) );
  NAND2XL U72 ( .A(n104), .B(n112), .Y(n125) );
  NAND2XL U73 ( .A(n213), .B(n23), .Y(n18) );
  NAND2XL U74 ( .A(n21), .B(n206), .Y(n213) );
  AOI21XL U75 ( .A0(n205), .A1(n209), .B0(n203), .Y(n208) );
  NOR2BXL U76 ( .AN(n165), .B(n169), .Y(n184) );
  NAND2XL U77 ( .A(n137), .B(n138), .Y(n133) );
  NOR2BXL U78 ( .AN(n146), .B(n136), .Y(n154) );
  NOR2BXL U79 ( .AN(n168), .B(n170), .Y(n187) );
  NOR2BXL U80 ( .AN(n210), .B(n204), .Y(n211) );
  INVXL U81 ( .A(n180), .Y(n191) );
  NAND2XL U82 ( .A(n199), .B(n200), .Y(n207) );
  INVXL U83 ( .A(n101), .Y(n103) );
  NOR2BXL U84 ( .AN(n20), .B(n13), .Y(n19) );
  NOR2BXL U85 ( .AN(n145), .B(n143), .Y(n157) );
  NOR2BXL U86 ( .AN(n27), .B(n28), .Y(n26) );
  INVXL U87 ( .A(n128), .Y(n130) );
  AND2X1 U88 ( .A(n144), .B(n137), .Y(n159) );
  NOR2BXL U89 ( .AN(n36), .B(n14), .Y(n38) );
  INVXL U90 ( .A(n34), .Y(n30) );
  NOR2BXL U91 ( .AN(n44), .B(n16), .Y(n43) );
  NOR2BXL U92 ( .AN(n71), .B(n148), .Y(n147) );
  NAND2XL U93 ( .A(B[11]), .B(A[11]), .Y(n199) );
  NAND2XL U94 ( .A(B[15]), .B(A[15]), .Y(n165) );
  NAND2XL U95 ( .A(B[18]), .B(A[18]), .Y(n146) );
  NAND2XL U96 ( .A(B[22]), .B(A[22]), .Y(n114) );
  NAND2XL U97 ( .A(B[19]), .B(A[19]), .Y(n142) );
  NAND2XL U98 ( .A(B[23]), .B(A[23]), .Y(n110) );
  NAND2XL U99 ( .A(B[7]), .B(A[7]), .Y(n27) );
  NAND2XL U100 ( .A(B[24]), .B(A[24]), .Y(n99) );
  NAND2XL U101 ( .A(B[3]), .B(A[3]), .Y(n44) );
  OR2XL U102 ( .A(A[2]), .B(B[2]), .Y(n68) );
  NOR2BXL U103 ( .AN(n142), .B(n11), .Y(n151) );
  NOR2BXL U104 ( .AN(n84), .B(n82), .Y(n98) );
  NOR2BXL U105 ( .AN(n110), .B(n115), .Y(n120) );
  NOR2BXL U106 ( .AN(n114), .B(n116), .Y(n123) );
  NOR2BXL U107 ( .AN(n113), .B(n111), .Y(n126) );
  INVX1 U108 ( .A(n177), .Y(n39) );
  NOR2X1 U109 ( .A(n115), .B(n116), .Y(n107) );
  NAND2BX1 U110 ( .AN(n173), .B(n174), .Y(n160) );
  AOI21X1 U111 ( .A0(n162), .A1(n163), .B0(n164), .Y(n161) );
  NOR2X1 U112 ( .A(n169), .B(n170), .Y(n162) );
  AOI21X1 U113 ( .A0(n172), .A1(n177), .B0(n178), .Y(n175) );
  INVX1 U114 ( .A(n179), .Y(n172) );
  INVX1 U115 ( .A(n171), .Y(n195) );
  OAI211X1 U116 ( .A0(n111), .A1(n112), .B0(n113), .C0(n114), .Y(n108) );
  INVX1 U117 ( .A(n117), .Y(n116) );
  INVX1 U118 ( .A(n110), .Y(n109) );
  INVX1 U119 ( .A(n124), .Y(n111) );
  INVX1 U120 ( .A(n118), .Y(n115) );
  NAND2X1 U121 ( .A(n131), .B(n132), .Y(n127) );
  AOI21X1 U122 ( .A0(n139), .A1(n140), .B0(n141), .Y(n131) );
  NAND3BX1 U123 ( .AN(n133), .B(n134), .C(n135), .Y(n132) );
  INVX1 U124 ( .A(n142), .Y(n141) );
  NOR2X1 U125 ( .A(n11), .B(n136), .Y(n139) );
  NOR2X1 U126 ( .A(n136), .B(n11), .Y(n135) );
  OAI211X1 U127 ( .A0(n12), .A1(n166), .B0(n167), .C0(n168), .Y(n163) );
  OAI211X1 U128 ( .A0(n143), .A1(n144), .B0(n145), .C0(n146), .Y(n140) );
  INVX1 U129 ( .A(n152), .Y(n136) );
  INVX1 U130 ( .A(n138), .Y(n143) );
  INVX1 U131 ( .A(n182), .Y(n169) );
  OAI21XL U132 ( .A0(n121), .A1(n116), .B0(n114), .Y(n119) );
  INVX1 U133 ( .A(n122), .Y(n121) );
  OAI2BB1X1 U134 ( .A0N(n124), .A1N(n125), .B0(n113), .Y(n122) );
  NAND4BXL U135 ( .AN(n12), .B(n180), .C(n181), .D(n182), .Y(n173) );
  OAI21XL U136 ( .A0(n215), .A1(n28), .B0(n27), .Y(n178) );
  AOI21X1 U137 ( .A0(n34), .A1(n217), .B0(n218), .Y(n215) );
  INVX1 U138 ( .A(n31), .Y(n218) );
  OAI21XL U139 ( .A0(n14), .A1(n40), .B0(n36), .Y(n217) );
  OAI21XL U140 ( .A0(n155), .A1(n143), .B0(n145), .Y(n153) );
  INVX1 U141 ( .A(n156), .Y(n155) );
  INVX1 U142 ( .A(n205), .Y(n204) );
  INVX1 U143 ( .A(n196), .Y(n176) );
  INVX1 U144 ( .A(n200), .Y(n198) );
  AOI21X1 U145 ( .A0(n201), .A1(n202), .B0(n203), .Y(n197) );
  NOR2X1 U146 ( .A(n13), .B(n204), .Y(n201) );
  NAND2X1 U147 ( .A(n158), .B(n144), .Y(n156) );
  NAND2X1 U148 ( .A(n23), .B(n20), .Y(n202) );
  OAI2BB1X1 U149 ( .A0N(n152), .A1N(n153), .B0(n146), .Y(n150) );
  INVX1 U150 ( .A(n165), .Y(n164) );
  OAI21XL U151 ( .A0(n219), .A1(n16), .B0(n44), .Y(n177) );
  AOI21X1 U152 ( .A0(n68), .A1(n220), .B0(n221), .Y(n219) );
  INVX1 U153 ( .A(n47), .Y(n221) );
  OAI21XL U154 ( .A0(n148), .A1(n149), .B0(n71), .Y(n220) );
  OAI21XL U155 ( .A0(n191), .A1(n192), .B0(n166), .Y(n189) );
  INVX1 U156 ( .A(n193), .Y(n192) );
  INVX1 U157 ( .A(n69), .Y(n148) );
  OAI21XL U158 ( .A0(n185), .A1(n170), .B0(n168), .Y(n183) );
  INVX1 U159 ( .A(n186), .Y(n185) );
  INVX1 U160 ( .A(n206), .Y(n24) );
  OAI21XL U161 ( .A0(n212), .A1(n13), .B0(n20), .Y(n209) );
  INVX1 U162 ( .A(n18), .Y(n212) );
  OAI21XL U163 ( .A0(n35), .A1(n14), .B0(n36), .Y(n32) );
  INVX1 U164 ( .A(n37), .Y(n35) );
  OAI21XL U165 ( .A0(n15), .A1(n39), .B0(n40), .Y(n37) );
  NOR2BX1 U166 ( .AN(n167), .B(n12), .Y(n190) );
  NOR2BX1 U167 ( .AN(n166), .B(n191), .Y(n194) );
  OAI21XL U168 ( .A0(n29), .A1(n30), .B0(n31), .Y(n25) );
  INVX1 U169 ( .A(n32), .Y(n29) );
  INVX1 U170 ( .A(n68), .Y(n46) );
  NOR2BX1 U171 ( .AN(n40), .B(n15), .Y(n41) );
  NOR2BX1 U172 ( .AN(n31), .B(n30), .Y(n33) );
  NOR2BX1 U173 ( .AN(n47), .B(n46), .Y(n67) );
  NOR2BX1 U174 ( .AN(n23), .B(n24), .Y(n22) );
  OAI21XL U175 ( .A0(n45), .A1(n46), .B0(n47), .Y(n42) );
  INVX1 U176 ( .A(n48), .Y(n45) );
  OAI2BB1X1 U177 ( .A0N(n69), .A1N(n70), .B0(n71), .Y(n48) );
  INVX1 U178 ( .A(n149), .Y(n70) );
  NOR2X1 U179 ( .A(A[19]), .B(B[19]), .Y(n11) );
  NAND2XL U180 ( .A(A[29]), .B(B[29]), .Y(n55) );
  NAND2XL U181 ( .A(B[26]), .B(A[26]), .Y(n92) );
  OR2X2 U182 ( .A(A[24]), .B(B[24]), .Y(n101) );
  OR2X2 U183 ( .A(A[23]), .B(B[23]), .Y(n118) );
  OR2X2 U184 ( .A(A[22]), .B(B[22]), .Y(n117) );
  NAND2XL U185 ( .A(B[26]), .B(A[26]), .Y(n85) );
  NAND2X1 U186 ( .A(A[24]), .B(B[24]), .Y(n83) );
  OR2X2 U187 ( .A(A[21]), .B(B[21]), .Y(n124) );
  NAND2X1 U188 ( .A(B[16]), .B(A[16]), .Y(n144) );
  NAND2X1 U189 ( .A(B[20]), .B(A[20]), .Y(n112) );
  NAND2X1 U190 ( .A(B[17]), .B(A[17]), .Y(n145) );
  NAND2X1 U191 ( .A(B[21]), .B(A[21]), .Y(n113) );
  OR2X2 U192 ( .A(A[16]), .B(B[16]), .Y(n137) );
  OR2X2 U193 ( .A(A[15]), .B(B[15]), .Y(n182) );
  OR2X2 U194 ( .A(A[14]), .B(B[14]), .Y(n181) );
  OR2X2 U195 ( .A(A[17]), .B(B[17]), .Y(n138) );
  OR2X2 U196 ( .A(A[20]), .B(B[20]), .Y(n128) );
  OR2X2 U197 ( .A(A[18]), .B(B[18]), .Y(n152) );
  NOR2X1 U198 ( .A(A[9]), .B(B[9]), .Y(n13) );
  NAND2X1 U199 ( .A(B[12]), .B(A[12]), .Y(n166) );
  NAND2X1 U200 ( .A(B[10]), .B(A[10]), .Y(n210) );
  OR2X2 U201 ( .A(A[12]), .B(B[12]), .Y(n180) );
  NOR2X1 U202 ( .A(A[5]), .B(B[5]), .Y(n14) );
  NOR2X1 U203 ( .A(A[4]), .B(B[4]), .Y(n15) );
  NAND2X1 U204 ( .A(B[4]), .B(A[4]), .Y(n40) );
  NAND2X1 U205 ( .A(B[8]), .B(A[8]), .Y(n23) );
  NAND2X1 U206 ( .A(B[5]), .B(A[5]), .Y(n36) );
  NAND2X1 U207 ( .A(B[6]), .B(A[6]), .Y(n31) );
  NAND2X1 U208 ( .A(B[2]), .B(A[2]), .Y(n47) );
  OR2X2 U209 ( .A(A[6]), .B(B[6]), .Y(n34) );
  NOR2X1 U210 ( .A(A[3]), .B(B[3]), .Y(n16) );
  OR2X2 U211 ( .A(A[8]), .B(B[8]), .Y(n206) );
  OR2X2 U212 ( .A(A[1]), .B(B[1]), .Y(n69) );
  NAND2X1 U213 ( .A(B[1]), .B(A[1]), .Y(n71) );
  NAND2X1 U214 ( .A(B[0]), .B(A[0]), .Y(n149) );
  NOR2X1 U215 ( .A(A[0]), .B(B[0]), .Y(n17) );
  NAND2XL U216 ( .A(n59), .B(n63), .Y(n72) );
  XOR2X1 U217 ( .A(n97), .B(n98), .Y(SUM[25]) );
  XOR2X1 U218 ( .A(n93), .B(n94), .Y(SUM[26]) );
  NOR2BXL U219 ( .AN(n92), .B(n86), .Y(n94) );
  XOR2X1 U220 ( .A(n89), .B(n90), .Y(SUM[27]) );
  NOR2BXL U221 ( .AN(n81), .B(n2), .Y(n90) );
  XOR2X1 U222 ( .A(n66), .B(n75), .Y(SUM[28]) );
  NOR2BX1 U223 ( .AN(n65), .B(n64), .Y(n75) );
  XOR2X1 U224 ( .A(n122), .B(n123), .Y(SUM[22]) );
  XOR2X1 U225 ( .A(n119), .B(n120), .Y(SUM[23]) );
  XOR2X1 U226 ( .A(n100), .B(n102), .Y(SUM[24]) );
  NOR2BX1 U227 ( .AN(n99), .B(n103), .Y(n102) );
  NOR2BX1 U228 ( .AN(n149), .B(n17), .Y(SUM[0]) );
  XOR2X1 U229 ( .A(n70), .B(n147), .Y(SUM[1]) );
  XOR2X1 U230 ( .A(n48), .B(n67), .Y(SUM[2]) );
  XOR2X1 U231 ( .A(n42), .B(n43), .Y(SUM[3]) );
  XOR2X1 U232 ( .A(n177), .B(n41), .Y(SUM[4]) );
  XOR2X1 U233 ( .A(n37), .B(n38), .Y(SUM[5]) );
  XOR2X1 U234 ( .A(n32), .B(n33), .Y(SUM[6]) );
  XOR2X1 U235 ( .A(n25), .B(n26), .Y(SUM[7]) );
  XOR2X1 U236 ( .A(n21), .B(n22), .Y(SUM[8]) );
  XOR2X1 U237 ( .A(n18), .B(n19), .Y(SUM[9]) );
  XOR2X1 U238 ( .A(n209), .B(n211), .Y(SUM[10]) );
  XOR2X1 U239 ( .A(n207), .B(n208), .Y(SUM[11]) );
  XOR2X1 U240 ( .A(n193), .B(n194), .Y(SUM[12]) );
  XOR2X1 U241 ( .A(n189), .B(n190), .Y(SUM[13]) );
  XOR2X1 U242 ( .A(n186), .B(n187), .Y(SUM[14]) );
  XOR2X1 U243 ( .A(n183), .B(n184), .Y(SUM[15]) );
  XOR2X1 U244 ( .A(n134), .B(n159), .Y(SUM[16]) );
  XOR2X1 U245 ( .A(n156), .B(n157), .Y(SUM[17]) );
  XOR2X1 U246 ( .A(n153), .B(n154), .Y(SUM[18]) );
  XOR2X1 U247 ( .A(n150), .B(n151), .Y(SUM[19]) );
  XOR2X1 U248 ( .A(n127), .B(n129), .Y(SUM[20]) );
  NOR2BX1 U249 ( .AN(n112), .B(n130), .Y(n129) );
  XOR2X1 U250 ( .A(n125), .B(n126), .Y(SUM[21]) );
  NOR2X4 U251 ( .A(A[30]), .B(B[30]), .Y(n54) );
  OR2X4 U252 ( .A(A[29]), .B(B[29]), .Y(n59) );
  CLKINVX3 U253 ( .A(n87), .Y(n86) );
  OR2X4 U254 ( .A(A[26]), .B(B[26]), .Y(n87) );
endmodule


module message_schedule ( clk, reset, data, write_enable, inner_busy, Wt );
  input [31:0] data;
  output [31:0] Wt;
  input clk, reset, write_enable, inner_busy;
  wire   N622, N623, N624, N625, N626, N627, N628, n578, n613, n614, n615, N9,
         N8, N7, N67, N66, N65, N64, N63, N62, N61, N60, N6, N59, N58, N57,
         N56, N55, N54, N53, N52, N51, N50, N5, N49, N48, N47, N46, N45, N44,
         N43, N42, N41, N40, N4, N39, N38, N37, N36, N35, N34, N33, N32, N31,
         N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17,
         N16, N15, N14, N13, N12, N11, N10, n20, n21, n23, n376, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638;
  wire   [31:0] R14;
  wire   [31:0] sigma0;
  wire   [31:0] R1;
  wire   [31:0] sigma1;
  wire   [31:0] R15;
  wire   [31:0] R6;
  wire   [31:0] logic_result;
  wire   [6:0] counter;
  wire   [31:0] R2;
  wire   [31:0] R3;
  wire   [31:0] R4;
  wire   [31:0] R5;
  wire   [31:0] R7;
  wire   [31:0] R8;
  wire   [31:0] R9;
  wire   [31:0] R10;
  wire   [31:0] R11;
  wire   [31:0] R12;
  wire   [31:0] R13;

  DFFHQX4 Wt_reg_15_ ( .D(n622), .CK(clk), .Q(Wt[15]) );
  DFFHQX4 Wt_reg_14_ ( .D(n623), .CK(clk), .Q(Wt[14]) );
  DFFHQX4 Wt_reg_13_ ( .D(n624), .CK(clk), .Q(Wt[13]) );
  DFFHQX4 Wt_reg_12_ ( .D(n625), .CK(clk), .Q(Wt[12]) );
  DFFHQX4 Wt_reg_11_ ( .D(n626), .CK(clk), .Q(Wt[11]) );
  DFFHQX4 Wt_reg_10_ ( .D(n627), .CK(clk), .Q(Wt[10]) );
  DFFHQX4 Wt_reg_9_ ( .D(n628), .CK(clk), .Q(Wt[9]) );
  DFFHQX4 Wt_reg_8_ ( .D(n629), .CK(clk), .Q(Wt[8]) );
  DFFHQX4 Wt_reg_7_ ( .D(n630), .CK(clk), .Q(Wt[7]) );
  DFFHQX4 Wt_reg_6_ ( .D(n631), .CK(clk), .Q(Wt[6]) );
  DFFHQX4 Wt_reg_5_ ( .D(n632), .CK(clk), .Q(Wt[5]) );
  DFFHQX4 Wt_reg_4_ ( .D(n633), .CK(clk), .Q(Wt[4]) );
  DFFHQX4 Wt_reg_3_ ( .D(n634), .CK(clk), .Q(Wt[3]) );
  DFFHQX4 Wt_reg_2_ ( .D(n635), .CK(clk), .Q(Wt[2]) );
  DFFHQX4 Wt_reg_1_ ( .D(n636), .CK(clk), .Q(Wt[1]) );
  DFFTRX4 R6_reg_1_ ( .D(R5[1]), .RN(n498), .CK(clk), .Q(R6[1]) );
  DFFTRX4 R15_reg_1_ ( .D(R14[1]), .RN(n497), .CK(clk), .Q(R15[1]) );
  DFFHQX4 Wt_reg_0_ ( .D(n637), .CK(clk), .Q(Wt[0]) );
  DFFTRX4 R6_reg_0_ ( .D(R5[0]), .RN(n496), .CK(clk), .Q(R6[0]) );
  DFFTRX4 R15_reg_0_ ( .D(R14[0]), .RN(n496), .CK(clk), .Q(R15[0]) );
  message_schedule_DW01_inc_0 add_110 ( .A(counter), .SUM({N628, N627, N626, 
        N625, N624, N623, N622}) );
  message_schedule_DW01_add_2 add_2_root_add_0_root_add_34_3 ( .A(R15), .B(R6), 
        .SUM({N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, 
        N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, 
        N40, N39, N38, N37, N36}) );
  message_schedule_DW01_add_6 add_1_root_add_0_root_add_34_3 ( .A(sigma1), .B(
        sigma0), .SUM({N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4}) );
  message_schedule_DW01_add_8 add_0_root_add_0_root_add_34_3 ( .A({N67, N66, 
        N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, 
        N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, 
        N37, N36}), .B({N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4}), .SUM(logic_result) );
  DFFTRX1 R15_reg_31_ ( .D(R14[31]), .RN(n534), .CK(clk), .Q(R15[31]) );
  DFFTRX1 R15_reg_30_ ( .D(R14[30]), .RN(n533), .CK(clk), .Q(R15[30]) );
  DFFTRX1 counter_reg_6_ ( .D(N628), .RN(n534), .CK(clk), .Q(counter[6]) );
  DFFTRX1 R6_reg_31_ ( .D(R5[31]), .RN(n535), .CK(clk), .Q(R6[31]) );
  DFFTRX1 R6_reg_30_ ( .D(R5[30]), .RN(n534), .CK(clk), .Q(R6[30]) );
  DFFTRX1 counter_reg_1_ ( .D(N623), .RN(n531), .CK(clk), .Q(counter[1]) );
  DFFTRX1 counter_reg_0_ ( .D(N622), .RN(n532), .CK(clk), .Q(counter[0]) );
  DFFTRX1 R15_reg_29_ ( .D(R14[29]), .RN(n532), .CK(clk), .Q(R15[29]) );
  DFFTRX1 R15_reg_28_ ( .D(R14[28]), .RN(n531), .CK(clk), .Q(R15[28]) );
  DFFTRX1 R15_reg_27_ ( .D(R14[27]), .RN(n529), .CK(clk), .Q(R15[27]) );
  DFFTRX1 R15_reg_26_ ( .D(R14[26]), .RN(n528), .CK(clk), .Q(R15[26]) );
  DFFTRX1 R6_reg_29_ ( .D(R5[29]), .RN(n533), .CK(clk), .Q(R6[29]) );
  DFFTRX1 R6_reg_28_ ( .D(R5[28]), .RN(n531), .CK(clk), .Q(R6[28]) );
  DFFTRX1 R6_reg_27_ ( .D(R5[27]), .RN(n530), .CK(clk), .Q(R6[27]) );
  DFFTRX1 R6_reg_26_ ( .D(R5[26]), .RN(n529), .CK(clk), .Q(R6[26]) );
  DFFTRX1 counter_reg_5_ ( .D(N627), .RN(n535), .CK(clk), .Q(counter[5]) );
  DFFTRX1 counter_reg_3_ ( .D(N625), .RN(n535), .CK(clk), .Q(counter[3]) );
  DFFTRX1 counter_reg_4_ ( .D(N626), .RN(n534), .CK(clk), .Q(counter[4]) );
  DFFTRX1 counter_reg_2_ ( .D(N624), .RN(n533), .CK(clk), .Q(counter[2]) );
  DFFTRX1 R15_reg_25_ ( .D(R14[25]), .RN(n527), .CK(clk), .Q(R15[25]) );
  DFFTRX1 R15_reg_24_ ( .D(R14[24]), .RN(n526), .CK(clk), .Q(R15[24]) );
  DFFTRX1 R15_reg_23_ ( .D(R14[23]), .RN(n524), .CK(clk), .Q(R15[23]) );
  DFFTRX1 R15_reg_22_ ( .D(R14[22]), .RN(n523), .CK(clk), .Q(R15[22]) );
  DFFTRX1 R6_reg_25_ ( .D(R5[25]), .RN(n528), .CK(clk), .Q(R6[25]) );
  DFFTRX1 R6_reg_24_ ( .D(R5[24]), .RN(n526), .CK(clk), .Q(R6[24]) );
  DFFTRX1 R6_reg_23_ ( .D(R5[23]), .RN(n525), .CK(clk), .Q(R6[23]) );
  DFFTRX1 R6_reg_22_ ( .D(R5[22]), .RN(n524), .CK(clk), .Q(R6[22]) );
  DFFHQXL Wt_reg_31_ ( .D(n603), .CK(clk), .Q(Wt[31]) );
  DFFTRX1 R15_reg_21_ ( .D(R14[21]), .RN(n522), .CK(clk), .Q(R15[21]) );
  DFFTRX1 R15_reg_20_ ( .D(R14[20]), .RN(n521), .CK(clk), .Q(R15[20]) );
  DFFTRX1 R15_reg_19_ ( .D(R14[19]), .RN(n519), .CK(clk), .Q(R15[19]) );
  DFFTRX1 R15_reg_18_ ( .D(R14[18]), .RN(n518), .CK(clk), .Q(R15[18]) );
  DFFTRX1 R6_reg_21_ ( .D(R5[21]), .RN(n523), .CK(clk), .Q(R6[21]) );
  DFFTRX1 R6_reg_20_ ( .D(R5[20]), .RN(n521), .CK(clk), .Q(R6[20]) );
  DFFTRX1 R6_reg_19_ ( .D(R5[19]), .RN(n520), .CK(clk), .Q(R6[19]) );
  DFFTRX1 R6_reg_18_ ( .D(R5[18]), .RN(n519), .CK(clk), .Q(R6[18]) );
  DFFTRX1 R14_reg_2_ ( .D(R13[2]), .RN(n498), .CK(clk), .Q(R14[2]) );
  DFFTRX1 R1_reg_9_ ( .D(Wt[9]), .RN(n508), .CK(clk), .Q(R1[9]) );
  DFFTRX1 R1_reg_6_ ( .D(Wt[6]), .RN(n504), .CK(clk), .Q(R1[6]) );
  DFFTRX1 R1_reg_8_ ( .D(Wt[8]), .RN(n507), .CK(clk), .Q(R1[8]) );
  DFFTRX1 R1_reg_7_ ( .D(Wt[7]), .RN(n505), .CK(clk), .Q(R1[7]) );
  DFFHQXL Wt_reg_30_ ( .D(n604), .CK(clk), .Q(Wt[30]) );
  DFFTRX1 R15_reg_17_ ( .D(R14[17]), .RN(n517), .CK(clk), .Q(R15[17]) );
  DFFTRX1 R15_reg_16_ ( .D(R14[16]), .RN(n516), .CK(clk), .Q(R15[16]) );
  DFFTRX1 R15_reg_15_ ( .D(R14[15]), .RN(n514), .CK(clk), .Q(R15[15]) );
  DFFTRX1 R15_reg_14_ ( .D(R14[14]), .RN(n513), .CK(clk), .Q(R15[14]) );
  DFFTRX1 R6_reg_17_ ( .D(R5[17]), .RN(n518), .CK(clk), .Q(R6[17]) );
  DFFTRX1 R6_reg_16_ ( .D(R5[16]), .RN(n516), .CK(clk), .Q(R6[16]) );
  DFFTRX1 R6_reg_15_ ( .D(R5[15]), .RN(n515), .CK(clk), .Q(R6[15]) );
  DFFTRX1 R6_reg_14_ ( .D(R5[14]), .RN(n514), .CK(clk), .Q(R6[14]) );
  DFFTRX1 R14_reg_1_ ( .D(R13[1]), .RN(n497), .CK(clk), .Q(R14[1]) );
  DFFTRX1 R14_reg_0_ ( .D(R13[0]), .RN(n496), .CK(clk), .Q(R14[0]) );
  DFFTRX1 R1_reg_5_ ( .D(Wt[5]), .RN(n503), .CK(clk), .Q(R1[5]) );
  DFFTRX1 R1_reg_4_ ( .D(Wt[4]), .RN(n502), .CK(clk), .Q(R1[4]) );
  DFFTRX1 R1_reg_2_ ( .D(Wt[2]), .RN(n499), .CK(clk), .Q(R1[2]) );
  DFFTRX1 R1_reg_29_ ( .D(Wt[29]), .RN(n533), .CK(clk), .Q(R1[29]) );
  DFFTRX1 R1_reg_27_ ( .D(Wt[27]), .RN(n530), .CK(clk), .Q(R1[27]) );
  DFFTRX1 R14_reg_26_ ( .D(R13[26]), .RN(n528), .CK(clk), .Q(R14[26]) );
  DFFTRX1 R1_reg_31_ ( .D(Wt[31]), .RN(n535), .CK(clk), .Q(R1[31]) );
  DFFTRX1 R1_reg_30_ ( .D(Wt[30]), .RN(n534), .CK(clk), .Q(R1[30]) );
  DFFTRX1 R14_reg_15_ ( .D(R13[15]), .RN(n514), .CK(clk), .Q(R14[15]) );
  DFFTRX1 R14_reg_17_ ( .D(R13[17]), .RN(n517), .CK(clk), .Q(R14[17]) );
  DFFTRX1 R14_reg_31_ ( .D(R13[31]), .RN(n534), .CK(clk), .Q(R14[31]) );
  DFFTRX1 R14_reg_30_ ( .D(R13[30]), .RN(n533), .CK(clk), .Q(R14[30]) );
  DFFTRX1 R14_reg_29_ ( .D(R13[29]), .RN(n532), .CK(clk), .Q(R14[29]) );
  DFFTRX1 R1_reg_0_ ( .D(Wt[0]), .RN(n497), .CK(clk), .Q(R1[0]) );
  DFFTRX1 R1_reg_3_ ( .D(Wt[3]), .RN(n500), .CK(clk), .Q(R1[3]) );
  DFFTRX1 R15_reg_13_ ( .D(R14[13]), .RN(n512), .CK(clk), .Q(R15[13]) );
  DFFTRX1 R15_reg_12_ ( .D(R14[12]), .RN(n511), .CK(clk), .Q(R15[12]) );
  DFFTRX1 R15_reg_11_ ( .D(R14[11]), .RN(n509), .CK(clk), .Q(R15[11]) );
  DFFTRX1 R15_reg_10_ ( .D(R14[10]), .RN(n508), .CK(clk), .Q(R15[10]) );
  DFFTRX1 R6_reg_13_ ( .D(R5[13]), .RN(n513), .CK(clk), .Q(R6[13]) );
  DFFTRX1 R6_reg_12_ ( .D(R5[12]), .RN(n511), .CK(clk), .Q(R6[12]) );
  DFFTRX1 R6_reg_11_ ( .D(R5[11]), .RN(n510), .CK(clk), .Q(R6[11]) );
  DFFTRX1 R6_reg_10_ ( .D(R5[10]), .RN(n509), .CK(clk), .Q(R6[10]) );
  DFFTRX1 R14_reg_19_ ( .D(R13[19]), .RN(n519), .CK(clk), .Q(R14[19]) );
  DFFTRX1 R14_reg_18_ ( .D(R13[18]), .RN(n518), .CK(clk), .Q(R14[18]) );
  DFFHQX1 Wt_reg_23_ ( .D(n611), .CK(clk), .Q(Wt[23]) );
  DFFTRX1 R14_reg_3_ ( .D(R13[3]), .RN(n499), .CK(clk), .Q(R14[3]) );
  DFFTRX1 R14_reg_6_ ( .D(R13[6]), .RN(n503), .CK(clk), .Q(R14[6]) );
  DFFTRX1 R14_reg_5_ ( .D(R13[5]), .RN(n502), .CK(clk), .Q(R14[5]) );
  DFFTRX1 R14_reg_4_ ( .D(R13[4]), .RN(n501), .CK(clk), .Q(R14[4]) );
  DFFTRX1 R1_reg_28_ ( .D(Wt[28]), .RN(n532), .CK(clk), .Q(R1[28]) );
  DFFTRX1 R14_reg_27_ ( .D(R13[27]), .RN(n529), .CK(clk), .Q(R14[27]) );
  DFFTRX1 R1_reg_26_ ( .D(Wt[26]), .RN(n529), .CK(clk), .Q(R1[26]) );
  DFFTRX1 R1_reg_25_ ( .D(Wt[25]), .RN(n528), .CK(clk), .Q(R1[25]) );
  DFFTRX1 R14_reg_25_ ( .D(R13[25]), .RN(n527), .CK(clk), .Q(R14[25]) );
  DFFTRX1 R14_reg_24_ ( .D(R13[24]), .RN(n526), .CK(clk), .Q(R14[24]) );
  DFFTRX1 R14_reg_14_ ( .D(R13[14]), .RN(n513), .CK(clk), .Q(R14[14]) );
  DFFTRX1 R14_reg_13_ ( .D(R13[13]), .RN(n512), .CK(clk), .Q(R14[13]) );
  DFFTRX1 R1_reg_16_ ( .D(Wt[16]), .RN(n517), .CK(clk), .Q(R1[16]) );
  DFFTRX1 R1_reg_15_ ( .D(Wt[15]), .RN(n515), .CK(clk), .Q(R1[15]) );
  DFFTRX1 R1_reg_14_ ( .D(Wt[14]), .RN(n514), .CK(clk), .Q(R1[14]) );
  DFFTRX1 R1_reg_13_ ( .D(Wt[13]), .RN(n513), .CK(clk), .Q(R1[13]) );
  DFFTRX1 R1_reg_12_ ( .D(Wt[12]), .RN(n512), .CK(clk), .Q(R1[12]) );
  DFFTRX1 R1_reg_11_ ( .D(Wt[11]), .RN(n510), .CK(clk), .Q(R1[11]) );
  DFFTRX1 R1_reg_10_ ( .D(Wt[10]), .RN(n509), .CK(clk), .Q(R1[10]) );
  DFFTRX1 R14_reg_9_ ( .D(R13[9]), .RN(n507), .CK(clk), .Q(R14[9]) );
  DFFTRX1 R14_reg_7_ ( .D(R13[7]), .RN(n504), .CK(clk), .Q(R14[7]) );
  DFFTRX1 R14_reg_28_ ( .D(R13[28]), .RN(n531), .CK(clk), .Q(R14[28]) );
  DFFTRX1 R1_reg_18_ ( .D(Wt[18]), .RN(n519), .CK(clk), .Q(R1[18]) );
  DFFTRX1 R1_reg_17_ ( .D(Wt[17]), .RN(n518), .CK(clk), .Q(R1[17]) );
  DFFTRX1 R14_reg_16_ ( .D(R13[16]), .RN(n516), .CK(clk), .Q(R14[16]) );
  DFFTRX1 R15_reg_9_ ( .D(R14[9]), .RN(n507), .CK(clk), .Q(R15[9]) );
  DFFTRX1 R15_reg_8_ ( .D(R14[8]), .RN(n506), .CK(clk), .Q(R15[8]) );
  DFFTRX1 R15_reg_7_ ( .D(R14[7]), .RN(n504), .CK(clk), .Q(R15[7]) );
  DFFTRX1 R15_reg_6_ ( .D(R14[6]), .RN(n503), .CK(clk), .Q(R15[6]) );
  DFFTRX1 R6_reg_9_ ( .D(R5[9]), .RN(n508), .CK(clk), .Q(R6[9]) );
  DFFTRX1 R6_reg_8_ ( .D(R5[8]), .RN(n506), .CK(clk), .Q(R6[8]) );
  DFFTRX1 R6_reg_7_ ( .D(R5[7]), .RN(n505), .CK(clk), .Q(R6[7]) );
  DFFTRX1 R6_reg_6_ ( .D(R5[6]), .RN(n504), .CK(clk), .Q(R6[6]) );
  DFFHQX1 Wt_reg_20_ ( .D(n617), .CK(clk), .Q(Wt[20]) );
  DFFTRX1 R15_reg_5_ ( .D(R14[5]), .RN(n502), .CK(clk), .Q(R15[5]) );
  DFFTRX1 R15_reg_4_ ( .D(R14[4]), .RN(n501), .CK(clk), .Q(R15[4]) );
  DFFTRX1 R15_reg_3_ ( .D(R14[3]), .RN(n499), .CK(clk), .Q(R15[3]) );
  DFFTRX1 R6_reg_5_ ( .D(R5[5]), .RN(n503), .CK(clk), .Q(R6[5]) );
  DFFTRX1 R6_reg_4_ ( .D(R5[4]), .RN(n501), .CK(clk), .Q(R6[4]) );
  DFFTRX1 R6_reg_3_ ( .D(R5[3]), .RN(n500), .CK(clk), .Q(R6[3]) );
  DFFHQX1 Wt_reg_19_ ( .D(n618), .CK(clk), .Q(Wt[19]) );
  DFFHQX1 Wt_reg_18_ ( .D(n619), .CK(clk), .Q(Wt[18]) );
  DFFHQX1 Wt_reg_16_ ( .D(n621), .CK(clk), .Q(Wt[16]) );
  DFFTRX1 R2_reg_31_ ( .D(R1[31]), .RN(n535), .CK(clk), .Q(R2[31]) );
  DFFTRX1 R3_reg_31_ ( .D(R2[31]), .RN(n535), .CK(clk), .Q(R3[31]) );
  DFFTRX1 R4_reg_31_ ( .D(R3[31]), .RN(n535), .CK(clk), .Q(R4[31]) );
  DFFTRX1 R5_reg_31_ ( .D(R4[31]), .RN(n535), .CK(clk), .Q(R5[31]) );
  DFFTRX1 R7_reg_31_ ( .D(R6[31]), .RN(n535), .CK(clk), .Q(R7[31]) );
  DFFTRX1 R8_reg_31_ ( .D(R7[31]), .RN(n535), .CK(clk), .Q(R8[31]) );
  DFFTRX1 R9_reg_31_ ( .D(R8[31]), .RN(n535), .CK(clk), .Q(R9[31]) );
  DFFTRX1 R10_reg_31_ ( .D(R9[31]), .RN(n535), .CK(clk), .Q(R10[31]) );
  DFFTRX1 R11_reg_31_ ( .D(R10[31]), .RN(n535), .CK(clk), .Q(R11[31]) );
  DFFTRX1 R12_reg_31_ ( .D(R11[31]), .RN(n535), .CK(clk), .Q(R12[31]) );
  DFFTRX1 R13_reg_31_ ( .D(R12[31]), .RN(n534), .CK(clk), .Q(R13[31]) );
  DFFTRX1 R2_reg_30_ ( .D(R1[30]), .RN(n534), .CK(clk), .Q(R2[30]) );
  DFFTRX1 R3_reg_30_ ( .D(R2[30]), .RN(n534), .CK(clk), .Q(R3[30]) );
  DFFTRX1 R4_reg_30_ ( .D(R3[30]), .RN(n534), .CK(clk), .Q(R4[30]) );
  DFFTRX1 R5_reg_30_ ( .D(R4[30]), .RN(n534), .CK(clk), .Q(R5[30]) );
  DFFTRX1 R7_reg_30_ ( .D(R6[30]), .RN(n534), .CK(clk), .Q(R7[30]) );
  DFFTRX1 R8_reg_30_ ( .D(R7[30]), .RN(n534), .CK(clk), .Q(R8[30]) );
  DFFTRX1 R9_reg_30_ ( .D(R8[30]), .RN(n534), .CK(clk), .Q(R9[30]) );
  DFFTRX1 R10_reg_30_ ( .D(R9[30]), .RN(n533), .CK(clk), .Q(R10[30]) );
  DFFTRX1 R11_reg_30_ ( .D(R10[30]), .RN(n533), .CK(clk), .Q(R11[30]) );
  DFFTRX1 R12_reg_30_ ( .D(R11[30]), .RN(n533), .CK(clk), .Q(R12[30]) );
  DFFTRX1 R13_reg_30_ ( .D(R12[30]), .RN(n533), .CK(clk), .Q(R13[30]) );
  DFFTRX1 R2_reg_29_ ( .D(R1[29]), .RN(n533), .CK(clk), .Q(R2[29]) );
  DFFTRX1 R3_reg_29_ ( .D(R2[29]), .RN(n533), .CK(clk), .Q(R3[29]) );
  DFFTRX1 R4_reg_29_ ( .D(R3[29]), .RN(n533), .CK(clk), .Q(R4[29]) );
  DFFTRX1 R5_reg_29_ ( .D(R4[29]), .RN(n533), .CK(clk), .Q(R5[29]) );
  DFFTRX1 R7_reg_29_ ( .D(R6[29]), .RN(n532), .CK(clk), .Q(R7[29]) );
  DFFTRX1 R8_reg_29_ ( .D(R7[29]), .RN(n532), .CK(clk), .Q(R8[29]) );
  DFFTRX1 R9_reg_29_ ( .D(R8[29]), .RN(n532), .CK(clk), .Q(R9[29]) );
  DFFTRX1 R10_reg_29_ ( .D(R9[29]), .RN(n532), .CK(clk), .Q(R10[29]) );
  DFFTRX1 R11_reg_29_ ( .D(R10[29]), .RN(n532), .CK(clk), .Q(R11[29]) );
  DFFTRX1 R12_reg_29_ ( .D(R11[29]), .RN(n532), .CK(clk), .Q(R12[29]) );
  DFFTRX1 R13_reg_29_ ( .D(R12[29]), .RN(n532), .CK(clk), .Q(R13[29]) );
  DFFTRX1 R2_reg_28_ ( .D(R1[28]), .RN(n532), .CK(clk), .Q(R2[28]) );
  DFFTRX1 R3_reg_28_ ( .D(R2[28]), .RN(n532), .CK(clk), .Q(R3[28]) );
  DFFTRX1 R4_reg_28_ ( .D(R3[28]), .RN(n531), .CK(clk), .Q(R4[28]) );
  DFFTRX1 R5_reg_28_ ( .D(R4[28]), .RN(n531), .CK(clk), .Q(R5[28]) );
  DFFTRX1 R7_reg_28_ ( .D(R6[28]), .RN(n531), .CK(clk), .Q(R7[28]) );
  DFFTRX1 R8_reg_28_ ( .D(R7[28]), .RN(n531), .CK(clk), .Q(R8[28]) );
  DFFTRX1 R9_reg_28_ ( .D(R8[28]), .RN(n531), .CK(clk), .Q(R9[28]) );
  DFFTRX1 R10_reg_28_ ( .D(R9[28]), .RN(n531), .CK(clk), .Q(R10[28]) );
  DFFTRX1 R11_reg_28_ ( .D(R10[28]), .RN(n531), .CK(clk), .Q(R11[28]) );
  DFFTRX1 R12_reg_28_ ( .D(R11[28]), .RN(n531), .CK(clk), .Q(R12[28]) );
  DFFTRX1 R13_reg_28_ ( .D(R12[28]), .RN(n531), .CK(clk), .Q(R13[28]) );
  DFFTRX1 R4_reg_0_ ( .D(R3[0]), .RN(n496), .CK(clk), .Q(R4[0]) );
  DFFTRX1 R5_reg_0_ ( .D(R4[0]), .RN(n496), .CK(clk), .Q(R5[0]) );
  DFFTRX1 R8_reg_0_ ( .D(R7[0]), .RN(n496), .CK(clk), .Q(R8[0]) );
  DFFTRX1 R9_reg_0_ ( .D(R8[0]), .RN(n496), .CK(clk), .Q(R9[0]) );
  DFFTRX1 R10_reg_0_ ( .D(R9[0]), .RN(n496), .CK(clk), .Q(R10[0]) );
  DFFTRX1 R11_reg_0_ ( .D(R10[0]), .RN(n496), .CK(clk), .Q(R11[0]) );
  DFFTRX1 R12_reg_0_ ( .D(R11[0]), .RN(n496), .CK(clk), .Q(R12[0]) );
  DFFTRX1 R13_reg_0_ ( .D(R12[0]), .RN(n496), .CK(clk), .Q(R13[0]) );
  DFFTRX1 R2_reg_27_ ( .D(R1[27]), .RN(n530), .CK(clk), .Q(R2[27]) );
  DFFTRX1 R3_reg_27_ ( .D(R2[27]), .RN(n530), .CK(clk), .Q(R3[27]) );
  DFFTRX1 R4_reg_27_ ( .D(R3[27]), .RN(n530), .CK(clk), .Q(R4[27]) );
  DFFTRX1 R5_reg_27_ ( .D(R4[27]), .RN(n530), .CK(clk), .Q(R5[27]) );
  DFFTRX1 R7_reg_27_ ( .D(R6[27]), .RN(n530), .CK(clk), .Q(R7[27]) );
  DFFTRX1 R8_reg_27_ ( .D(R7[27]), .RN(n530), .CK(clk), .Q(R8[27]) );
  DFFTRX1 R9_reg_27_ ( .D(R8[27]), .RN(n530), .CK(clk), .Q(R9[27]) );
  DFFTRX1 R10_reg_27_ ( .D(R9[27]), .RN(n530), .CK(clk), .Q(R10[27]) );
  DFFTRX1 R11_reg_27_ ( .D(R10[27]), .RN(n530), .CK(clk), .Q(R11[27]) );
  DFFTRX1 R12_reg_27_ ( .D(R11[27]), .RN(n530), .CK(clk), .Q(R12[27]) );
  DFFTRX1 R13_reg_27_ ( .D(R12[27]), .RN(n529), .CK(clk), .Q(R13[27]) );
  DFFTRX1 R2_reg_26_ ( .D(R1[26]), .RN(n529), .CK(clk), .Q(R2[26]) );
  DFFTRX1 R3_reg_26_ ( .D(R2[26]), .RN(n529), .CK(clk), .Q(R3[26]) );
  DFFTRX1 R4_reg_26_ ( .D(R3[26]), .RN(n529), .CK(clk), .Q(R4[26]) );
  DFFTRX1 R5_reg_26_ ( .D(R4[26]), .RN(n529), .CK(clk), .Q(R5[26]) );
  DFFTRX1 R7_reg_26_ ( .D(R6[26]), .RN(n529), .CK(clk), .Q(R7[26]) );
  DFFTRX1 R8_reg_26_ ( .D(R7[26]), .RN(n529), .CK(clk), .Q(R8[26]) );
  DFFTRX1 R9_reg_26_ ( .D(R8[26]), .RN(n529), .CK(clk), .Q(R9[26]) );
  DFFTRX1 R10_reg_26_ ( .D(R9[26]), .RN(n528), .CK(clk), .Q(R10[26]) );
  DFFTRX1 R11_reg_26_ ( .D(R10[26]), .RN(n528), .CK(clk), .Q(R11[26]) );
  DFFTRX1 R12_reg_26_ ( .D(R11[26]), .RN(n528), .CK(clk), .Q(R12[26]) );
  DFFTRX1 R13_reg_26_ ( .D(R12[26]), .RN(n528), .CK(clk), .Q(R13[26]) );
  DFFTRX1 R2_reg_25_ ( .D(R1[25]), .RN(n528), .CK(clk), .Q(R2[25]) );
  DFFTRX1 R3_reg_25_ ( .D(R2[25]), .RN(n528), .CK(clk), .Q(R3[25]) );
  DFFTRX1 R4_reg_25_ ( .D(R3[25]), .RN(n528), .CK(clk), .Q(R4[25]) );
  DFFTRX1 R5_reg_25_ ( .D(R4[25]), .RN(n528), .CK(clk), .Q(R5[25]) );
  DFFTRX1 R7_reg_25_ ( .D(R6[25]), .RN(n527), .CK(clk), .Q(R7[25]) );
  DFFTRX1 R8_reg_25_ ( .D(R7[25]), .RN(n527), .CK(clk), .Q(R8[25]) );
  DFFTRX1 R9_reg_25_ ( .D(R8[25]), .RN(n527), .CK(clk), .Q(R9[25]) );
  DFFTRX1 R10_reg_25_ ( .D(R9[25]), .RN(n527), .CK(clk), .Q(R10[25]) );
  DFFTRX1 R11_reg_25_ ( .D(R10[25]), .RN(n527), .CK(clk), .Q(R11[25]) );
  DFFTRX1 R12_reg_25_ ( .D(R11[25]), .RN(n527), .CK(clk), .Q(R12[25]) );
  DFFTRX1 R13_reg_25_ ( .D(R12[25]), .RN(n527), .CK(clk), .Q(R13[25]) );
  DFFTRX1 R2_reg_24_ ( .D(R1[24]), .RN(n527), .CK(clk), .Q(R2[24]) );
  DFFTRX1 R3_reg_24_ ( .D(R2[24]), .RN(n527), .CK(clk), .Q(R3[24]) );
  DFFTRX1 R4_reg_24_ ( .D(R3[24]), .RN(n526), .CK(clk), .Q(R4[24]) );
  DFFTRX1 R5_reg_24_ ( .D(R4[24]), .RN(n526), .CK(clk), .Q(R5[24]) );
  DFFTRX1 R7_reg_24_ ( .D(R6[24]), .RN(n526), .CK(clk), .Q(R7[24]) );
  DFFTRX1 R8_reg_24_ ( .D(R7[24]), .RN(n526), .CK(clk), .Q(R8[24]) );
  DFFTRX1 R9_reg_24_ ( .D(R8[24]), .RN(n526), .CK(clk), .Q(R9[24]) );
  DFFTRX1 R10_reg_24_ ( .D(R9[24]), .RN(n526), .CK(clk), .Q(R10[24]) );
  DFFTRX1 R11_reg_24_ ( .D(R10[24]), .RN(n526), .CK(clk), .Q(R11[24]) );
  DFFTRX1 R12_reg_24_ ( .D(R11[24]), .RN(n526), .CK(clk), .Q(R12[24]) );
  DFFTRX1 R13_reg_24_ ( .D(R12[24]), .RN(n526), .CK(clk), .Q(R13[24]) );
  DFFTRX1 R2_reg_23_ ( .D(R1[23]), .RN(n525), .CK(clk), .Q(R2[23]) );
  DFFTRX1 R3_reg_23_ ( .D(R2[23]), .RN(n525), .CK(clk), .Q(R3[23]) );
  DFFTRX1 R4_reg_23_ ( .D(R3[23]), .RN(n525), .CK(clk), .Q(R4[23]) );
  DFFTRX1 R5_reg_23_ ( .D(R4[23]), .RN(n525), .CK(clk), .Q(R5[23]) );
  DFFTRX1 R7_reg_23_ ( .D(R6[23]), .RN(n525), .CK(clk), .Q(R7[23]) );
  DFFTRX1 R8_reg_23_ ( .D(R7[23]), .RN(n525), .CK(clk), .Q(R8[23]) );
  DFFTRX1 R9_reg_23_ ( .D(R8[23]), .RN(n525), .CK(clk), .Q(R9[23]) );
  DFFTRX1 R10_reg_23_ ( .D(R9[23]), .RN(n525), .CK(clk), .Q(R10[23]) );
  DFFTRX1 R11_reg_23_ ( .D(R10[23]), .RN(n525), .CK(clk), .Q(R11[23]) );
  DFFTRX1 R12_reg_23_ ( .D(R11[23]), .RN(n525), .CK(clk), .Q(R12[23]) );
  DFFTRX1 R13_reg_23_ ( .D(R12[23]), .RN(n524), .CK(clk), .Q(R13[23]) );
  DFFTRX1 R2_reg_22_ ( .D(R1[22]), .RN(n524), .CK(clk), .Q(R2[22]) );
  DFFTRX1 R3_reg_22_ ( .D(R2[22]), .RN(n524), .CK(clk), .Q(R3[22]) );
  DFFTRX1 R4_reg_22_ ( .D(R3[22]), .RN(n524), .CK(clk), .Q(R4[22]) );
  DFFTRX1 R5_reg_22_ ( .D(R4[22]), .RN(n524), .CK(clk), .Q(R5[22]) );
  DFFTRX1 R7_reg_22_ ( .D(R6[22]), .RN(n524), .CK(clk), .Q(R7[22]) );
  DFFTRX1 R8_reg_22_ ( .D(R7[22]), .RN(n524), .CK(clk), .Q(R8[22]) );
  DFFTRX1 R9_reg_22_ ( .D(R8[22]), .RN(n524), .CK(clk), .Q(R9[22]) );
  DFFTRX1 R10_reg_22_ ( .D(R9[22]), .RN(n523), .CK(clk), .Q(R10[22]) );
  DFFTRX1 R11_reg_22_ ( .D(R10[22]), .RN(n523), .CK(clk), .Q(R11[22]) );
  DFFTRX1 R12_reg_22_ ( .D(R11[22]), .RN(n523), .CK(clk), .Q(R12[22]) );
  DFFTRX1 R13_reg_22_ ( .D(R12[22]), .RN(n523), .CK(clk), .Q(R13[22]) );
  DFFTRX1 R2_reg_21_ ( .D(R1[21]), .RN(n523), .CK(clk), .Q(R2[21]) );
  DFFTRX1 R3_reg_21_ ( .D(R2[21]), .RN(n523), .CK(clk), .Q(R3[21]) );
  DFFTRX1 R4_reg_21_ ( .D(R3[21]), .RN(n523), .CK(clk), .Q(R4[21]) );
  DFFTRX1 R5_reg_21_ ( .D(R4[21]), .RN(n523), .CK(clk), .Q(R5[21]) );
  DFFTRX1 R7_reg_21_ ( .D(R6[21]), .RN(n522), .CK(clk), .Q(R7[21]) );
  DFFTRX1 R8_reg_21_ ( .D(R7[21]), .RN(n522), .CK(clk), .Q(R8[21]) );
  DFFTRX1 R9_reg_21_ ( .D(R8[21]), .RN(n522), .CK(clk), .Q(R9[21]) );
  DFFTRX1 R10_reg_21_ ( .D(R9[21]), .RN(n522), .CK(clk), .Q(R10[21]) );
  DFFTRX1 R11_reg_21_ ( .D(R10[21]), .RN(n522), .CK(clk), .Q(R11[21]) );
  DFFTRX1 R12_reg_21_ ( .D(R11[21]), .RN(n522), .CK(clk), .Q(R12[21]) );
  DFFTRX1 R13_reg_21_ ( .D(R12[21]), .RN(n522), .CK(clk), .Q(R13[21]) );
  DFFTRX1 R2_reg_20_ ( .D(R1[20]), .RN(n522), .CK(clk), .Q(R2[20]) );
  DFFTRX1 R3_reg_20_ ( .D(R2[20]), .RN(n522), .CK(clk), .Q(R3[20]) );
  DFFTRX1 R4_reg_20_ ( .D(R3[20]), .RN(n521), .CK(clk), .Q(R4[20]) );
  DFFTRX1 R5_reg_20_ ( .D(R4[20]), .RN(n521), .CK(clk), .Q(R5[20]) );
  DFFTRX1 R7_reg_20_ ( .D(R6[20]), .RN(n521), .CK(clk), .Q(R7[20]) );
  DFFTRX1 R8_reg_20_ ( .D(R7[20]), .RN(n521), .CK(clk), .Q(R8[20]) );
  DFFTRX1 R9_reg_20_ ( .D(R8[20]), .RN(n521), .CK(clk), .Q(R9[20]) );
  DFFTRX1 R10_reg_20_ ( .D(R9[20]), .RN(n521), .CK(clk), .Q(R10[20]) );
  DFFTRX1 R11_reg_20_ ( .D(R10[20]), .RN(n521), .CK(clk), .Q(R11[20]) );
  DFFTRX1 R12_reg_20_ ( .D(R11[20]), .RN(n521), .CK(clk), .Q(R12[20]) );
  DFFTRX1 R13_reg_20_ ( .D(R12[20]), .RN(n521), .CK(clk), .Q(R13[20]) );
  DFFTRX1 R2_reg_19_ ( .D(R1[19]), .RN(n520), .CK(clk), .Q(R2[19]) );
  DFFTRX1 R3_reg_19_ ( .D(R2[19]), .RN(n520), .CK(clk), .Q(R3[19]) );
  DFFTRX1 R4_reg_19_ ( .D(R3[19]), .RN(n520), .CK(clk), .Q(R4[19]) );
  DFFTRX1 R5_reg_19_ ( .D(R4[19]), .RN(n520), .CK(clk), .Q(R5[19]) );
  DFFTRX1 R7_reg_19_ ( .D(R6[19]), .RN(n520), .CK(clk), .Q(R7[19]) );
  DFFTRX1 R8_reg_19_ ( .D(R7[19]), .RN(n520), .CK(clk), .Q(R8[19]) );
  DFFTRX1 R9_reg_19_ ( .D(R8[19]), .RN(n520), .CK(clk), .Q(R9[19]) );
  DFFTRX1 R10_reg_19_ ( .D(R9[19]), .RN(n520), .CK(clk), .Q(R10[19]) );
  DFFTRX1 R11_reg_19_ ( .D(R10[19]), .RN(n520), .CK(clk), .Q(R11[19]) );
  DFFTRX1 R12_reg_19_ ( .D(R11[19]), .RN(n520), .CK(clk), .Q(R12[19]) );
  DFFTRX1 R13_reg_19_ ( .D(R12[19]), .RN(n519), .CK(clk), .Q(R13[19]) );
  DFFTRX1 R2_reg_18_ ( .D(R1[18]), .RN(n519), .CK(clk), .Q(R2[18]) );
  DFFTRX1 R3_reg_18_ ( .D(R2[18]), .RN(n519), .CK(clk), .Q(R3[18]) );
  DFFTRX1 R4_reg_18_ ( .D(R3[18]), .RN(n519), .CK(clk), .Q(R4[18]) );
  DFFTRX1 R5_reg_18_ ( .D(R4[18]), .RN(n519), .CK(clk), .Q(R5[18]) );
  DFFTRX1 R7_reg_18_ ( .D(R6[18]), .RN(n519), .CK(clk), .Q(R7[18]) );
  DFFTRX1 R8_reg_18_ ( .D(R7[18]), .RN(n519), .CK(clk), .Q(R8[18]) );
  DFFTRX1 R9_reg_18_ ( .D(R8[18]), .RN(n519), .CK(clk), .Q(R9[18]) );
  DFFTRX1 R10_reg_18_ ( .D(R9[18]), .RN(n518), .CK(clk), .Q(R10[18]) );
  DFFTRX1 R11_reg_18_ ( .D(R10[18]), .RN(n518), .CK(clk), .Q(R11[18]) );
  DFFTRX1 R12_reg_18_ ( .D(R11[18]), .RN(n518), .CK(clk), .Q(R12[18]) );
  DFFTRX1 R13_reg_18_ ( .D(R12[18]), .RN(n518), .CK(clk), .Q(R13[18]) );
  DFFTRX1 R2_reg_17_ ( .D(R1[17]), .RN(n518), .CK(clk), .Q(R2[17]) );
  DFFTRX1 R3_reg_17_ ( .D(R2[17]), .RN(n518), .CK(clk), .Q(R3[17]) );
  DFFTRX1 R4_reg_17_ ( .D(R3[17]), .RN(n518), .CK(clk), .Q(R4[17]) );
  DFFTRX1 R5_reg_17_ ( .D(R4[17]), .RN(n518), .CK(clk), .Q(R5[17]) );
  DFFTRX1 R7_reg_17_ ( .D(R6[17]), .RN(n517), .CK(clk), .Q(R7[17]) );
  DFFTRX1 R8_reg_17_ ( .D(R7[17]), .RN(n517), .CK(clk), .Q(R8[17]) );
  DFFTRX1 R9_reg_17_ ( .D(R8[17]), .RN(n517), .CK(clk), .Q(R9[17]) );
  DFFTRX1 R10_reg_17_ ( .D(R9[17]), .RN(n517), .CK(clk), .Q(R10[17]) );
  DFFTRX1 R11_reg_17_ ( .D(R10[17]), .RN(n517), .CK(clk), .Q(R11[17]) );
  DFFTRX1 R12_reg_17_ ( .D(R11[17]), .RN(n517), .CK(clk), .Q(R12[17]) );
  DFFTRX1 R13_reg_17_ ( .D(R12[17]), .RN(n517), .CK(clk), .Q(R13[17]) );
  DFFTRX1 R2_reg_16_ ( .D(R1[16]), .RN(n517), .CK(clk), .Q(R2[16]) );
  DFFTRX1 R3_reg_16_ ( .D(R2[16]), .RN(n517), .CK(clk), .Q(R3[16]) );
  DFFTRX1 R4_reg_16_ ( .D(R3[16]), .RN(n516), .CK(clk), .Q(R4[16]) );
  DFFTRX1 R5_reg_16_ ( .D(R4[16]), .RN(n516), .CK(clk), .Q(R5[16]) );
  DFFTRX1 R7_reg_16_ ( .D(R6[16]), .RN(n516), .CK(clk), .Q(R7[16]) );
  DFFTRX1 R8_reg_16_ ( .D(R7[16]), .RN(n516), .CK(clk), .Q(R8[16]) );
  DFFTRX1 R9_reg_16_ ( .D(R8[16]), .RN(n516), .CK(clk), .Q(R9[16]) );
  DFFTRX1 R10_reg_16_ ( .D(R9[16]), .RN(n516), .CK(clk), .Q(R10[16]) );
  DFFTRX1 R11_reg_16_ ( .D(R10[16]), .RN(n516), .CK(clk), .Q(R11[16]) );
  DFFTRX1 R12_reg_16_ ( .D(R11[16]), .RN(n516), .CK(clk), .Q(R12[16]) );
  DFFTRX1 R13_reg_16_ ( .D(R12[16]), .RN(n516), .CK(clk), .Q(R13[16]) );
  DFFTRX1 R2_reg_15_ ( .D(R1[15]), .RN(n515), .CK(clk), .Q(R2[15]) );
  DFFTRX1 R3_reg_15_ ( .D(R2[15]), .RN(n515), .CK(clk), .Q(R3[15]) );
  DFFTRX1 R4_reg_15_ ( .D(R3[15]), .RN(n515), .CK(clk), .Q(R4[15]) );
  DFFTRX1 R5_reg_15_ ( .D(R4[15]), .RN(n515), .CK(clk), .Q(R5[15]) );
  DFFTRX1 R7_reg_15_ ( .D(R6[15]), .RN(n515), .CK(clk), .Q(R7[15]) );
  DFFTRX1 R8_reg_15_ ( .D(R7[15]), .RN(n515), .CK(clk), .Q(R8[15]) );
  DFFTRX1 R9_reg_15_ ( .D(R8[15]), .RN(n515), .CK(clk), .Q(R9[15]) );
  DFFTRX1 R10_reg_15_ ( .D(R9[15]), .RN(n515), .CK(clk), .Q(R10[15]) );
  DFFTRX1 R11_reg_15_ ( .D(R10[15]), .RN(n515), .CK(clk), .Q(R11[15]) );
  DFFTRX1 R12_reg_15_ ( .D(R11[15]), .RN(n515), .CK(clk), .Q(R12[15]) );
  DFFTRX1 R13_reg_15_ ( .D(R12[15]), .RN(n514), .CK(clk), .Q(R13[15]) );
  DFFTRX1 R2_reg_14_ ( .D(R1[14]), .RN(n514), .CK(clk), .Q(R2[14]) );
  DFFTRX1 R3_reg_14_ ( .D(R2[14]), .RN(n514), .CK(clk), .Q(R3[14]) );
  DFFTRX1 R4_reg_14_ ( .D(R3[14]), .RN(n514), .CK(clk), .Q(R4[14]) );
  DFFTRX1 R5_reg_14_ ( .D(R4[14]), .RN(n514), .CK(clk), .Q(R5[14]) );
  DFFTRX1 R7_reg_14_ ( .D(R6[14]), .RN(n514), .CK(clk), .Q(R7[14]) );
  DFFTRX1 R8_reg_14_ ( .D(R7[14]), .RN(n514), .CK(clk), .Q(R8[14]) );
  DFFTRX1 R9_reg_14_ ( .D(R8[14]), .RN(n514), .CK(clk), .Q(R9[14]) );
  DFFTRX1 R10_reg_14_ ( .D(R9[14]), .RN(n513), .CK(clk), .Q(R10[14]) );
  DFFTRX1 R11_reg_14_ ( .D(R10[14]), .RN(n513), .CK(clk), .Q(R11[14]) );
  DFFTRX1 R12_reg_14_ ( .D(R11[14]), .RN(n513), .CK(clk), .Q(R12[14]) );
  DFFTRX1 R13_reg_14_ ( .D(R12[14]), .RN(n513), .CK(clk), .Q(R13[14]) );
  DFFTRX1 R2_reg_13_ ( .D(R1[13]), .RN(n513), .CK(clk), .Q(R2[13]) );
  DFFTRX1 R3_reg_13_ ( .D(R2[13]), .RN(n513), .CK(clk), .Q(R3[13]) );
  DFFTRX1 R4_reg_13_ ( .D(R3[13]), .RN(n513), .CK(clk), .Q(R4[13]) );
  DFFTRX1 R5_reg_13_ ( .D(R4[13]), .RN(n513), .CK(clk), .Q(R5[13]) );
  DFFTRX1 R7_reg_13_ ( .D(R6[13]), .RN(n512), .CK(clk), .Q(R7[13]) );
  DFFTRX1 R8_reg_13_ ( .D(R7[13]), .RN(n512), .CK(clk), .Q(R8[13]) );
  DFFTRX1 R9_reg_13_ ( .D(R8[13]), .RN(n512), .CK(clk), .Q(R9[13]) );
  DFFTRX1 R10_reg_13_ ( .D(R9[13]), .RN(n512), .CK(clk), .Q(R10[13]) );
  DFFTRX1 R11_reg_13_ ( .D(R10[13]), .RN(n512), .CK(clk), .Q(R11[13]) );
  DFFTRX1 R12_reg_13_ ( .D(R11[13]), .RN(n512), .CK(clk), .Q(R12[13]) );
  DFFTRX1 R13_reg_13_ ( .D(R12[13]), .RN(n512), .CK(clk), .Q(R13[13]) );
  DFFTRX1 R2_reg_12_ ( .D(R1[12]), .RN(n512), .CK(clk), .Q(R2[12]) );
  DFFTRX1 R3_reg_12_ ( .D(R2[12]), .RN(n512), .CK(clk), .Q(R3[12]) );
  DFFTRX1 R4_reg_12_ ( .D(R3[12]), .RN(n511), .CK(clk), .Q(R4[12]) );
  DFFTRX1 R5_reg_12_ ( .D(R4[12]), .RN(n511), .CK(clk), .Q(R5[12]) );
  DFFTRX1 R7_reg_12_ ( .D(R6[12]), .RN(n511), .CK(clk), .Q(R7[12]) );
  DFFTRX1 R8_reg_12_ ( .D(R7[12]), .RN(n511), .CK(clk), .Q(R8[12]) );
  DFFTRX1 R9_reg_12_ ( .D(R8[12]), .RN(n511), .CK(clk), .Q(R9[12]) );
  DFFTRX1 R10_reg_12_ ( .D(R9[12]), .RN(n511), .CK(clk), .Q(R10[12]) );
  DFFTRX1 R11_reg_12_ ( .D(R10[12]), .RN(n511), .CK(clk), .Q(R11[12]) );
  DFFTRX1 R12_reg_12_ ( .D(R11[12]), .RN(n511), .CK(clk), .Q(R12[12]) );
  DFFTRX1 R13_reg_12_ ( .D(R12[12]), .RN(n511), .CK(clk), .Q(R13[12]) );
  DFFTRX1 R2_reg_11_ ( .D(R1[11]), .RN(n510), .CK(clk), .Q(R2[11]) );
  DFFTRX1 R3_reg_11_ ( .D(R2[11]), .RN(n510), .CK(clk), .Q(R3[11]) );
  DFFTRX1 R4_reg_11_ ( .D(R3[11]), .RN(n510), .CK(clk), .Q(R4[11]) );
  DFFTRX1 R5_reg_11_ ( .D(R4[11]), .RN(n510), .CK(clk), .Q(R5[11]) );
  DFFTRX1 R7_reg_11_ ( .D(R6[11]), .RN(n510), .CK(clk), .Q(R7[11]) );
  DFFTRX1 R8_reg_11_ ( .D(R7[11]), .RN(n510), .CK(clk), .Q(R8[11]) );
  DFFTRX1 R9_reg_11_ ( .D(R8[11]), .RN(n510), .CK(clk), .Q(R9[11]) );
  DFFTRX1 R10_reg_11_ ( .D(R9[11]), .RN(n510), .CK(clk), .Q(R10[11]) );
  DFFTRX1 R11_reg_11_ ( .D(R10[11]), .RN(n510), .CK(clk), .Q(R11[11]) );
  DFFTRX1 R12_reg_11_ ( .D(R11[11]), .RN(n510), .CK(clk), .Q(R12[11]) );
  DFFTRX1 R13_reg_11_ ( .D(R12[11]), .RN(n509), .CK(clk), .Q(R13[11]) );
  DFFTRX1 R2_reg_10_ ( .D(R1[10]), .RN(n509), .CK(clk), .Q(R2[10]) );
  DFFTRX1 R3_reg_10_ ( .D(R2[10]), .RN(n509), .CK(clk), .Q(R3[10]) );
  DFFTRX1 R4_reg_10_ ( .D(R3[10]), .RN(n509), .CK(clk), .Q(R4[10]) );
  DFFTRX1 R5_reg_10_ ( .D(R4[10]), .RN(n509), .CK(clk), .Q(R5[10]) );
  DFFTRX1 R7_reg_10_ ( .D(R6[10]), .RN(n509), .CK(clk), .Q(R7[10]) );
  DFFTRX1 R8_reg_10_ ( .D(R7[10]), .RN(n509), .CK(clk), .Q(R8[10]) );
  DFFTRX1 R9_reg_10_ ( .D(R8[10]), .RN(n509), .CK(clk), .Q(R9[10]) );
  DFFTRX1 R10_reg_10_ ( .D(R9[10]), .RN(n508), .CK(clk), .Q(R10[10]) );
  DFFTRX1 R11_reg_10_ ( .D(R10[10]), .RN(n508), .CK(clk), .Q(R11[10]) );
  DFFTRX1 R12_reg_10_ ( .D(R11[10]), .RN(n508), .CK(clk), .Q(R12[10]) );
  DFFTRX1 R13_reg_10_ ( .D(R12[10]), .RN(n508), .CK(clk), .Q(R13[10]) );
  DFFTRX1 R2_reg_9_ ( .D(R1[9]), .RN(n508), .CK(clk), .Q(R2[9]) );
  DFFTRX1 R3_reg_9_ ( .D(R2[9]), .RN(n508), .CK(clk), .Q(R3[9]) );
  DFFTRX1 R4_reg_9_ ( .D(R3[9]), .RN(n508), .CK(clk), .Q(R4[9]) );
  DFFTRX1 R5_reg_9_ ( .D(R4[9]), .RN(n508), .CK(clk), .Q(R5[9]) );
  DFFTRX1 R7_reg_9_ ( .D(R6[9]), .RN(n507), .CK(clk), .Q(R7[9]) );
  DFFTRX1 R8_reg_9_ ( .D(R7[9]), .RN(n507), .CK(clk), .Q(R8[9]) );
  DFFTRX1 R9_reg_9_ ( .D(R8[9]), .RN(n507), .CK(clk), .Q(R9[9]) );
  DFFTRX1 R10_reg_9_ ( .D(R9[9]), .RN(n507), .CK(clk), .Q(R10[9]) );
  DFFTRX1 R11_reg_9_ ( .D(R10[9]), .RN(n507), .CK(clk), .Q(R11[9]) );
  DFFTRX1 R12_reg_9_ ( .D(R11[9]), .RN(n507), .CK(clk), .Q(R12[9]) );
  DFFTRX1 R13_reg_9_ ( .D(R12[9]), .RN(n507), .CK(clk), .Q(R13[9]) );
  DFFTRX1 R2_reg_8_ ( .D(R1[8]), .RN(n507), .CK(clk), .Q(R2[8]) );
  DFFTRX1 R3_reg_8_ ( .D(R2[8]), .RN(n507), .CK(clk), .Q(R3[8]) );
  DFFTRX1 R4_reg_8_ ( .D(R3[8]), .RN(n506), .CK(clk), .Q(R4[8]) );
  DFFTRX1 R5_reg_8_ ( .D(R4[8]), .RN(n506), .CK(clk), .Q(R5[8]) );
  DFFTRX1 R7_reg_8_ ( .D(R6[8]), .RN(n506), .CK(clk), .Q(R7[8]) );
  DFFTRX1 R8_reg_8_ ( .D(R7[8]), .RN(n506), .CK(clk), .Q(R8[8]) );
  DFFTRX1 R9_reg_8_ ( .D(R8[8]), .RN(n506), .CK(clk), .Q(R9[8]) );
  DFFTRX1 R10_reg_8_ ( .D(R9[8]), .RN(n506), .CK(clk), .Q(R10[8]) );
  DFFTRX1 R11_reg_8_ ( .D(R10[8]), .RN(n506), .CK(clk), .Q(R11[8]) );
  DFFTRX1 R12_reg_8_ ( .D(R11[8]), .RN(n506), .CK(clk), .Q(R12[8]) );
  DFFTRX1 R13_reg_8_ ( .D(R12[8]), .RN(n506), .CK(clk), .Q(R13[8]) );
  DFFTRX1 R2_reg_7_ ( .D(R1[7]), .RN(n505), .CK(clk), .Q(R2[7]) );
  DFFTRX1 R3_reg_7_ ( .D(R2[7]), .RN(n505), .CK(clk), .Q(R3[7]) );
  DFFTRX1 R4_reg_7_ ( .D(R3[7]), .RN(n505), .CK(clk), .Q(R4[7]) );
  DFFTRX1 R5_reg_7_ ( .D(R4[7]), .RN(n505), .CK(clk), .Q(R5[7]) );
  DFFTRX1 R7_reg_7_ ( .D(R6[7]), .RN(n505), .CK(clk), .Q(R7[7]) );
  DFFTRX1 R8_reg_7_ ( .D(R7[7]), .RN(n505), .CK(clk), .Q(R8[7]) );
  DFFTRX1 R9_reg_7_ ( .D(R8[7]), .RN(n505), .CK(clk), .Q(R9[7]) );
  DFFTRX1 R10_reg_7_ ( .D(R9[7]), .RN(n505), .CK(clk), .Q(R10[7]) );
  DFFTRX1 R11_reg_7_ ( .D(R10[7]), .RN(n505), .CK(clk), .Q(R11[7]) );
  DFFTRX1 R12_reg_7_ ( .D(R11[7]), .RN(n505), .CK(clk), .Q(R12[7]) );
  DFFTRX1 R13_reg_7_ ( .D(R12[7]), .RN(n504), .CK(clk), .Q(R13[7]) );
  DFFTRX1 R2_reg_6_ ( .D(R1[6]), .RN(n504), .CK(clk), .Q(R2[6]) );
  DFFTRX1 R3_reg_6_ ( .D(R2[6]), .RN(n504), .CK(clk), .Q(R3[6]) );
  DFFTRX1 R4_reg_6_ ( .D(R3[6]), .RN(n504), .CK(clk), .Q(R4[6]) );
  DFFTRX1 R5_reg_6_ ( .D(R4[6]), .RN(n504), .CK(clk), .Q(R5[6]) );
  DFFTRX1 R7_reg_6_ ( .D(R6[6]), .RN(n504), .CK(clk), .Q(R7[6]) );
  DFFTRX1 R8_reg_6_ ( .D(R7[6]), .RN(n504), .CK(clk), .Q(R8[6]) );
  DFFTRX1 R9_reg_6_ ( .D(R8[6]), .RN(n504), .CK(clk), .Q(R9[6]) );
  DFFTRX1 R10_reg_6_ ( .D(R9[6]), .RN(n503), .CK(clk), .Q(R10[6]) );
  DFFTRX1 R11_reg_6_ ( .D(R10[6]), .RN(n503), .CK(clk), .Q(R11[6]) );
  DFFTRX1 R12_reg_6_ ( .D(R11[6]), .RN(n503), .CK(clk), .Q(R12[6]) );
  DFFTRX1 R13_reg_6_ ( .D(R12[6]), .RN(n503), .CK(clk), .Q(R13[6]) );
  DFFTRX1 R2_reg_5_ ( .D(R1[5]), .RN(n503), .CK(clk), .Q(R2[5]) );
  DFFTRX1 R3_reg_5_ ( .D(R2[5]), .RN(n503), .CK(clk), .Q(R3[5]) );
  DFFTRX1 R4_reg_5_ ( .D(R3[5]), .RN(n503), .CK(clk), .Q(R4[5]) );
  DFFTRX1 R5_reg_5_ ( .D(R4[5]), .RN(n503), .CK(clk), .Q(R5[5]) );
  DFFTRX1 R7_reg_5_ ( .D(R6[5]), .RN(n502), .CK(clk), .Q(R7[5]) );
  DFFTRX1 R8_reg_5_ ( .D(R7[5]), .RN(n502), .CK(clk), .Q(R8[5]) );
  DFFTRX1 R9_reg_5_ ( .D(R8[5]), .RN(n502), .CK(clk), .Q(R9[5]) );
  DFFTRX1 R10_reg_5_ ( .D(R9[5]), .RN(n502), .CK(clk), .Q(R10[5]) );
  DFFTRX1 R11_reg_5_ ( .D(R10[5]), .RN(n502), .CK(clk), .Q(R11[5]) );
  DFFTRX1 R12_reg_5_ ( .D(R11[5]), .RN(n502), .CK(clk), .Q(R12[5]) );
  DFFTRX1 R13_reg_5_ ( .D(R12[5]), .RN(n502), .CK(clk), .Q(R13[5]) );
  DFFTRX1 R2_reg_4_ ( .D(R1[4]), .RN(n502), .CK(clk), .Q(R2[4]) );
  DFFTRX1 R3_reg_4_ ( .D(R2[4]), .RN(n502), .CK(clk), .Q(R3[4]) );
  DFFTRX1 R4_reg_4_ ( .D(R3[4]), .RN(n501), .CK(clk), .Q(R4[4]) );
  DFFTRX1 R5_reg_4_ ( .D(R4[4]), .RN(n501), .CK(clk), .Q(R5[4]) );
  DFFTRX1 R7_reg_4_ ( .D(R6[4]), .RN(n501), .CK(clk), .Q(R7[4]) );
  DFFTRX1 R8_reg_4_ ( .D(R7[4]), .RN(n501), .CK(clk), .Q(R8[4]) );
  DFFTRX1 R9_reg_4_ ( .D(R8[4]), .RN(n501), .CK(clk), .Q(R9[4]) );
  DFFTRX1 R10_reg_4_ ( .D(R9[4]), .RN(n501), .CK(clk), .Q(R10[4]) );
  DFFTRX1 R11_reg_4_ ( .D(R10[4]), .RN(n501), .CK(clk), .Q(R11[4]) );
  DFFTRX1 R12_reg_4_ ( .D(R11[4]), .RN(n501), .CK(clk), .Q(R12[4]) );
  DFFTRX1 R13_reg_4_ ( .D(R12[4]), .RN(n501), .CK(clk), .Q(R13[4]) );
  DFFTRX1 R2_reg_3_ ( .D(R1[3]), .RN(n500), .CK(clk), .Q(R2[3]) );
  DFFTRX1 R3_reg_3_ ( .D(R2[3]), .RN(n500), .CK(clk), .Q(R3[3]) );
  DFFTRX1 R4_reg_3_ ( .D(R3[3]), .RN(n500), .CK(clk), .Q(R4[3]) );
  DFFTRX1 R5_reg_3_ ( .D(R4[3]), .RN(n500), .CK(clk), .Q(R5[3]) );
  DFFTRX1 R7_reg_3_ ( .D(R6[3]), .RN(n500), .CK(clk), .Q(R7[3]) );
  DFFTRX1 R8_reg_3_ ( .D(R7[3]), .RN(n500), .CK(clk), .Q(R8[3]) );
  DFFTRX1 R9_reg_3_ ( .D(R8[3]), .RN(n500), .CK(clk), .Q(R9[3]) );
  DFFTRX1 R10_reg_3_ ( .D(R9[3]), .RN(n500), .CK(clk), .Q(R10[3]) );
  DFFTRX1 R11_reg_3_ ( .D(R10[3]), .RN(n500), .CK(clk), .Q(R11[3]) );
  DFFTRX1 R12_reg_3_ ( .D(R11[3]), .RN(n500), .CK(clk), .Q(R12[3]) );
  DFFTRX1 R13_reg_3_ ( .D(R12[3]), .RN(n499), .CK(clk), .Q(R13[3]) );
  DFFTRX1 R2_reg_2_ ( .D(R1[2]), .RN(n499), .CK(clk), .Q(R2[2]) );
  DFFTRX1 R3_reg_2_ ( .D(R2[2]), .RN(n499), .CK(clk), .Q(R3[2]) );
  DFFTRX1 R4_reg_2_ ( .D(R3[2]), .RN(n499), .CK(clk), .Q(R4[2]) );
  DFFTRX1 R5_reg_2_ ( .D(R4[2]), .RN(n499), .CK(clk), .Q(R5[2]) );
  DFFTRX1 R7_reg_2_ ( .D(R6[2]), .RN(n499), .CK(clk), .Q(R7[2]) );
  DFFTRX1 R8_reg_2_ ( .D(R7[2]), .RN(n499), .CK(clk), .Q(R8[2]) );
  DFFTRX1 R9_reg_2_ ( .D(R8[2]), .RN(n499), .CK(clk), .Q(R9[2]) );
  DFFTRX1 R10_reg_2_ ( .D(R9[2]), .RN(n498), .CK(clk), .Q(R10[2]) );
  DFFTRX1 R11_reg_2_ ( .D(R10[2]), .RN(n498), .CK(clk), .Q(R11[2]) );
  DFFTRX1 R12_reg_2_ ( .D(R11[2]), .RN(n498), .CK(clk), .Q(R12[2]) );
  DFFTRX1 R13_reg_2_ ( .D(R12[2]), .RN(n498), .CK(clk), .Q(R13[2]) );
  DFFTRX1 R2_reg_1_ ( .D(R1[1]), .RN(n498), .CK(clk), .Q(R2[1]) );
  DFFTRX1 R3_reg_1_ ( .D(R2[1]), .RN(n498), .CK(clk), .Q(R3[1]) );
  DFFTRX1 R4_reg_1_ ( .D(R3[1]), .RN(n498), .CK(clk), .Q(R4[1]) );
  DFFTRX1 R5_reg_1_ ( .D(R4[1]), .RN(n498), .CK(clk), .Q(R5[1]) );
  DFFTRX1 R7_reg_1_ ( .D(R6[1]), .RN(n497), .CK(clk), .Q(R7[1]) );
  DFFTRX1 R8_reg_1_ ( .D(R7[1]), .RN(n497), .CK(clk), .Q(R8[1]) );
  DFFTRX1 R9_reg_1_ ( .D(R8[1]), .RN(n497), .CK(clk), .Q(R9[1]) );
  DFFTRX1 R10_reg_1_ ( .D(R9[1]), .RN(n497), .CK(clk), .Q(R10[1]) );
  DFFTRX1 R11_reg_1_ ( .D(R10[1]), .RN(n497), .CK(clk), .Q(R11[1]) );
  DFFTRX1 R12_reg_1_ ( .D(R11[1]), .RN(n497), .CK(clk), .Q(R12[1]) );
  DFFTRX1 R13_reg_1_ ( .D(R12[1]), .RN(n497), .CK(clk), .Q(R13[1]) );
  DFFTRX1 R2_reg_0_ ( .D(R1[0]), .RN(n497), .CK(clk), .Q(R2[0]) );
  DFFTRX1 R3_reg_0_ ( .D(R2[0]), .RN(n497), .CK(clk), .Q(R3[0]) );
  DFFHQXL Wt_reg_25_ ( .D(n609), .CK(clk), .Q(Wt[25]) );
  DFFHQX1 Wt_reg_24_ ( .D(n610), .CK(clk), .Q(Wt[24]) );
  DFFHQXL Wt_reg_27_ ( .D(n607), .CK(clk), .Q(Wt[27]) );
  DFFHQXL Wt_reg_28_ ( .D(n606), .CK(clk), .Q(Wt[28]) );
  DFFHQXL Wt_reg_26_ ( .D(n608), .CK(clk), .Q(Wt[26]) );
  DFFTRX2 R14_reg_22_ ( .D(R13[22]), .RN(n523), .CK(clk), .Q(R14[22]) );
  DFFHQX2 Wt_reg_17_ ( .D(n620), .CK(clk), .Q(Wt[17]) );
  DFFHQXL Wt_reg_29_ ( .D(n605), .CK(clk), .Q(Wt[29]) );
  DFFTRX1 R6_reg_2_ ( .D(R5[2]), .RN(n499), .CK(clk), .Q(R6[2]) );
  DFFTRX1 R15_reg_2_ ( .D(R14[2]), .RN(n498), .CK(clk), .Q(R15[2]) );
  DFFTRX2 R1_reg_21_ ( .D(Wt[21]), .RN(n523), .CK(clk), .Q(R1[21]) );
  DFFHQX1 Wt_reg_21_ ( .D(n616), .CK(clk), .Q(Wt[21]) );
  DFFTRX1 R1_reg_20_ ( .D(Wt[20]), .RN(n522), .CK(clk), .Q(R1[20]) );
  DFFTRX1 R14_reg_11_ ( .D(R13[11]), .RN(n509), .CK(clk), .Q(R14[11]) );
  DFFHQX1 Wt_reg_22_ ( .D(n612), .CK(clk), .Q(Wt[22]) );
  DFFTRX1 R1_reg_23_ ( .D(Wt[23]), .RN(n525), .CK(clk), .Q(R1[23]) );
  DFFTRX1 R1_reg_19_ ( .D(Wt[19]), .RN(n520), .CK(clk), .Q(R1[19]) );
  DFFTRX1 R14_reg_10_ ( .D(R13[10]), .RN(n508), .CK(clk), .Q(R14[10]) );
  DFFTRX1 R1_reg_1_ ( .D(Wt[1]), .RN(n498), .CK(clk), .Q(R1[1]) );
  DFFTRX1 R7_reg_0_ ( .D(R6[0]), .RN(n496), .CK(clk), .Q(R7[0]) );
  DFFTRX2 R14_reg_23_ ( .D(R13[23]), .RN(n524), .CK(clk), .Q(R14[23]) );
  DFFTRX2 R1_reg_22_ ( .D(Wt[22]), .RN(n524), .CK(clk), .Q(R1[22]) );
  DFFTRX2 R14_reg_12_ ( .D(R13[12]), .RN(n511), .CK(clk), .Q(R14[12]) );
  DFFTRX2 R1_reg_24_ ( .D(Wt[24]), .RN(n527), .CK(clk), .Q(R1[24]) );
  DFFTRX2 R14_reg_21_ ( .D(R13[21]), .RN(n522), .CK(clk), .Q(R14[21]) );
  DFFTRX2 R14_reg_8_ ( .D(R13[8]), .RN(n506), .CK(clk), .Q(R14[8]) );
  DFFTRX2 R14_reg_20_ ( .D(R13[20]), .RN(n521), .CK(clk), .Q(R14[20]) );
  XOR3X4 U3 ( .A(R1[22]), .B(R1[24]), .C(R1[15]), .Y(sigma1[5]) );
  XOR3X4 U4 ( .A(R14[23]), .B(R14[12]), .C(R14[8]), .Y(sigma0[5]) );
  XOR3X4 U5 ( .A(R1[20]), .B(R1[22]), .C(R1[13]), .Y(sigma1[3]) );
  XOR3X2 U6 ( .A(R1[19]), .B(R1[21]), .C(R1[12]), .Y(sigma1[2]) );
  XOR3X2 U7 ( .A(R14[22]), .B(R14[11]), .C(R14[7]), .Y(sigma0[4]) );
  XOR3X2 U8 ( .A(R1[21]), .B(R1[23]), .C(R1[14]), .Y(sigma1[4]) );
  OAI2BB1X2 U9 ( .A0N(n491), .A1N(logic_result[29]), .B0(n599), .Y(n605) );
  CLKINVX3 U10 ( .A(n376), .Y(n589) );
  OAI2BB1X4 U11 ( .A0N(logic_result[27]), .A1N(n491), .B0(n597), .Y(n607) );
  XOR2X1 U12 ( .A(R1[13]), .B(R1[15]), .Y(sigma1[28]) );
  OAI2BB1X4 U13 ( .A0N(logic_result[31]), .A1N(n491), .B0(n602), .Y(n603) );
  OAI2BB1X4 U14 ( .A0N(n491), .A1N(logic_result[30]), .B0(n600), .Y(n604) );
  NAND2XL U15 ( .A(inner_busy), .B(n613), .Y(n578) );
  XOR2XL U16 ( .A(R1[16]), .B(R1[18]), .Y(sigma1[31]) );
  NAND2XL U17 ( .A(write_enable), .B(n548), .Y(n20) );
  NAND2XL U18 ( .A(write_enable), .B(n548), .Y(n21) );
  NAND2XL U19 ( .A(write_enable), .B(n548), .Y(n23) );
  XOR2XL U20 ( .A(R1[10]), .B(R1[12]), .Y(sigma1[25]) );
  XOR2XL U21 ( .A(R1[8]), .B(R1[10]), .Y(sigma1[23]) );
  XOR2XL U22 ( .A(R1[9]), .B(R1[11]), .Y(sigma1[24]) );
  XOR2XL U23 ( .A(R1[11]), .B(R1[13]), .Y(sigma1[26]) );
  INVX1 U24 ( .A(n536), .Y(n499) );
  INVX1 U25 ( .A(n546), .Y(n501) );
  INVX1 U26 ( .A(n546), .Y(n502) );
  INVX1 U27 ( .A(n545), .Y(n503) );
  INVX1 U28 ( .A(n545), .Y(n504) );
  INVX1 U29 ( .A(n544), .Y(n505) );
  INVX1 U30 ( .A(n544), .Y(n506) );
  INVX1 U31 ( .A(n543), .Y(n507) );
  INVX1 U32 ( .A(n543), .Y(n508) );
  INVX1 U33 ( .A(n542), .Y(n509) );
  INVX1 U34 ( .A(n542), .Y(n510) );
  INVX1 U35 ( .A(n541), .Y(n511) );
  INVX1 U36 ( .A(n541), .Y(n512) );
  INVX1 U37 ( .A(n540), .Y(n513) );
  INVX1 U38 ( .A(n540), .Y(n514) );
  INVX1 U39 ( .A(n540), .Y(n515) );
  INVX1 U40 ( .A(n540), .Y(n516) );
  INVX1 U41 ( .A(n537), .Y(n517) );
  INVX1 U42 ( .A(n536), .Y(n518) );
  INVX1 U43 ( .A(n539), .Y(n519) );
  INVX1 U44 ( .A(n539), .Y(n520) );
  INVX1 U45 ( .A(n539), .Y(n521) );
  INVX1 U46 ( .A(n539), .Y(n522) );
  INVX1 U47 ( .A(n537), .Y(n523) );
  INVX1 U48 ( .A(n536), .Y(n524) );
  INVX1 U49 ( .A(n538), .Y(n525) );
  INVX1 U50 ( .A(n538), .Y(n526) );
  INVX1 U51 ( .A(n536), .Y(n527) );
  INVX1 U52 ( .A(n538), .Y(n528) );
  INVX1 U53 ( .A(n537), .Y(n529) );
  INVX1 U54 ( .A(n536), .Y(n530) );
  INVX1 U55 ( .A(n537), .Y(n497) );
  INVX1 U56 ( .A(n536), .Y(n498) );
  INVX1 U57 ( .A(n537), .Y(n500) );
  INVX1 U58 ( .A(n547), .Y(n496) );
  INVX1 U59 ( .A(n494), .Y(n547) );
  INVX1 U60 ( .A(n537), .Y(n531) );
  INVX1 U61 ( .A(n537), .Y(n532) );
  INVX1 U62 ( .A(n537), .Y(n533) );
  INVX1 U63 ( .A(n536), .Y(n534) );
  INVX1 U64 ( .A(n536), .Y(n535) );
  INVX1 U65 ( .A(n494), .Y(n546) );
  INVX1 U66 ( .A(n494), .Y(n545) );
  INVX1 U67 ( .A(n494), .Y(n544) );
  INVX1 U68 ( .A(n493), .Y(n543) );
  INVX1 U69 ( .A(n493), .Y(n542) );
  INVX1 U70 ( .A(n493), .Y(n541) );
  INVX1 U71 ( .A(n493), .Y(n540) );
  INVX1 U72 ( .A(n492), .Y(n539) );
  INVX1 U73 ( .A(n492), .Y(n538) );
  INVX1 U74 ( .A(n495), .Y(n494) );
  INVX1 U75 ( .A(n495), .Y(n493) );
  INVX1 U76 ( .A(n495), .Y(n492) );
  INVX1 U77 ( .A(n638), .Y(n537) );
  INVX1 U78 ( .A(n638), .Y(n536) );
  INVX1 U79 ( .A(n638), .Y(n495) );
  INVX1 U80 ( .A(n578), .Y(n548) );
  INVX1 U81 ( .A(n578), .Y(n638) );
  INVX1 U82 ( .A(n20), .Y(n601) );
  BUFX3 U83 ( .A(n376), .Y(n491) );
  NAND2X1 U84 ( .A(data[30]), .B(n601), .Y(n600) );
  NAND2X1 U85 ( .A(data[31]), .B(n601), .Y(n602) );
  NAND2X1 U86 ( .A(data[29]), .B(n601), .Y(n599) );
  OAI2BB1X1 U87 ( .A0N(logic_result[25]), .A1N(n491), .B0(n595), .Y(n609) );
  NAND2X1 U88 ( .A(data[25]), .B(n601), .Y(n595) );
  OAI2BB1X1 U89 ( .A0N(logic_result[26]), .A1N(n491), .B0(n596), .Y(n608) );
  NAND2X1 U90 ( .A(data[26]), .B(n601), .Y(n596) );
  NAND2X1 U91 ( .A(data[27]), .B(n601), .Y(n597) );
  OAI2BB1X1 U92 ( .A0N(logic_result[28]), .A1N(n491), .B0(n598), .Y(n606) );
  NAND2X1 U93 ( .A(data[28]), .B(n601), .Y(n598) );
  OAI2BB1X1 U94 ( .A0N(logic_result[22]), .A1N(n491), .B0(n592), .Y(n612) );
  NAND2X1 U95 ( .A(data[22]), .B(n601), .Y(n592) );
  OAI2BB1X1 U96 ( .A0N(logic_result[23]), .A1N(n491), .B0(n593), .Y(n611) );
  NAND2X1 U97 ( .A(data[23]), .B(n601), .Y(n593) );
  OAI2BB1X1 U98 ( .A0N(logic_result[24]), .A1N(n491), .B0(n594), .Y(n610) );
  NAND2X1 U99 ( .A(data[24]), .B(n601), .Y(n594) );
  XOR3X2 U100 ( .A(R14[18]), .B(R14[7]), .C(R14[3]), .Y(sigma0[0]) );
  XOR3X2 U101 ( .A(R1[19]), .B(R1[17]), .C(R1[10]), .Y(sigma1[0]) );
  AOI31X1 U102 ( .A0(n614), .A1(counter[6]), .A2(n615), .B0(reset), .Y(n613)
         );
  NOR2X1 U103 ( .A(counter[1]), .B(counter[0]), .Y(n614) );
  NOR4X1 U104 ( .A(counter[5]), .B(counter[4]), .C(counter[3]), .D(counter[2]), 
        .Y(n615) );
  OAI22XL U105 ( .A0(n23), .A1(n550), .B0(n589), .B1(n549), .Y(n637) );
  INVX1 U106 ( .A(logic_result[0]), .Y(n549) );
  INVX1 U107 ( .A(data[0]), .Y(n550) );
  OAI22XL U108 ( .A0(n20), .A1(n552), .B0(n589), .B1(n551), .Y(n636) );
  INVX1 U109 ( .A(logic_result[1]), .Y(n551) );
  INVX1 U110 ( .A(data[1]), .Y(n552) );
  OAI22XL U111 ( .A0(n21), .A1(n554), .B0(n589), .B1(n553), .Y(n635) );
  INVX1 U112 ( .A(logic_result[2]), .Y(n553) );
  INVX1 U113 ( .A(data[2]), .Y(n554) );
  OAI22XL U114 ( .A0(n21), .A1(n556), .B0(n589), .B1(n555), .Y(n634) );
  INVX1 U115 ( .A(logic_result[3]), .Y(n555) );
  INVX1 U116 ( .A(data[3]), .Y(n556) );
  OAI22XL U117 ( .A0(n23), .A1(n558), .B0(n589), .B1(n557), .Y(n633) );
  INVX1 U118 ( .A(logic_result[4]), .Y(n557) );
  INVX1 U119 ( .A(data[4]), .Y(n558) );
  OAI22XL U120 ( .A0(n20), .A1(n560), .B0(n589), .B1(n559), .Y(n632) );
  INVX1 U121 ( .A(logic_result[5]), .Y(n559) );
  INVX1 U122 ( .A(data[5]), .Y(n560) );
  OAI22XL U123 ( .A0(n20), .A1(n562), .B0(n589), .B1(n561), .Y(n631) );
  INVX1 U124 ( .A(logic_result[6]), .Y(n561) );
  INVX1 U125 ( .A(data[6]), .Y(n562) );
  OAI22XL U126 ( .A0(n21), .A1(n564), .B0(n589), .B1(n563), .Y(n630) );
  INVX1 U127 ( .A(logic_result[7]), .Y(n563) );
  INVX1 U128 ( .A(data[7]), .Y(n564) );
  OAI22XL U129 ( .A0(n23), .A1(n566), .B0(n589), .B1(n565), .Y(n629) );
  INVX1 U130 ( .A(logic_result[8]), .Y(n565) );
  INVX1 U131 ( .A(data[8]), .Y(n566) );
  OAI22XL U132 ( .A0(n23), .A1(n568), .B0(n589), .B1(n567), .Y(n628) );
  INVX1 U133 ( .A(logic_result[9]), .Y(n567) );
  INVX1 U134 ( .A(data[9]), .Y(n568) );
  OAI22XL U135 ( .A0(n20), .A1(n570), .B0(n589), .B1(n569), .Y(n627) );
  INVX1 U136 ( .A(logic_result[10]), .Y(n569) );
  INVX1 U137 ( .A(data[10]), .Y(n570) );
  OAI22XL U138 ( .A0(n21), .A1(n572), .B0(n589), .B1(n571), .Y(n626) );
  INVX1 U139 ( .A(logic_result[11]), .Y(n571) );
  INVX1 U140 ( .A(data[11]), .Y(n572) );
  OAI22XL U141 ( .A0(n21), .A1(n574), .B0(n589), .B1(n573), .Y(n625) );
  INVX1 U142 ( .A(logic_result[12]), .Y(n573) );
  INVX1 U143 ( .A(data[12]), .Y(n574) );
  OAI22XL U144 ( .A0(n23), .A1(n576), .B0(n589), .B1(n575), .Y(n624) );
  INVX1 U145 ( .A(logic_result[13]), .Y(n575) );
  INVX1 U146 ( .A(data[13]), .Y(n576) );
  OAI22XL U147 ( .A0(n20), .A1(n579), .B0(n589), .B1(n577), .Y(n623) );
  INVX1 U148 ( .A(logic_result[14]), .Y(n577) );
  INVX1 U149 ( .A(data[14]), .Y(n579) );
  OAI22XL U150 ( .A0(n20), .A1(n581), .B0(n589), .B1(n580), .Y(n622) );
  INVX1 U151 ( .A(logic_result[15]), .Y(n580) );
  INVX1 U152 ( .A(data[15]), .Y(n581) );
  OAI22XL U153 ( .A0(n21), .A1(n583), .B0(n589), .B1(n582), .Y(n621) );
  INVX1 U154 ( .A(logic_result[16]), .Y(n582) );
  INVX1 U155 ( .A(data[16]), .Y(n583) );
  OAI22XL U156 ( .A0(n23), .A1(n585), .B0(n589), .B1(n584), .Y(n620) );
  INVX1 U157 ( .A(logic_result[17]), .Y(n584) );
  INVX1 U158 ( .A(data[17]), .Y(n585) );
  OAI22XL U159 ( .A0(n23), .A1(n587), .B0(n589), .B1(n586), .Y(n619) );
  INVX1 U160 ( .A(data[18]), .Y(n587) );
  INVX1 U161 ( .A(logic_result[18]), .Y(n586) );
  NOR2BX1 U162 ( .AN(n548), .B(write_enable), .Y(n376) );
  XOR3X2 U163 ( .A(R14[28]), .B(R14[17]), .C(R14[13]), .Y(sigma0[10]) );
  XOR3X2 U164 ( .A(R14[27]), .B(R14[16]), .C(R14[12]), .Y(sigma0[9]) );
  XOR3X2 U165 ( .A(R14[21]), .B(R14[10]), .C(R14[6]), .Y(sigma0[3]) );
  XOR3X2 U166 ( .A(R14[20]), .B(R14[9]), .C(R14[5]), .Y(sigma0[2]) );
  XOR3X2 U167 ( .A(R14[19]), .B(R14[8]), .C(R14[4]), .Y(sigma0[1]) );
  XOR3X2 U168 ( .A(R14[25]), .B(R14[14]), .C(R14[10]), .Y(sigma0[7]) );
  XOR3X2 U169 ( .A(R14[24]), .B(R14[13]), .C(R14[9]), .Y(sigma0[6]) );
  XOR3X2 U170 ( .A(R1[20]), .B(R1[18]), .C(R1[11]), .Y(sigma1[1]) );
  XOR3X2 U171 ( .A(R1[24]), .B(R1[26]), .C(R1[17]), .Y(sigma1[7]) );
  XOR3X2 U172 ( .A(R1[26]), .B(R1[28]), .C(R1[19]), .Y(sigma1[9]) );
  XOR3X2 U173 ( .A(R1[23]), .B(R1[25]), .C(R1[16]), .Y(sigma1[6]) );
  OAI2BB2X1 U174 ( .B0(n589), .B1(n588), .A0N(data[19]), .A1N(n601), .Y(n618)
         );
  INVX1 U175 ( .A(logic_result[19]), .Y(n588) );
  OAI2BB1X1 U176 ( .A0N(logic_result[20]), .A1N(n491), .B0(n590), .Y(n617) );
  NAND2X1 U177 ( .A(data[20]), .B(n601), .Y(n590) );
  OAI2BB1X1 U178 ( .A0N(logic_result[21]), .A1N(n491), .B0(n591), .Y(n616) );
  NAND2X1 U179 ( .A(data[21]), .B(n601), .Y(n591) );
  XOR3X2 U180 ( .A(R14[18]), .B(R14[29]), .C(R14[14]), .Y(sigma0[11]) );
  XOR3X2 U181 ( .A(R14[19]), .B(R14[30]), .C(R14[15]), .Y(sigma0[12]) );
  XOR3X2 U182 ( .A(R14[20]), .B(R14[31]), .C(R14[16]), .Y(sigma0[13]) );
  XOR3X2 U183 ( .A(R14[21]), .B(R14[17]), .C(R14[0]), .Y(sigma0[14]) );
  XOR3X2 U184 ( .A(R14[26]), .B(R14[15]), .C(R14[11]), .Y(sigma0[8]) );
  XOR3X2 U185 ( .A(R1[26]), .B(R1[3]), .C(R1[1]), .Y(sigma1[16]) );
  XOR3X2 U186 ( .A(R14[18]), .B(R14[22]), .C(R14[1]), .Y(sigma0[15]) );
  XOR3X2 U187 ( .A(R14[20]), .B(R14[24]), .C(R14[3]), .Y(sigma0[17]) );
  XOR3X2 U188 ( .A(R14[22]), .B(R14[26]), .C(R14[5]), .Y(sigma0[19]) );
  XOR3X2 U189 ( .A(R14[19]), .B(R14[23]), .C(R14[2]), .Y(sigma0[16]) );
  XOR3X2 U190 ( .A(R14[21]), .B(R14[25]), .C(R14[4]), .Y(sigma0[18]) );
  XOR3X2 U191 ( .A(R1[28]), .B(R1[30]), .C(R1[21]), .Y(sigma1[11]) );
  XOR3X2 U192 ( .A(R1[24]), .B(R1[31]), .C(R1[1]), .Y(sigma1[14]) );
  XOR3X2 U193 ( .A(R1[29]), .B(R1[31]), .C(R1[22]), .Y(sigma1[12]) );
  XOR3X2 U194 ( .A(R1[23]), .B(R1[30]), .C(R1[0]), .Y(sigma1[13]) );
  XOR3X2 U195 ( .A(R1[25]), .B(R1[27]), .C(R1[18]), .Y(sigma1[8]) );
  XOR3X2 U196 ( .A(R1[27]), .B(R1[29]), .C(R1[20]), .Y(sigma1[10]) );
  XOR3X2 U197 ( .A(R1[25]), .B(R1[2]), .C(R1[0]), .Y(sigma1[15]) );
  XOR3X2 U198 ( .A(R1[27]), .B(R1[4]), .C(R1[2]), .Y(sigma1[17]) );
  XOR3X2 U199 ( .A(R1[29]), .B(R1[6]), .C(R1[4]), .Y(sigma1[19]) );
  XOR3X2 U200 ( .A(R1[28]), .B(R1[5]), .C(R1[3]), .Y(sigma1[18]) );
  XOR2X1 U201 ( .A(R14[6]), .B(R14[17]), .Y(sigma0[31]) );
  XOR3X2 U202 ( .A(R14[26]), .B(R14[30]), .C(R14[9]), .Y(sigma0[23]) );
  XOR3X2 U203 ( .A(R14[27]), .B(R14[31]), .C(R14[10]), .Y(sigma0[24]) );
  XOR3X2 U204 ( .A(R14[25]), .B(R14[29]), .C(R14[8]), .Y(sigma0[22]) );
  XOR3X2 U205 ( .A(R14[24]), .B(R14[28]), .C(R14[7]), .Y(sigma0[21]) );
  XOR3X2 U206 ( .A(R14[23]), .B(R14[27]), .C(R14[6]), .Y(sigma0[20]) );
  XOR3X2 U207 ( .A(R1[30]), .B(R1[7]), .C(R1[5]), .Y(sigma1[20]) );
  XOR3X2 U208 ( .A(R1[31]), .B(R1[8]), .C(R1[6]), .Y(sigma1[21]) );
  XOR2X1 U209 ( .A(R1[7]), .B(R1[9]), .Y(sigma1[22]) );
  XOR3X2 U210 ( .A(R14[13]), .B(R14[30]), .C(R14[2]), .Y(sigma0[27]) );
  XOR3X2 U211 ( .A(R14[12]), .B(R14[29]), .C(R14[1]), .Y(sigma0[26]) );
  XOR3X2 U212 ( .A(R14[11]), .B(R14[28]), .C(R14[0]), .Y(sigma0[25]) );
  XOR2X1 U213 ( .A(R1[12]), .B(R1[14]), .Y(sigma1[27]) );
  XOR3X2 U214 ( .A(R14[14]), .B(R14[31]), .C(R14[3]), .Y(sigma0[28]) );
  XOR2X1 U215 ( .A(R14[4]), .B(R14[15]), .Y(sigma0[29]) );
  XOR2X1 U216 ( .A(R14[5]), .B(R14[16]), .Y(sigma0[30]) );
  XOR2X1 U217 ( .A(R1[14]), .B(R1[16]), .Y(sigma1[29]) );
  XOR2X1 U218 ( .A(R1[15]), .B(R1[17]), .Y(sigma1[30]) );
endmodule


module hash_core_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  wire   [31:2] carry;

  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX4 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n18), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX4 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX4 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX4 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX4 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX4 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX4 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  NAND2X4 U1 ( .A(n1), .B(n16), .Y(carry[25]) );
  NAND2X2 U2 ( .A(A[20]), .B(n3), .Y(n6) );
  ADDFHX1 U3 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(n3) );
  NAND3X4 U4 ( .A(n12), .B(n10), .C(n11), .Y(carry[6]) );
  NAND2X2 U5 ( .A(B[5]), .B(carry[5]), .Y(n10) );
  NAND2X2 U6 ( .A(A[5]), .B(carry[5]), .Y(n11) );
  NAND2X2 U7 ( .A(B[20]), .B(carry[20]), .Y(n7) );
  INVX1 U8 ( .A(A[24]), .Y(n2) );
  NAND2X1 U9 ( .A(B[24]), .B(A[24]), .Y(n17) );
  AND2X2 U10 ( .A(B[0]), .B(A[0]), .Y(n18) );
  ADDFX2 U11 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(n4) );
  ADDFX2 U12 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(n13) );
  NAND2X1 U13 ( .A(A[5]), .B(B[5]), .Y(n12) );
  AND2X4 U14 ( .A(n17), .B(n15), .Y(n1) );
  NAND2BX4 U15 ( .AN(n2), .B(carry[24]), .Y(n15) );
  XOR2X1 U16 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U17 ( .A(A[20]), .B(B[20]), .Y(n5) );
  XOR2X1 U18 ( .A(n4), .B(n5), .Y(SUM[20]) );
  NAND2X4 U19 ( .A(B[20]), .B(A[20]), .Y(n8) );
  NAND3X4 U20 ( .A(n8), .B(n6), .C(n7), .Y(carry[21]) );
  XOR2X1 U21 ( .A(B[5]), .B(A[5]), .Y(n9) );
  XOR2X1 U22 ( .A(carry[5]), .B(n9), .Y(SUM[5]) );
  NAND2X1 U23 ( .A(B[24]), .B(carry[24]), .Y(n16) );
  XOR2X1 U24 ( .A(A[24]), .B(B[24]), .Y(n14) );
  XOR2X1 U25 ( .A(n13), .B(n14), .Y(SUM[24]) );
endmodule


module hash_core_DW01_add_1 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22;
  wire   [31:2] carry;

  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n17), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX4 U1_26 ( .A(A[26]), .B(B[26]), .CI(n16), .CO(carry[27]), .S(SUM[26])
         );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX4 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX4 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX4 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX4 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX4 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  NAND2X2 U1 ( .A(B[4]), .B(carry[4]), .Y(n6) );
  NAND3X4 U2 ( .A(n11), .B(n9), .C(n10), .Y(carry[19]) );
  NAND2X4 U3 ( .A(B[27]), .B(carry[27]), .Y(n20) );
  NAND2X4 U4 ( .A(A[18]), .B(n2), .Y(n9) );
  ADDFHX4 U5 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(n2) );
  NAND2X4 U6 ( .A(B[18]), .B(carry[18]), .Y(n10) );
  NAND2X4 U7 ( .A(A[25]), .B(carry[25]), .Y(n14) );
  ADDFHX2 U8 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(n1) );
  NAND2X1 U9 ( .A(B[18]), .B(A[18]), .Y(n11) );
  ADDFX2 U10 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(n3) );
  AND2X2 U11 ( .A(B[0]), .B(A[0]), .Y(n17) );
  XOR2X1 U12 ( .A(A[4]), .B(B[4]), .Y(n4) );
  XOR2X1 U13 ( .A(carry[4]), .B(n4), .Y(SUM[4]) );
  NAND2X4 U14 ( .A(A[4]), .B(n1), .Y(n5) );
  NAND2X4 U15 ( .A(B[4]), .B(A[4]), .Y(n7) );
  NAND3X4 U16 ( .A(n7), .B(n5), .C(n6), .Y(carry[5]) );
  XOR2X1 U17 ( .A(A[18]), .B(B[18]), .Y(n8) );
  XOR2X1 U18 ( .A(n3), .B(n8), .Y(SUM[18]) );
  AND2X4 U19 ( .A(n22), .B(n20), .Y(n12) );
  NAND2X2 U20 ( .A(n12), .B(n21), .Y(carry[28]) );
  NAND2X4 U21 ( .A(B[25]), .B(carry[25]), .Y(n13) );
  NAND2X4 U22 ( .A(A[25]), .B(B[25]), .Y(n15) );
  NAND3X4 U23 ( .A(n15), .B(n13), .C(n14), .Y(n16) );
  NAND2X1 U24 ( .A(A[27]), .B(B[27]), .Y(n22) );
  CMPR32X1 U25 ( .A(A[26]), .B(B[26]), .C(carry[26]), .CO(n18) );
  NAND2X1 U26 ( .A(A[27]), .B(carry[27]), .Y(n21) );
  XOR2X1 U27 ( .A(B[27]), .B(A[27]), .Y(n19) );
  XOR2X1 U28 ( .A(n18), .B(n19), .Y(SUM[27]) );
  XOR2X1 U29 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module hash_core_DW01_add_2 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [31:2] carry;

  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n16), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX4 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX4 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX4 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX4 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX4 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX4 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  XOR3X2 U1 ( .A(carry[22]), .B(B[22]), .C(A[22]), .Y(SUM[22]) );
  NAND2X2 U2 ( .A(A[22]), .B(carry[22]), .Y(n1) );
  NAND2X2 U3 ( .A(B[22]), .B(carry[22]), .Y(n2) );
  NAND2X1 U4 ( .A(B[22]), .B(A[22]), .Y(n3) );
  NAND3X2 U5 ( .A(n3), .B(n1), .C(n2), .Y(carry[23]) );
  NAND3X4 U6 ( .A(n9), .B(n10), .C(n11), .Y(carry[27]) );
  NAND2X4 U7 ( .A(A[26]), .B(carry[26]), .Y(n10) );
  ADDFHX2 U8 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(n4) );
  ADDFHX4 U9 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(n7) );
  NAND3X4 U10 ( .A(n14), .B(n13), .C(n15), .Y(carry[31]) );
  NAND2BX4 U11 ( .AN(n6), .B(n7), .Y(n14) );
  AND2X4 U12 ( .A(B[0]), .B(A[0]), .Y(n16) );
  NAND2X2 U13 ( .A(B[26]), .B(n4), .Y(n9) );
  INVX1 U14 ( .A(B[30]), .Y(n6) );
  NAND2X2 U15 ( .A(A[30]), .B(carry[30]), .Y(n13) );
  INVX1 U16 ( .A(A[31]), .Y(n5) );
  XNOR3X4 U17 ( .A(n5), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  XOR2XL U18 ( .A(B[26]), .B(A[26]), .Y(n8) );
  XOR2X1 U19 ( .A(carry[26]), .B(n8), .Y(SUM[26]) );
  NAND2X1 U20 ( .A(A[26]), .B(B[26]), .Y(n11) );
  XOR2X1 U21 ( .A(A[30]), .B(B[30]), .Y(n12) );
  XOR2X2 U22 ( .A(n7), .B(n12), .Y(SUM[30]) );
  NAND2XL U23 ( .A(B[30]), .B(A[30]), .Y(n15) );
  XOR2XL U24 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module hash_core_DW01_add_4 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2;
  wire   [31:1] carry;

  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX4 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX4 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX4 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX4 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX4 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX4 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX4 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX4 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  XOR2X4 U1 ( .A(carry[31]), .B(n1), .Y(SUM[31]) );
  CLKINVX3 U2 ( .A(n2), .Y(carry[1]) );
  NAND2X4 U3 ( .A(B[0]), .B(A[0]), .Y(n2) );
  XOR2XL U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U5 ( .A(A[31]), .B(B[31]), .Y(n1) );
endmodule


module hash_core_DW01_add_5 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;
  wire   [31:2] carry;

  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n15), .CO(carry[2]), .S(SUM[1]) );
  XOR3X4 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX4 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX4 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX4 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX4 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX4 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX4 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  XOR2X1 U1 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  NAND3X4 U2 ( .A(n13), .B(n12), .C(n14), .Y(carry[19]) );
  NAND3X4 U3 ( .A(n8), .B(n9), .C(n10), .Y(carry[17]) );
  NAND3X2 U4 ( .A(n5), .B(n3), .C(n4), .Y(carry[8]) );
  INVX1 U5 ( .A(A[18]), .Y(n1) );
  NAND2X1 U6 ( .A(B[7]), .B(carry[7]), .Y(n4) );
  ADDFX2 U7 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(n6) );
  NAND2X1 U8 ( .A(B[7]), .B(A[7]), .Y(n5) );
  NAND2X1 U9 ( .A(A[7]), .B(carry[7]), .Y(n3) );
  NAND2X2 U10 ( .A(B[16]), .B(carry[16]), .Y(n9) );
  NAND2X2 U11 ( .A(A[16]), .B(carry[16]), .Y(n8) );
  NAND2BX2 U12 ( .AN(n1), .B(carry[18]), .Y(n12) );
  NAND2X2 U13 ( .A(B[18]), .B(carry[18]), .Y(n13) );
  XOR2XL U14 ( .A(A[7]), .B(B[7]), .Y(n2) );
  XOR2X1 U15 ( .A(carry[7]), .B(n2), .Y(SUM[7]) );
  NAND2X1 U16 ( .A(B[16]), .B(A[16]), .Y(n10) );
  XOR2X1 U17 ( .A(A[16]), .B(B[16]), .Y(n7) );
  XOR2X1 U18 ( .A(n6), .B(n7), .Y(SUM[16]) );
  AND2X4 U19 ( .A(B[0]), .B(A[0]), .Y(n15) );
  NAND2X1 U20 ( .A(B[18]), .B(A[18]), .Y(n14) );
  XOR2X1 U21 ( .A(A[18]), .B(B[18]), .Y(n11) );
  XOR2X1 U22 ( .A(carry[18]), .B(n11), .Y(SUM[18]) );
endmodule


module hash_core_DW01_add_6 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [31:2] carry;

  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n24), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX4 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX4 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX4 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX4 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX4 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX4 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX4 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX4 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX4 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX4 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  NAND2X4 U1 ( .A(n10), .B(n8), .Y(n1) );
  NAND2X4 U2 ( .A(n2), .B(n9), .Y(carry[24]) );
  CLKINVX8 U3 ( .A(n1), .Y(n2) );
  NAND2X4 U4 ( .A(B[23]), .B(A[23]), .Y(n10) );
  NAND2X4 U5 ( .A(A[23]), .B(carry[23]), .Y(n8) );
  NAND2X4 U6 ( .A(n14), .B(n12), .Y(n3) );
  NAND2X4 U7 ( .A(n4), .B(n13), .Y(carry[11]) );
  CLKINVX8 U8 ( .A(n3), .Y(n4) );
  NAND2X4 U9 ( .A(B[10]), .B(A[10]), .Y(n14) );
  NAND2X4 U10 ( .A(A[10]), .B(carry[10]), .Y(n12) );
  ADDFHXL U11 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(n6) );
  ADDFHX4 U12 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(n5) );
  NAND3X4 U13 ( .A(n22), .B(n20), .C(n21), .Y(carry[18]) );
  NAND2X4 U14 ( .A(A[28]), .B(n5), .Y(n16) );
  NAND3X4 U15 ( .A(n18), .B(n16), .C(n17), .Y(carry[29]) );
  NAND2X4 U16 ( .A(B[28]), .B(carry[28]), .Y(n17) );
  NAND2X2 U17 ( .A(B[17]), .B(carry[17]), .Y(n21) );
  NAND2X1 U18 ( .A(B[23]), .B(carry[23]), .Y(n9) );
  NAND2X1 U19 ( .A(B[10]), .B(carry[10]), .Y(n13) );
  NAND2X1 U20 ( .A(B[28]), .B(A[28]), .Y(n18) );
  NAND2X1 U21 ( .A(B[17]), .B(A[17]), .Y(n22) );
  NAND2X2 U22 ( .A(A[17]), .B(carry[17]), .Y(n20) );
  XOR2X1 U23 ( .A(A[23]), .B(B[23]), .Y(n7) );
  XOR2X1 U24 ( .A(carry[23]), .B(n7), .Y(SUM[23]) );
  XOR2X1 U25 ( .A(A[10]), .B(B[10]), .Y(n11) );
  XOR2X1 U26 ( .A(carry[10]), .B(n11), .Y(SUM[10]) );
  XOR2XL U27 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  AND2X4 U28 ( .A(A[0]), .B(B[0]), .Y(n24) );
  XOR2X1 U29 ( .A(A[28]), .B(B[28]), .Y(n15) );
  XOR2X1 U30 ( .A(n6), .B(n15), .Y(SUM[28]) );
  XOR2X1 U31 ( .A(A[17]), .B(B[17]), .Y(n19) );
  XOR2X1 U32 ( .A(carry[17]), .B(n19), .Y(SUM[17]) );
  XOR2X4 U33 ( .A(carry[31]), .B(n23), .Y(SUM[31]) );
  XOR2X1 U34 ( .A(A[31]), .B(B[31]), .Y(n23) );
endmodule


module hash_core_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module hash_core_DW01_add_16 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232;

  NOR2BX2 U2 ( .AN(n210), .B(n211), .Y(n204) );
  CLKINVX3 U3 ( .A(n212), .Y(n211) );
  CLKINVX3 U4 ( .A(n163), .Y(n162) );
  OAI21X4 U5 ( .A0(n73), .A1(n74), .B0(n75), .Y(n7) );
  NOR2X4 U6 ( .A(A[25]), .B(B[25]), .Y(n91) );
  OR2X2 U7 ( .A(n229), .B(n230), .Y(n1) );
  NAND2X2 U8 ( .A(n1), .B(n54), .Y(n184) );
  XOR2X4 U9 ( .A(n97), .B(n98), .Y(SUM[27]) );
  AOI21X4 U10 ( .A0(n144), .A1(n145), .B0(n146), .Y(n135) );
  AND2X4 U11 ( .A(n75), .B(n76), .Y(n22) );
  NAND2X4 U12 ( .A(B[28]), .B(A[28]), .Y(n75) );
  NAND2X4 U13 ( .A(n84), .B(n106), .Y(n104) );
  AND2X2 U14 ( .A(n106), .B(n108), .Y(n109) );
  NAND2X1 U15 ( .A(B[24]), .B(A[24]), .Y(n106) );
  INVX4 U16 ( .A(n129), .Y(n117) );
  NAND4BBX2 U17 ( .AN(n46), .BN(n24), .C(n44), .D(n38), .Y(n187) );
  CLKINVX3 U18 ( .A(n172), .Y(n171) );
  OR2X2 U19 ( .A(A[9]), .B(B[9]), .Y(n208) );
  OR2X2 U20 ( .A(A[6]), .B(B[6]), .Y(n44) );
  OAI21X2 U21 ( .A0(n65), .A1(n66), .B0(n67), .Y(n64) );
  NOR2X2 U22 ( .A(n68), .B(n65), .Y(n62) );
  NAND2X2 U23 ( .A(B[20]), .B(n4), .Y(n118) );
  NAND2X1 U24 ( .A(n165), .B(n149), .Y(n163) );
  NAND2X1 U25 ( .A(B[13]), .B(A[13]), .Y(n174) );
  NAND2X2 U26 ( .A(B[10]), .B(A[10]), .Y(n210) );
  NAND2X1 U27 ( .A(n30), .B(n213), .Y(n221) );
  NAND2X1 U28 ( .A(B[9]), .B(A[9]), .Y(n28) );
  INVX1 U29 ( .A(n48), .Y(n45) );
  NAND2X1 U30 ( .A(B[6]), .B(A[6]), .Y(n41) );
  INVX1 U31 ( .A(n58), .Y(n231) );
  INVX1 U32 ( .A(n147), .Y(n146) );
  XOR2X1 U33 ( .A(n194), .B(n195), .Y(SUM[14]) );
  OAI21X2 U34 ( .A0(n203), .A1(n178), .B0(n183), .Y(n201) );
  XOR2X1 U35 ( .A(n159), .B(n161), .Y(SUM[18]) );
  NOR2BX1 U36 ( .AN(n94), .B(n2), .Y(n101) );
  NAND2X1 U37 ( .A(B[15]), .B(A[15]), .Y(n172) );
  NOR2X4 U38 ( .A(A[26]), .B(B[26]), .Y(n2) );
  OR2X2 U39 ( .A(A[25]), .B(B[25]), .Y(n103) );
  INVX3 U40 ( .A(n190), .Y(n176) );
  NAND3X2 U41 ( .A(n103), .B(n3), .C(n96), .Y(n85) );
  NOR2BXL U42 ( .AN(n116), .B(n25), .Y(n125) );
  OR2X1 U43 ( .A(A[26]), .B(B[26]), .Y(n3) );
  NOR2X2 U44 ( .A(A[13]), .B(B[13]), .Y(n23) );
  NAND2X4 U45 ( .A(B[26]), .B(A[26]), .Y(n94) );
  NAND2X1 U46 ( .A(B[5]), .B(A[5]), .Y(n47) );
  BUFX3 U47 ( .A(A[20]), .Y(n4) );
  NAND2X2 U48 ( .A(B[21]), .B(A[21]), .Y(n119) );
  NAND3X4 U49 ( .A(n129), .B(n122), .C(n123), .Y(n5) );
  NAND3XL U50 ( .A(n129), .B(n122), .C(n123), .Y(n111) );
  INVX4 U51 ( .A(n116), .Y(n115) );
  OAI21X2 U52 ( .A0(n220), .A1(n29), .B0(n28), .Y(n216) );
  NAND2X1 U53 ( .A(B[29]), .B(A[29]), .Y(n72) );
  NAND2X1 U54 ( .A(A[29]), .B(B[29]), .Y(n66) );
  OAI21X4 U55 ( .A0(n110), .A1(n5), .B0(n112), .Y(n6) );
  OAI21XL U56 ( .A0(n111), .A1(n110), .B0(n112), .Y(n107) );
  NAND4BBX4 U57 ( .AN(n33), .BN(n29), .C(n207), .D(n206), .Y(n178) );
  AOI21X2 U58 ( .A0(n179), .A1(n184), .B0(n185), .Y(n182) );
  XOR2X2 U59 ( .A(n156), .B(n157), .Y(SUM[19]) );
  AOI21X2 U60 ( .A0(n158), .A1(n159), .B0(n160), .Y(n157) );
  NAND2X2 U61 ( .A(B[19]), .B(A[19]), .Y(n147) );
  INVX2 U62 ( .A(n75), .Y(n19) );
  OAI21X4 U63 ( .A0(n99), .A1(n2), .B0(n94), .Y(n97) );
  OAI21X2 U64 ( .A0(n24), .A1(n227), .B0(n50), .Y(n48) );
  OAI2BB1X4 U65 ( .A0N(n204), .A1N(n205), .B0(n206), .Y(n183) );
  NAND2XL U66 ( .A(n22), .B(n74), .Y(n10) );
  NAND2X2 U67 ( .A(n8), .B(n9), .Y(n11) );
  NAND2X2 U68 ( .A(n10), .B(n11), .Y(SUM[28]) );
  INVXL U69 ( .A(n22), .Y(n8) );
  INVXL U70 ( .A(n74), .Y(n9) );
  INVX8 U71 ( .A(n83), .Y(n74) );
  NAND2X4 U72 ( .A(n60), .B(n13), .Y(n14) );
  NAND2X2 U73 ( .A(n61), .B(n12), .Y(n15) );
  NAND2X4 U74 ( .A(n14), .B(n15), .Y(SUM[31]) );
  CLKINVX3 U75 ( .A(n60), .Y(n12) );
  INVX4 U76 ( .A(n61), .Y(n13) );
  XNOR2X2 U77 ( .A(B[31]), .B(A[31]), .Y(n60) );
  XOR2X4 U78 ( .A(n20), .B(n70), .Y(SUM[30]) );
  XNOR2X1 U79 ( .A(B[30]), .B(A[30]), .Y(n20) );
  INVX2 U80 ( .A(n30), .Y(n203) );
  OAI21X2 U81 ( .A0(n227), .A1(n187), .B0(n186), .Y(n30) );
  OAI21X4 U82 ( .A0(n126), .A1(n121), .B0(n120), .Y(n124) );
  INVX4 U83 ( .A(n127), .Y(n126) );
  NAND2X4 U84 ( .A(B[7]), .B(A[7]), .Y(n36) );
  OAI21X2 U85 ( .A0(n162), .A1(n148), .B0(n150), .Y(n159) );
  NAND2X1 U86 ( .A(n110), .B(n118), .Y(n130) );
  OAI2BB1X4 U87 ( .A0N(n129), .A1N(n130), .B0(n119), .Y(n127) );
  NOR2X2 U88 ( .A(n196), .B(n23), .Y(n16) );
  INVXL U89 ( .A(n174), .Y(n17) );
  OR2X4 U90 ( .A(n16), .B(n17), .Y(n194) );
  INVX2 U91 ( .A(n197), .Y(n196) );
  INVX4 U92 ( .A(n194), .Y(n193) );
  NAND2X1 U93 ( .A(B[17]), .B(A[17]), .Y(n150) );
  OR2X1 U94 ( .A(A[2]), .B(B[2]), .Y(n78) );
  NAND2BX4 U95 ( .AN(n180), .B(n181), .Y(n167) );
  NAND2X2 U96 ( .A(A[24]), .B(B[24]), .Y(n92) );
  NAND2X2 U97 ( .A(B[27]), .B(A[27]), .Y(n90) );
  OAI21X4 U98 ( .A0(n182), .A1(n178), .B0(n183), .Y(n181) );
  INVX4 U99 ( .A(n100), .Y(n99) );
  OAI21X2 U100 ( .A0(n193), .A1(n177), .B0(n175), .Y(n191) );
  INVX2 U101 ( .A(n224), .Y(n46) );
  NOR2BXL U102 ( .AN(n172), .B(n176), .Y(n192) );
  OAI21XL U103 ( .A0(n45), .A1(n46), .B0(n47), .Y(n42) );
  OR2X4 U104 ( .A(A[7]), .B(B[7]), .Y(n38) );
  NOR2X1 U105 ( .A(A[4]), .B(B[4]), .Y(n24) );
  OR2X2 U106 ( .A(n4), .B(B[20]), .Y(n133) );
  NAND2X1 U107 ( .A(B[2]), .B(A[2]), .Y(n58) );
  OAI21X2 U108 ( .A0(n199), .A1(n200), .B0(n173), .Y(n197) );
  INVX2 U109 ( .A(n201), .Y(n200) );
  OAI2BB1X2 U110 ( .A0N(n222), .A1N(n223), .B0(n38), .Y(n186) );
  NAND2XL U111 ( .A(n147), .B(n152), .Y(n156) );
  INVXL U112 ( .A(n151), .Y(n160) );
  NAND2XL U113 ( .A(n221), .B(n32), .Y(n26) );
  AOI21XL U114 ( .A0(n207), .A1(n216), .B0(n217), .Y(n215) );
  AOI21XL U115 ( .A0(n76), .A1(n83), .B0(n19), .Y(n18) );
  OAI211X2 U116 ( .A0(n23), .A1(n173), .B0(n174), .C0(n175), .Y(n170) );
  NOR2BXL U117 ( .AN(n28), .B(n29), .Y(n27) );
  NAND4BX2 U118 ( .AN(n23), .B(n188), .C(n189), .D(n190), .Y(n180) );
  NOR2BXL U119 ( .AN(n90), .B(n95), .Y(n98) );
  NOR2BXL U120 ( .AN(n120), .B(n121), .Y(n128) );
  INVXL U121 ( .A(n188), .Y(n199) );
  AND2X1 U122 ( .A(n118), .B(n133), .Y(n134) );
  INVXL U123 ( .A(n44), .Y(n40) );
  NOR2BXL U124 ( .AN(n47), .B(n46), .Y(n49) );
  AND2X1 U125 ( .A(n149), .B(n142), .Y(n166) );
  INVXL U126 ( .A(n228), .Y(n55) );
  NOR2BXL U127 ( .AN(n81), .B(n154), .Y(n153) );
  INVXL U128 ( .A(n155), .Y(n80) );
  NAND2X4 U129 ( .A(B[11]), .B(A[11]), .Y(n212) );
  NAND2X2 U130 ( .A(B[14]), .B(A[14]), .Y(n175) );
  NAND2XL U131 ( .A(B[3]), .B(A[3]), .Y(n54) );
  OR2X4 U132 ( .A(A[16]), .B(B[16]), .Y(n142) );
  NAND2XL U133 ( .A(B[1]), .B(A[1]), .Y(n81) );
  NOR2BX1 U134 ( .AN(n155), .B(n21), .Y(SUM[0]) );
  NOR2XL U135 ( .A(A[0]), .B(B[0]), .Y(n21) );
  INVX1 U136 ( .A(n186), .Y(n185) );
  INVX1 U137 ( .A(n187), .Y(n179) );
  INVX1 U138 ( .A(n184), .Y(n227) );
  INVX1 U139 ( .A(n59), .Y(n56) );
  INVX1 U140 ( .A(n208), .Y(n29) );
  INVX1 U141 ( .A(n90), .Y(n89) );
  NOR2BXL U142 ( .AN(n119), .B(n117), .Y(n131) );
  NAND3X2 U143 ( .A(n207), .B(n208), .C(n209), .Y(n205) );
  INVX1 U144 ( .A(n213), .Y(n33) );
  NAND3X1 U145 ( .A(n224), .B(n44), .C(n225), .Y(n223) );
  NOR2BX1 U146 ( .AN(n41), .B(n226), .Y(n222) );
  NAND2X1 U147 ( .A(n47), .B(n50), .Y(n225) );
  NOR2BXL U148 ( .AN(n175), .B(n177), .Y(n195) );
  XOR2X1 U149 ( .A(n163), .B(n164), .Y(SUM[17]) );
  NOR2BXL U150 ( .AN(n150), .B(n148), .Y(n164) );
  NAND2X1 U151 ( .A(n28), .B(n32), .Y(n209) );
  INVX1 U152 ( .A(n36), .Y(n226) );
  XOR2X1 U153 ( .A(n82), .B(n18), .Y(SUM[29]) );
  XOR2X1 U154 ( .A(n124), .B(n125), .Y(SUM[23]) );
  XOR2X1 U155 ( .A(n127), .B(n128), .Y(SUM[22]) );
  NOR2BXL U156 ( .AN(n93), .B(n91), .Y(n105) );
  NAND2XL U157 ( .A(n69), .B(n72), .Y(n82) );
  XOR2X1 U158 ( .A(n100), .B(n101), .Y(SUM[26]) );
  INVX4 U159 ( .A(n152), .Y(n141) );
  NAND2XL U160 ( .A(n142), .B(n143), .Y(n137) );
  INVX8 U161 ( .A(n122), .Y(n121) );
  INVX1 U162 ( .A(n26), .Y(n220) );
  NAND2X1 U163 ( .A(n78), .B(n228), .Y(n230) );
  NOR2X1 U164 ( .A(n231), .B(n232), .Y(n229) );
  INVX1 U165 ( .A(n210), .Y(n217) );
  NOR2BX1 U166 ( .AN(n174), .B(n23), .Y(n198) );
  INVX1 U167 ( .A(n79), .Y(n154) );
  OAI21XL U168 ( .A0(n154), .A1(n155), .B0(n81), .Y(n232) );
  XOR2X1 U169 ( .A(n201), .B(n202), .Y(SUM[12]) );
  NOR2BX1 U170 ( .AN(n173), .B(n199), .Y(n202) );
  XOR2X1 U171 ( .A(n216), .B(n218), .Y(SUM[10]) );
  NOR2BX1 U172 ( .AN(n210), .B(n219), .Y(n218) );
  INVX1 U173 ( .A(n207), .Y(n219) );
  XOR2X1 U174 ( .A(n26), .B(n27), .Y(SUM[9]) );
  NAND2XL U175 ( .A(n206), .B(n212), .Y(n214) );
  XOR2X1 U176 ( .A(n30), .B(n31), .Y(SUM[8]) );
  NOR2BX1 U177 ( .AN(n32), .B(n33), .Y(n31) );
  XOR2X1 U178 ( .A(n48), .B(n49), .Y(SUM[5]) );
  XOR2X1 U179 ( .A(n42), .B(n43), .Y(SUM[6]) );
  NOR2BX1 U180 ( .AN(n41), .B(n40), .Y(n43) );
  INVX1 U181 ( .A(n38), .Y(n37) );
  XOR2X1 U182 ( .A(n34), .B(n35), .Y(SUM[7]) );
  OAI21XL U183 ( .A0(n39), .A1(n40), .B0(n41), .Y(n34) );
  NOR2BX1 U184 ( .AN(n36), .B(n37), .Y(n35) );
  INVX1 U185 ( .A(n42), .Y(n39) );
  INVX1 U186 ( .A(n78), .Y(n57) );
  XOR2X1 U187 ( .A(n80), .B(n153), .Y(SUM[1]) );
  XOR2X1 U188 ( .A(n59), .B(n77), .Y(SUM[2]) );
  NOR2BX1 U189 ( .AN(n58), .B(n57), .Y(n77) );
  OAI2BB1X1 U190 ( .A0N(n79), .A1N(n80), .B0(n81), .Y(n59) );
  XOR2X1 U191 ( .A(n184), .B(n51), .Y(SUM[4]) );
  NOR2BX1 U192 ( .AN(n50), .B(n24), .Y(n51) );
  XOR2X1 U193 ( .A(n52), .B(n53), .Y(SUM[3]) );
  NOR2BX1 U194 ( .AN(n54), .B(n55), .Y(n53) );
  OAI21XL U195 ( .A0(n56), .A1(n57), .B0(n58), .Y(n52) );
  NAND2X2 U196 ( .A(B[12]), .B(A[12]), .Y(n173) );
  NAND2X1 U197 ( .A(B[8]), .B(A[8]), .Y(n32) );
  NAND2X2 U198 ( .A(B[22]), .B(A[22]), .Y(n120) );
  NAND2X2 U199 ( .A(B[18]), .B(A[18]), .Y(n151) );
  OR2X2 U200 ( .A(A[12]), .B(B[12]), .Y(n188) );
  OR2X2 U201 ( .A(A[24]), .B(B[24]), .Y(n108) );
  OR2X2 U202 ( .A(A[8]), .B(B[8]), .Y(n213) );
  NAND2X2 U203 ( .A(A[30]), .B(B[30]), .Y(n67) );
  OR2X2 U204 ( .A(A[5]), .B(B[5]), .Y(n224) );
  XOR2X1 U205 ( .A(n191), .B(n192), .Y(SUM[15]) );
  XOR2X1 U206 ( .A(n130), .B(n131), .Y(SUM[21]) );
  NAND2X1 U207 ( .A(B[4]), .B(A[4]), .Y(n50) );
  OR2X2 U208 ( .A(A[3]), .B(B[3]), .Y(n228) );
  OR2X2 U209 ( .A(A[1]), .B(B[1]), .Y(n79) );
  XOR2X1 U210 ( .A(n214), .B(n215), .Y(SUM[11]) );
  XOR2X1 U211 ( .A(n197), .B(n198), .Y(SUM[13]) );
  NAND2X1 U212 ( .A(B[0]), .B(A[0]), .Y(n155) );
  NAND2X4 U213 ( .A(n167), .B(n168), .Y(n138) );
  NAND2X2 U214 ( .A(B[23]), .B(A[23]), .Y(n116) );
  NOR2BX1 U215 ( .AN(n151), .B(n140), .Y(n161) );
  INVX4 U216 ( .A(n158), .Y(n140) );
  NAND2X1 U217 ( .A(n138), .B(n142), .Y(n165) );
  NOR2X4 U218 ( .A(B[23]), .B(A[23]), .Y(n25) );
  XOR2X1 U219 ( .A(n138), .B(n166), .Y(SUM[16]) );
  CLKINVX8 U220 ( .A(n96), .Y(n95) );
  XOR2X1 U221 ( .A(n132), .B(n134), .Y(SUM[20]) );
  XOR2X1 U222 ( .A(n104), .B(n105), .Y(SUM[25]) );
  XOR2X1 U223 ( .A(n107), .B(n109), .Y(SUM[24]) );
  AOI21X4 U224 ( .A0(n62), .A1(n7), .B0(n64), .Y(n61) );
  NOR2X4 U225 ( .A(A[30]), .B(B[30]), .Y(n65) );
  CLKINVX3 U226 ( .A(n69), .Y(n68) );
  AOI21X4 U227 ( .A0(n69), .A1(n63), .B0(n71), .Y(n70) );
  CLKINVX3 U228 ( .A(n72), .Y(n71) );
  OAI21X4 U229 ( .A0(n73), .A1(n74), .B0(n75), .Y(n63) );
  CLKINVX3 U230 ( .A(n76), .Y(n73) );
  OR2X4 U231 ( .A(A[29]), .B(B[29]), .Y(n69) );
  OAI21X4 U232 ( .A0(n84), .A1(n85), .B0(n86), .Y(n83) );
  AOI21X4 U233 ( .A0(n87), .A1(n88), .B0(n89), .Y(n86) );
  OAI211X2 U234 ( .A0(n91), .A1(n92), .B0(n93), .C0(n94), .Y(n88) );
  NOR2X4 U235 ( .A(n95), .B(n2), .Y(n87) );
  OR2X4 U236 ( .A(A[28]), .B(B[28]), .Y(n76) );
  OR2X4 U237 ( .A(A[27]), .B(B[27]), .Y(n96) );
  NAND2X4 U238 ( .A(n102), .B(n93), .Y(n100) );
  NAND2X4 U239 ( .A(n103), .B(n104), .Y(n102) );
  NAND2X4 U240 ( .A(B[25]), .B(A[25]), .Y(n93) );
  NAND2X4 U241 ( .A(n6), .B(n108), .Y(n84) );
  AOI21X4 U242 ( .A0(n113), .A1(n114), .B0(n115), .Y(n112) );
  OAI211X2 U243 ( .A0(n117), .A1(n118), .B0(n119), .C0(n120), .Y(n114) );
  NOR2X4 U244 ( .A(n25), .B(n121), .Y(n113) );
  OR2X4 U245 ( .A(A[23]), .B(B[23]), .Y(n123) );
  OR2X4 U246 ( .A(A[22]), .B(B[22]), .Y(n122) );
  OR2X4 U247 ( .A(A[21]), .B(B[21]), .Y(n129) );
  NAND2X4 U248 ( .A(n132), .B(n133), .Y(n110) );
  NAND2X4 U249 ( .A(n135), .B(n136), .Y(n132) );
  NAND3BX4 U250 ( .AN(n137), .B(n138), .C(n139), .Y(n136) );
  NOR2X4 U251 ( .A(n140), .B(n141), .Y(n139) );
  OAI211X2 U252 ( .A0(n148), .A1(n149), .B0(n150), .C0(n151), .Y(n145) );
  NOR2X4 U253 ( .A(n141), .B(n140), .Y(n144) );
  OR2X4 U254 ( .A(A[19]), .B(B[19]), .Y(n152) );
  OR2X4 U255 ( .A(A[18]), .B(B[18]), .Y(n158) );
  CLKINVX3 U256 ( .A(n143), .Y(n148) );
  OR2X4 U257 ( .A(A[17]), .B(B[17]), .Y(n143) );
  NAND2X4 U258 ( .A(B[16]), .B(A[16]), .Y(n149) );
  AOI21X4 U259 ( .A0(n169), .A1(n170), .B0(n171), .Y(n168) );
  NOR2X4 U260 ( .A(n176), .B(n177), .Y(n169) );
  OR2X4 U261 ( .A(A[15]), .B(B[15]), .Y(n190) );
  CLKINVX3 U262 ( .A(n189), .Y(n177) );
  OR2X4 U263 ( .A(A[14]), .B(B[14]), .Y(n189) );
  OR2X4 U264 ( .A(A[11]), .B(B[11]), .Y(n206) );
  OR2X4 U265 ( .A(A[10]), .B(B[10]), .Y(n207) );
endmodule


module hash_core_DW01_add_18 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240;

  AOI21X4 U2 ( .A0(n153), .A1(n154), .B0(n155), .Y(n144) );
  NOR2X4 U3 ( .A(n150), .B(n149), .Y(n153) );
  NAND2X2 U4 ( .A(B[15]), .B(A[15]), .Y(n181) );
  NAND2X4 U5 ( .A(n89), .B(n114), .Y(n112) );
  NAND2X1 U6 ( .A(n133), .B(n2), .Y(n3) );
  NAND2X2 U7 ( .A(n1), .B(n134), .Y(n4) );
  NAND2X2 U8 ( .A(n3), .B(n4), .Y(SUM[23]) );
  CLKINVX3 U9 ( .A(n133), .Y(n1) );
  INVXL U10 ( .A(n134), .Y(n2) );
  NAND2X2 U11 ( .A(n17), .B(n9), .Y(n133) );
  NOR2BX1 U12 ( .AN(n124), .B(n129), .Y(n134) );
  NAND2X2 U13 ( .A(n88), .B(n6), .Y(n7) );
  NAND2XL U14 ( .A(n5), .B(n77), .Y(n8) );
  NAND2X2 U15 ( .A(n7), .B(n8), .Y(SUM[28]) );
  INVX1 U16 ( .A(n88), .Y(n5) );
  INVXL U17 ( .A(n77), .Y(n6) );
  NAND2X2 U18 ( .A(n78), .B(n79), .Y(n88) );
  OR2X4 U19 ( .A(A[27]), .B(B[27]), .Y(n104) );
  NAND2X4 U20 ( .A(B[20]), .B(A[20]), .Y(n126) );
  INVX2 U21 ( .A(n156), .Y(n155) );
  AOI21X2 U22 ( .A0(n79), .A1(n86), .B0(n87), .Y(n85) );
  OAI21X2 U23 ( .A0(n205), .A1(n24), .B0(n183), .Y(n203) );
  INVX4 U24 ( .A(n206), .Y(n205) );
  NOR2BX4 U25 ( .AN(n12), .B(n102), .Y(n113) );
  DLY1X1 U26 ( .A(n98), .Y(n12) );
  AOI21X4 U27 ( .A0(n65), .A1(n72), .B0(n74), .Y(n73) );
  INVX4 U28 ( .A(n193), .Y(n235) );
  AOI21X2 U29 ( .A0(n188), .A1(n193), .B0(n194), .Y(n191) );
  OAI21X4 U30 ( .A0(n237), .A1(n238), .B0(n56), .Y(n193) );
  XNOR2X2 U31 ( .A(n23), .B(n85), .Y(SUM[29]) );
  NAND2X4 U32 ( .A(n21), .B(n22), .Y(SUM[31]) );
  NAND3X2 U33 ( .A(n111), .B(n10), .C(n104), .Y(n90) );
  CLKINVX4 U34 ( .A(n101), .Y(n10) );
  NOR2X2 U35 ( .A(n70), .B(n71), .Y(n64) );
  INVX4 U36 ( .A(n152), .Y(n157) );
  OAI2BB1X2 U37 ( .A0N(n230), .A1N(n231), .B0(n40), .Y(n195) );
  OR2X2 U38 ( .A(A[12]), .B(B[12]), .Y(n197) );
  NOR2X2 U39 ( .A(A[30]), .B(B[30]), .Y(n71) );
  NAND2X2 U40 ( .A(B[30]), .B(A[30]), .Y(n69) );
  NOR2X2 U41 ( .A(A[30]), .B(B[30]), .Y(n67) );
  CLKINVX3 U42 ( .A(n95), .Y(n94) );
  NAND2X1 U43 ( .A(A[25]), .B(B[25]), .Y(n98) );
  NAND3X1 U44 ( .A(n216), .B(n217), .C(n218), .Y(n214) );
  INVX1 U45 ( .A(n181), .Y(n180) );
  INVX4 U46 ( .A(n131), .Y(n130) );
  CLKINVX3 U47 ( .A(n199), .Y(n185) );
  NAND2X1 U48 ( .A(B[12]), .B(A[12]), .Y(n182) );
  CLKINVX3 U49 ( .A(n138), .Y(n125) );
  INVX1 U50 ( .A(n75), .Y(n74) );
  NAND2X1 U51 ( .A(B[29]), .B(A[29]), .Y(n75) );
  CLKINVX4 U52 ( .A(n104), .Y(n100) );
  OR2X2 U53 ( .A(A[25]), .B(B[25]), .Y(n111) );
  OAI21XL U54 ( .A0(n47), .A1(n48), .B0(n49), .Y(n44) );
  OR2X2 U55 ( .A(n171), .B(n157), .Y(n18) );
  CLKINVX3 U56 ( .A(n172), .Y(n171) );
  OR2X2 U57 ( .A(A[20]), .B(B[20]), .Y(n142) );
  INVX1 U58 ( .A(n28), .Y(n228) );
  OAI21X1 U59 ( .A0(n202), .A1(n186), .B0(n184), .Y(n200) );
  INVX4 U60 ( .A(n198), .Y(n186) );
  NAND2BX4 U61 ( .AN(n189), .B(n190), .Y(n176) );
  NAND2XL U62 ( .A(n147), .B(n151), .Y(n174) );
  OR2X2 U63 ( .A(A[8]), .B(B[8]), .Y(n221) );
  DLY1X1 U64 ( .A(n128), .Y(n9) );
  NOR2BX1 U65 ( .AN(n9), .B(n130), .Y(n137) );
  INVX8 U66 ( .A(n161), .Y(n150) );
  CLKINVX3 U67 ( .A(n62), .Y(n19) );
  INVX8 U68 ( .A(n103), .Y(n101) );
  NAND2BX4 U69 ( .AN(A[26]), .B(n11), .Y(n103) );
  CLKINVX20 U70 ( .A(B[26]), .Y(n11) );
  INVX1 U71 ( .A(A[30]), .Y(n14) );
  NAND2X4 U72 ( .A(B[26]), .B(A[26]), .Y(n99) );
  NAND2X2 U73 ( .A(n111), .B(n112), .Y(n110) );
  INVX4 U74 ( .A(n111), .Y(n102) );
  NAND2X1 U75 ( .A(A[29]), .B(B[29]), .Y(n68) );
  OAI21X4 U76 ( .A0(n107), .A1(n101), .B0(n99), .Y(n105) );
  INVX2 U77 ( .A(n108), .Y(n107) );
  NAND2X2 U78 ( .A(n110), .B(n12), .Y(n108) );
  XOR2X2 U79 ( .A(n112), .B(n113), .Y(SUM[25]) );
  NAND2X1 U80 ( .A(B[30]), .B(n14), .Y(n15) );
  NAND2XL U81 ( .A(n13), .B(A[30]), .Y(n16) );
  NAND2X2 U82 ( .A(n15), .B(n16), .Y(n26) );
  INVX1 U83 ( .A(B[30]), .Y(n13) );
  OR2X4 U84 ( .A(n135), .B(n130), .Y(n17) );
  INVX3 U85 ( .A(n136), .Y(n135) );
  NAND2X2 U86 ( .A(n18), .B(n159), .Y(n168) );
  AOI21X2 U87 ( .A0(n167), .A1(n168), .B0(n169), .Y(n166) );
  NAND2X2 U88 ( .A(n62), .B(n20), .Y(n21) );
  NAND2X2 U89 ( .A(n63), .B(n19), .Y(n22) );
  INVX4 U90 ( .A(n63), .Y(n20) );
  XNOR2X2 U91 ( .A(B[31]), .B(A[31]), .Y(n62) );
  OAI21X2 U92 ( .A0(n235), .A1(n196), .B0(n195), .Y(n32) );
  NOR2X2 U93 ( .A(A[25]), .B(B[25]), .Y(n96) );
  OR2X4 U94 ( .A(A[5]), .B(B[5]), .Y(n232) );
  NAND2X4 U95 ( .A(B[5]), .B(A[5]), .Y(n49) );
  NAND2X2 U96 ( .A(B[24]), .B(A[24]), .Y(n114) );
  OR2X4 U97 ( .A(A[24]), .B(B[24]), .Y(n116) );
  NAND2X2 U98 ( .A(n118), .B(n126), .Y(n139) );
  NAND2X2 U99 ( .A(B[6]), .B(A[6]), .Y(n43) );
  NAND2X4 U100 ( .A(B[7]), .B(A[7]), .Y(n38) );
  NAND2X1 U101 ( .A(B[17]), .B(A[17]), .Y(n159) );
  NAND2X2 U102 ( .A(B[13]), .B(A[13]), .Y(n183) );
  NAND2X2 U103 ( .A(B[8]), .B(A[8]), .Y(n34) );
  NOR2X2 U104 ( .A(A[13]), .B(B[13]), .Y(n24) );
  OR2X2 U105 ( .A(A[7]), .B(B[7]), .Y(n40) );
  NAND4BBX2 U106 ( .AN(n48), .BN(n25), .C(n46), .D(n40), .Y(n196) );
  OR2X1 U107 ( .A(A[2]), .B(B[2]), .Y(n81) );
  CLKINVX3 U108 ( .A(n60), .Y(n239) );
  NAND2X2 U109 ( .A(B[9]), .B(A[9]), .Y(n30) );
  NOR2X1 U110 ( .A(A[4]), .B(B[4]), .Y(n25) );
  OAI21X2 U111 ( .A0(n191), .A1(n187), .B0(n192), .Y(n190) );
  INVX2 U112 ( .A(n232), .Y(n48) );
  OAI21XL U113 ( .A0(n228), .A1(n31), .B0(n30), .Y(n224) );
  NOR2BX1 U114 ( .AN(n182), .B(n208), .Y(n211) );
  NAND2X1 U115 ( .A(B[2]), .B(A[2]), .Y(n60) );
  OAI21X2 U116 ( .A0(n212), .A1(n187), .B0(n192), .Y(n210) );
  INVX2 U117 ( .A(n203), .Y(n202) );
  OAI21X2 U118 ( .A0(n208), .A1(n209), .B0(n182), .Y(n206) );
  INVX2 U119 ( .A(n210), .Y(n209) );
  INVXL U120 ( .A(n160), .Y(n169) );
  OAI2BB1X2 U121 ( .A0N(n138), .A1N(n139), .B0(n127), .Y(n136) );
  AND2X1 U122 ( .A(n72), .B(n75), .Y(n23) );
  AND2X2 U123 ( .A(n219), .B(n220), .Y(n213) );
  NAND2X2 U124 ( .A(n174), .B(n158), .Y(n172) );
  NOR2BXL U125 ( .AN(n30), .B(n31), .Y(n29) );
  NOR2BXL U126 ( .AN(n34), .B(n35), .Y(n33) );
  AND2X1 U127 ( .A(n158), .B(n151), .Y(n175) );
  AND2X1 U128 ( .A(n114), .B(n116), .Y(n117) );
  INVXL U129 ( .A(n46), .Y(n42) );
  AND2X1 U130 ( .A(n126), .B(n142), .Y(n143) );
  INVXL U131 ( .A(n236), .Y(n57) );
  NOR2BXL U132 ( .AN(n84), .B(n163), .Y(n162) );
  INVXL U133 ( .A(n164), .Y(n83) );
  NAND2X2 U134 ( .A(B[10]), .B(A[10]), .Y(n219) );
  OR2X4 U135 ( .A(A[9]), .B(B[9]), .Y(n217) );
  NAND2X2 U136 ( .A(B[14]), .B(A[14]), .Y(n184) );
  NAND2XL U137 ( .A(B[1]), .B(A[1]), .Y(n84) );
  NAND2XL U138 ( .A(B[3]), .B(A[3]), .Y(n56) );
  NOR2XL U139 ( .A(A[0]), .B(B[0]), .Y(n27) );
  INVX1 U140 ( .A(n32), .Y(n212) );
  INVX1 U141 ( .A(n195), .Y(n194) );
  INVX1 U142 ( .A(n196), .Y(n188) );
  XOR2X1 U143 ( .A(n108), .B(n109), .Y(SUM[26]) );
  INVX1 U144 ( .A(n61), .Y(n58) );
  INVX1 U145 ( .A(n217), .Y(n31) );
  INVX1 U146 ( .A(n197), .Y(n208) );
  INVXL U147 ( .A(n78), .Y(n87) );
  NOR2BXL U148 ( .AN(n127), .B(n125), .Y(n140) );
  OAI2BB1X2 U149 ( .A0N(n213), .A1N(n214), .B0(n215), .Y(n192) );
  INVX1 U150 ( .A(n221), .Y(n35) );
  NAND3X1 U151 ( .A(n232), .B(n46), .C(n233), .Y(n231) );
  NOR2BX1 U152 ( .AN(n43), .B(n234), .Y(n230) );
  NAND2X1 U153 ( .A(n49), .B(n52), .Y(n233) );
  NAND4BX2 U154 ( .AN(n24), .B(n197), .C(n198), .D(n199), .Y(n189) );
  XOR2X1 U155 ( .A(n200), .B(n201), .Y(SUM[15]) );
  XOR2X1 U156 ( .A(n203), .B(n204), .Y(SUM[14]) );
  NOR2BXL U157 ( .AN(n184), .B(n186), .Y(n204) );
  XOR2X1 U158 ( .A(n165), .B(n166), .Y(SUM[19]) );
  NAND2XL U159 ( .A(n156), .B(n161), .Y(n165) );
  NAND2X1 U160 ( .A(n30), .B(n34), .Y(n218) );
  INVX1 U161 ( .A(n38), .Y(n234) );
  XOR2X1 U162 ( .A(n136), .B(n137), .Y(SUM[22]) );
  XOR2X1 U163 ( .A(n139), .B(n140), .Y(SUM[21]) );
  NAND2XL U164 ( .A(n151), .B(n152), .Y(n146) );
  XOR2X1 U165 ( .A(n141), .B(n143), .Y(SUM[20]) );
  XOR2X1 U166 ( .A(n172), .B(n173), .Y(SUM[17]) );
  XOR2X1 U167 ( .A(n168), .B(n170), .Y(SUM[18]) );
  NAND2X1 U168 ( .A(n81), .B(n236), .Y(n238) );
  NOR2X1 U169 ( .A(n239), .B(n240), .Y(n237) );
  AOI21XL U170 ( .A0(n216), .A1(n224), .B0(n225), .Y(n223) );
  INVX1 U171 ( .A(n219), .Y(n225) );
  INVX1 U172 ( .A(n82), .Y(n163) );
  NOR2BXL U173 ( .AN(n159), .B(n157), .Y(n173) );
  OAI21XL U174 ( .A0(n163), .A1(n164), .B0(n84), .Y(n240) );
  NAND2X1 U175 ( .A(n229), .B(n34), .Y(n28) );
  NAND2X1 U176 ( .A(n32), .B(n221), .Y(n229) );
  XOR2X1 U177 ( .A(n224), .B(n226), .Y(SUM[10]) );
  NOR2BX1 U178 ( .AN(n219), .B(n227), .Y(n226) );
  INVXL U179 ( .A(n216), .Y(n227) );
  XOR2X1 U180 ( .A(n210), .B(n211), .Y(SUM[12]) );
  XOR2X1 U181 ( .A(n206), .B(n207), .Y(SUM[13]) );
  NOR2BX1 U182 ( .AN(n183), .B(n24), .Y(n207) );
  XOR2X1 U183 ( .A(n28), .B(n29), .Y(SUM[9]) );
  NAND2XL U184 ( .A(n215), .B(n220), .Y(n222) );
  XOR2X1 U185 ( .A(n32), .B(n33), .Y(SUM[8]) );
  XOR2X1 U186 ( .A(n222), .B(n223), .Y(SUM[11]) );
  NOR2BX1 U187 ( .AN(n164), .B(n27), .Y(SUM[0]) );
  OAI21XL U188 ( .A0(n25), .A1(n235), .B0(n52), .Y(n50) );
  INVX1 U189 ( .A(n50), .Y(n47) );
  XOR2X1 U190 ( .A(n50), .B(n51), .Y(SUM[5]) );
  NOR2BX1 U191 ( .AN(n49), .B(n48), .Y(n51) );
  XOR2X1 U192 ( .A(n44), .B(n45), .Y(SUM[6]) );
  NOR2BX1 U193 ( .AN(n43), .B(n42), .Y(n45) );
  INVX1 U194 ( .A(n40), .Y(n39) );
  XOR2X1 U195 ( .A(n36), .B(n37), .Y(SUM[7]) );
  OAI21XL U196 ( .A0(n41), .A1(n42), .B0(n43), .Y(n36) );
  NOR2BX1 U197 ( .AN(n38), .B(n39), .Y(n37) );
  INVX1 U198 ( .A(n44), .Y(n41) );
  INVX1 U199 ( .A(n81), .Y(n59) );
  XOR2X1 U200 ( .A(n83), .B(n162), .Y(SUM[1]) );
  XOR2X1 U201 ( .A(n61), .B(n80), .Y(SUM[2]) );
  NOR2BX1 U202 ( .AN(n60), .B(n59), .Y(n80) );
  OAI2BB1X1 U203 ( .A0N(n82), .A1N(n83), .B0(n84), .Y(n61) );
  XOR2X1 U204 ( .A(n193), .B(n53), .Y(SUM[4]) );
  NOR2BX1 U205 ( .AN(n52), .B(n25), .Y(n53) );
  XOR2X1 U206 ( .A(n54), .B(n55), .Y(SUM[3]) );
  NOR2BX1 U207 ( .AN(n56), .B(n57), .Y(n55) );
  OAI21XL U208 ( .A0(n58), .A1(n59), .B0(n60), .Y(n54) );
  NAND2X2 U209 ( .A(B[22]), .B(A[22]), .Y(n128) );
  OR2X2 U210 ( .A(A[6]), .B(B[6]), .Y(n46) );
  NAND2X1 U211 ( .A(B[21]), .B(A[21]), .Y(n127) );
  NAND2X1 U212 ( .A(B[18]), .B(A[18]), .Y(n160) );
  NAND2X2 U213 ( .A(B[11]), .B(A[11]), .Y(n220) );
  XNOR2X4 U214 ( .A(n26), .B(n73), .Y(SUM[30]) );
  NAND2X1 U215 ( .A(B[4]), .B(A[4]), .Y(n52) );
  OR2X2 U216 ( .A(A[3]), .B(B[3]), .Y(n236) );
  OR2X2 U217 ( .A(A[1]), .B(B[1]), .Y(n82) );
  NAND2X1 U218 ( .A(B[0]), .B(A[0]), .Y(n164) );
  NAND2X4 U219 ( .A(n176), .B(n177), .Y(n147) );
  NOR2BX1 U220 ( .AN(n160), .B(n149), .Y(n170) );
  INVX2 U221 ( .A(n167), .Y(n149) );
  NAND2XL U222 ( .A(B[19]), .B(A[19]), .Y(n156) );
  XOR2X1 U223 ( .A(n147), .B(n175), .Y(SUM[16]) );
  NOR2BX1 U224 ( .AN(n95), .B(n100), .Y(n106) );
  NAND3BX2 U225 ( .AN(n125), .B(n131), .C(n132), .Y(n119) );
  NOR2X4 U226 ( .A(n100), .B(n101), .Y(n92) );
  NAND2X2 U227 ( .A(A[24]), .B(B[24]), .Y(n97) );
  NOR2BXL U228 ( .AN(n181), .B(n185), .Y(n201) );
  INVX2 U229 ( .A(n124), .Y(n123) );
  NAND2X1 U230 ( .A(B[27]), .B(A[27]), .Y(n95) );
  NAND2X1 U231 ( .A(B[23]), .B(A[23]), .Y(n124) );
  NOR2BXL U232 ( .AN(n99), .B(n101), .Y(n109) );
  XOR2X1 U233 ( .A(n115), .B(n117), .Y(SUM[24]) );
  INVX8 U234 ( .A(n86), .Y(n77) );
  INVX8 U235 ( .A(n132), .Y(n129) );
  AOI21X4 U236 ( .A0(n64), .A1(n65), .B0(n66), .Y(n63) );
  OAI21X4 U237 ( .A0(n67), .A1(n68), .B0(n69), .Y(n66) );
  CLKINVX3 U238 ( .A(n72), .Y(n70) );
  OAI21X4 U239 ( .A0(n76), .A1(n77), .B0(n78), .Y(n65) );
  CLKINVX3 U240 ( .A(n79), .Y(n76) );
  OR2X4 U241 ( .A(A[29]), .B(B[29]), .Y(n72) );
  OAI21X4 U242 ( .A0(n89), .A1(n90), .B0(n91), .Y(n86) );
  AOI21X4 U243 ( .A0(n92), .A1(n93), .B0(n94), .Y(n91) );
  OAI211X2 U244 ( .A0(n96), .A1(n97), .B0(n98), .C0(n99), .Y(n93) );
  OR2X4 U245 ( .A(A[28]), .B(B[28]), .Y(n79) );
  NAND2X4 U246 ( .A(B[28]), .B(A[28]), .Y(n78) );
  XOR2X4 U247 ( .A(n105), .B(n106), .Y(SUM[27]) );
  NAND2X4 U248 ( .A(n115), .B(n116), .Y(n89) );
  OAI21X4 U249 ( .A0(n118), .A1(n119), .B0(n120), .Y(n115) );
  AOI21X4 U250 ( .A0(n121), .A1(n122), .B0(n123), .Y(n120) );
  OAI211X2 U251 ( .A0(n125), .A1(n126), .B0(n127), .C0(n128), .Y(n122) );
  NOR2X4 U252 ( .A(n129), .B(n130), .Y(n121) );
  OR2X4 U253 ( .A(A[23]), .B(B[23]), .Y(n132) );
  OR2X4 U254 ( .A(A[22]), .B(B[22]), .Y(n131) );
  OR2X4 U255 ( .A(A[21]), .B(B[21]), .Y(n138) );
  NAND2X4 U256 ( .A(n141), .B(n142), .Y(n118) );
  NAND2X4 U257 ( .A(n144), .B(n145), .Y(n141) );
  NAND3BX4 U258 ( .AN(n146), .B(n147), .C(n148), .Y(n145) );
  NOR2X4 U259 ( .A(n149), .B(n150), .Y(n148) );
  OAI211X2 U260 ( .A0(n157), .A1(n158), .B0(n159), .C0(n160), .Y(n154) );
  OR2X4 U261 ( .A(A[19]), .B(B[19]), .Y(n161) );
  OR2X4 U262 ( .A(A[18]), .B(B[18]), .Y(n167) );
  OR2X4 U263 ( .A(A[17]), .B(B[17]), .Y(n152) );
  OR2X4 U264 ( .A(A[16]), .B(B[16]), .Y(n151) );
  NAND2X4 U265 ( .A(B[16]), .B(A[16]), .Y(n158) );
  AOI21X4 U266 ( .A0(n178), .A1(n179), .B0(n180), .Y(n177) );
  OAI211X2 U267 ( .A0(n24), .A1(n182), .B0(n183), .C0(n184), .Y(n179) );
  NOR2X4 U268 ( .A(n185), .B(n186), .Y(n178) );
  OR2X4 U269 ( .A(A[15]), .B(B[15]), .Y(n199) );
  OR2X4 U270 ( .A(A[14]), .B(B[14]), .Y(n198) );
  NAND4BBX4 U271 ( .AN(n35), .BN(n31), .C(n216), .D(n215), .Y(n187) );
  OR2X4 U272 ( .A(A[11]), .B(B[11]), .Y(n215) );
  OR2X4 U273 ( .A(A[10]), .B(B[10]), .Y(n216) );
endmodule


module hash_core_DW01_add_26 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n215, n216, n217, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214;

  NAND4BX1 U2 ( .AN(n104), .B(n105), .C(n106), .D(n107), .Y(n103) );
  AOI21X2 U3 ( .A0(n173), .A1(n174), .B0(n167), .Y(n171) );
  XOR2X2 U4 ( .A(n32), .B(n33), .Y(SUM[7]) );
  OAI21X4 U5 ( .A0(n155), .A1(n156), .B0(n157), .Y(n151) );
  NOR2X2 U6 ( .A(n171), .B(n172), .Y(n155) );
  NAND4BX1 U7 ( .AN(n17), .B(n198), .C(n193), .D(n194), .Y(n167) );
  OAI21X2 U8 ( .A0(n17), .A1(n188), .B0(n31), .Y(n25) );
  NOR2X1 U9 ( .A(A[8]), .B(B[8]), .Y(n17) );
  NAND2X2 U10 ( .A(n121), .B(n116), .Y(n119) );
  OAI21X1 U11 ( .A0(n64), .A1(n65), .B0(n66), .Y(n62) );
  BUFX3 U12 ( .A(n215), .Y(SUM[30]) );
  BUFX4 U13 ( .A(n217), .Y(SUM[25]) );
  OAI21X4 U14 ( .A0(n19), .A1(n185), .B0(n165), .Y(n183) );
  INVX4 U15 ( .A(n186), .Y(n185) );
  BUFX3 U16 ( .A(n216), .Y(SUM[29]) );
  XOR2X4 U17 ( .A(n95), .B(n15), .Y(SUM[26]) );
  BUFX3 U18 ( .A(n62), .Y(n4) );
  XOR2X4 U19 ( .A(n93), .B(n94), .Y(SUM[27]) );
  NAND3BXL U20 ( .AN(n20), .B(n140), .C(n141), .Y(n129) );
  OAI21X1 U21 ( .A0(n159), .A1(n18), .B0(n160), .Y(n158) );
  CLKINVX3 U22 ( .A(n29), .Y(n188) );
  NAND2X1 U23 ( .A(n6), .B(n130), .Y(n124) );
  NOR2BX1 U24 ( .AN(n139), .B(n131), .Y(n130) );
  NAND2X1 U25 ( .A(n124), .B(n125), .Y(n104) );
  NAND2X1 U26 ( .A(n100), .B(n101), .Y(n80) );
  INVX1 U27 ( .A(n198), .Y(n28) );
  CLKINVX3 U28 ( .A(n5), .Y(n7) );
  NAND2X1 U29 ( .A(n97), .B(n92), .Y(n95) );
  NAND2X1 U30 ( .A(n81), .B(n98), .Y(n97) );
  XOR2X2 U31 ( .A(n178), .B(n179), .Y(SUM[15]) );
  OAI2BB1X2 U32 ( .A0N(n161), .A1N(n180), .B0(n164), .Y(n178) );
  INVX1 U33 ( .A(n209), .Y(n37) );
  AND2X2 U34 ( .A(B[4]), .B(A[4]), .Y(n5) );
  NAND2X1 U35 ( .A(B[2]), .B(A[2]), .Y(n58) );
  XOR2X2 U36 ( .A(n143), .B(n144), .Y(SUM[19]) );
  XOR2X4 U37 ( .A(n199), .B(n200), .Y(SUM[11]) );
  INVX2 U38 ( .A(n183), .Y(n182) );
  INVX2 U39 ( .A(n25), .Y(n205) );
  XOR2X2 U40 ( .A(n201), .B(n203), .Y(SUM[10]) );
  AOI21X2 U41 ( .A0(n74), .A1(n75), .B0(n76), .Y(n65) );
  AOI21X1 U42 ( .A0(n194), .A1(n201), .B0(n202), .Y(n200) );
  OR2XL U43 ( .A(n128), .B(n129), .Y(n6) );
  NAND2X4 U44 ( .A(n151), .B(n152), .Y(n128) );
  OAI21X4 U45 ( .A0(n182), .A1(n16), .B0(n166), .Y(n180) );
  XOR2X2 U46 ( .A(n180), .B(n181), .Y(SUM[14]) );
  NAND3BX4 U47 ( .AN(n177), .B(n54), .C(n176), .Y(n46) );
  NAND3X2 U48 ( .A(n211), .B(n70), .C(n212), .Y(n176) );
  NOR2XL U49 ( .A(n16), .B(n19), .Y(n168) );
  NAND2XL U50 ( .A(n104), .B(n115), .Y(n122) );
  OAI21X2 U51 ( .A0(n16), .A1(n165), .B0(n166), .Y(n162) );
  XNOR2X1 U52 ( .A(n119), .B(n13), .Y(SUM[22]) );
  XNOR2X1 U53 ( .A(n4), .B(n10), .Y(n215) );
  OR2X1 U54 ( .A(A[1]), .B(B[1]), .Y(n70) );
  OAI21XL U55 ( .A0(n36), .A1(n37), .B0(n38), .Y(n32) );
  OAI21XL U56 ( .A0(n56), .A1(n57), .B0(n58), .Y(n52) );
  NOR2BXL U57 ( .AN(n54), .B(n55), .Y(n53) );
  NOR2BX1 U58 ( .AN(n7), .B(n51), .Y(n50) );
  NOR2BXL U59 ( .AN(n54), .B(n177), .Y(n175) );
  NAND3XL U60 ( .A(n44), .B(n209), .C(n210), .Y(n207) );
  INVX1 U61 ( .A(n88), .Y(n96) );
  AOI21X1 U62 ( .A0(n83), .A1(n95), .B0(n96), .Y(n94) );
  INVX1 U63 ( .A(n164), .Y(n163) );
  NAND2X1 U64 ( .A(B[5]), .B(A[5]), .Y(n42) );
  NAND2X1 U65 ( .A(B[6]), .B(A[6]), .Y(n38) );
  NAND2X1 U66 ( .A(B[1]), .B(A[1]), .Y(n71) );
  OR2X2 U67 ( .A(A[5]), .B(B[5]), .Y(n44) );
  OR2X2 U68 ( .A(A[17]), .B(B[17]), .Y(n141) );
  OAI21X1 U69 ( .A0(n188), .A1(n167), .B0(n189), .Y(n186) );
  AND2X2 U70 ( .A(n8), .B(n9), .Y(n14) );
  NOR2X1 U71 ( .A(n47), .B(n51), .Y(n8) );
  NOR2X1 U72 ( .A(n35), .B(n37), .Y(n9) );
  NAND2XL U73 ( .A(n58), .B(n72), .Y(n68) );
  OAI21X1 U74 ( .A0(n205), .A1(n28), .B0(n27), .Y(n201) );
  OAI21X2 U75 ( .A0(n190), .A1(n191), .B0(n192), .Y(n172) );
  NAND2XL U76 ( .A(n193), .B(n194), .Y(n191) );
  NOR2BXL U77 ( .AN(n164), .B(n170), .Y(n181) );
  INVXL U78 ( .A(n194), .Y(n204) );
  NAND2X1 U79 ( .A(n60), .B(n63), .Y(n10) );
  NAND2XL U80 ( .A(n192), .B(n193), .Y(n199) );
  INVXL U81 ( .A(n197), .Y(n202) );
  NOR2BXL U82 ( .AN(n34), .B(n35), .Y(n33) );
  NOR2XL U83 ( .A(n7), .B(n47), .Y(n41) );
  NAND3XL U84 ( .A(n44), .B(n45), .C(n46), .Y(n43) );
  AND2X2 U85 ( .A(n38), .B(n34), .Y(n206) );
  XNOR2X1 U86 ( .A(n100), .B(n11), .Y(SUM[24]) );
  NAND2X1 U87 ( .A(n91), .B(n101), .Y(n11) );
  XNOR2X1 U88 ( .A(n74), .B(n12), .Y(SUM[28]) );
  NAND2X1 U89 ( .A(n77), .B(n75), .Y(n12) );
  NOR2BXL U90 ( .AN(n27), .B(n28), .Y(n26) );
  NOR2BXL U91 ( .AN(n38), .B(n37), .Y(n40) );
  NOR2BXL U92 ( .AN(n133), .B(n134), .Y(n147) );
  XOR2XL U93 ( .A(n73), .B(n65), .Y(n216) );
  NOR2BXL U94 ( .AN(n139), .B(n20), .Y(n144) );
  NAND2X1 U95 ( .A(n112), .B(n107), .Y(n13) );
  NAND2XL U96 ( .A(n128), .B(n137), .Y(n149) );
  NAND2XL U97 ( .A(n4), .B(n63), .Y(n61) );
  NAND2XL U98 ( .A(B[9]), .B(A[9]), .Y(n27) );
  NOR2XL U99 ( .A(A[12]), .B(B[12]), .Y(n19) );
  NAND2XL U100 ( .A(B[13]), .B(A[13]), .Y(n166) );
  NAND2XL U101 ( .A(B[11]), .B(A[11]), .Y(n192) );
  NAND2XL U102 ( .A(B[7]), .B(A[7]), .Y(n34) );
  NAND2XL U103 ( .A(B[18]), .B(A[18]), .Y(n133) );
  NAND2XL U104 ( .A(B[19]), .B(A[19]), .Y(n139) );
  NAND2XL U105 ( .A(B[15]), .B(A[15]), .Y(n160) );
  OR2XL U106 ( .A(A[16]), .B(B[16]), .Y(n152) );
  INVX1 U107 ( .A(n172), .Y(n189) );
  OAI2BB1X1 U108 ( .A0N(n14), .A1N(n46), .B0(n174), .Y(n29) );
  NAND2X1 U109 ( .A(n168), .B(n169), .Y(n156) );
  INVX1 U110 ( .A(n158), .Y(n157) );
  NOR2BX1 U111 ( .AN(n160), .B(n18), .Y(n179) );
  INVX1 U112 ( .A(n72), .Y(n57) );
  INVX1 U113 ( .A(n213), .Y(n55) );
  NOR2BX1 U114 ( .AN(n197), .B(n204), .Y(n203) );
  NOR2X1 U115 ( .A(n195), .B(n196), .Y(n190) );
  NAND2X1 U116 ( .A(n27), .B(n197), .Y(n196) );
  NAND3BX1 U117 ( .AN(n41), .B(n42), .C(n43), .Y(n39) );
  INVX1 U118 ( .A(n44), .Y(n47) );
  INVX1 U119 ( .A(n45), .Y(n51) );
  INVX1 U120 ( .A(n208), .Y(n35) );
  XOR2X1 U121 ( .A(n46), .B(n50), .Y(SUM[4]) );
  XOR2X1 U122 ( .A(n183), .B(n184), .Y(SUM[13]) );
  NOR2BX1 U123 ( .AN(n166), .B(n16), .Y(n184) );
  XOR2X1 U124 ( .A(n25), .B(n26), .Y(SUM[9]) );
  XOR2X1 U125 ( .A(n186), .B(n187), .Y(SUM[12]) );
  NOR2BX1 U126 ( .AN(n165), .B(n19), .Y(n187) );
  XOR2X1 U127 ( .A(n39), .B(n40), .Y(SUM[6]) );
  INVX1 U128 ( .A(n39), .Y(n36) );
  OAI21XL U129 ( .A0(n145), .A1(n134), .B0(n133), .Y(n143) );
  INVX1 U130 ( .A(n146), .Y(n145) );
  XOR2X1 U131 ( .A(n52), .B(n53), .Y(SUM[3]) );
  XOR2X1 U132 ( .A(n68), .B(n56), .Y(SUM[2]) );
  XOR2X1 U133 ( .A(n48), .B(n49), .Y(SUM[5]) );
  NAND2X1 U134 ( .A(n44), .B(n42), .Y(n48) );
  AOI21X1 U135 ( .A0(n46), .A1(n45), .B0(n5), .Y(n49) );
  XOR2X1 U136 ( .A(n29), .B(n30), .Y(SUM[8]) );
  NOR2BX1 U137 ( .AN(n31), .B(n17), .Y(n30) );
  OAI2BB1X1 U138 ( .A0N(n175), .A1N(n176), .B0(n14), .Y(n173) );
  AOI21X1 U139 ( .A0(n161), .A1(n162), .B0(n163), .Y(n159) );
  NAND2X1 U140 ( .A(n105), .B(n122), .Y(n121) );
  OAI2BB1X1 U141 ( .A0N(n206), .A1N(n207), .B0(n208), .Y(n174) );
  NOR2X1 U142 ( .A(n28), .B(n31), .Y(n195) );
  NAND2X1 U143 ( .A(n148), .B(n138), .Y(n146) );
  NAND2X1 U144 ( .A(n141), .B(n149), .Y(n148) );
  INVX1 U145 ( .A(n214), .Y(n177) );
  NAND2BX1 U146 ( .AN(n58), .B(n213), .Y(n214) );
  NAND2X1 U147 ( .A(n7), .B(n42), .Y(n210) );
  NAND2X1 U148 ( .A(n71), .B(n70), .Y(n142) );
  INVX1 U149 ( .A(n77), .Y(n76) );
  NAND2X1 U150 ( .A(n86), .B(n82), .Y(n93) );
  INVX1 U151 ( .A(n67), .Y(n64) );
  INVX1 U152 ( .A(n140), .Y(n134) );
  XOR2X1 U153 ( .A(n124), .B(n126), .Y(SUM[20]) );
  NOR2BX1 U154 ( .AN(n115), .B(n127), .Y(n126) );
  INVX1 U155 ( .A(n125), .Y(n127) );
  AND2X2 U156 ( .A(n88), .B(n83), .Y(n15) );
  XOR2X1 U157 ( .A(n117), .B(n118), .Y(SUM[23]) );
  NAND2X1 U158 ( .A(n110), .B(n106), .Y(n117) );
  AOI21X1 U159 ( .A0(n107), .A1(n119), .B0(n120), .Y(n118) );
  INVX1 U160 ( .A(n112), .Y(n120) );
  XOR2X1 U161 ( .A(n122), .B(n123), .Y(SUM[21]) );
  NOR2BX1 U162 ( .AN(n116), .B(n114), .Y(n123) );
  INVX1 U163 ( .A(n141), .Y(n136) );
  INVX1 U164 ( .A(n161), .Y(n170) );
  AOI21X1 U165 ( .A0(n132), .A1(n133), .B0(n20), .Y(n131) );
  NAND2BX1 U166 ( .AN(n134), .B(n135), .Y(n132) );
  OAI21XL U167 ( .A0(n136), .A1(n137), .B0(n138), .Y(n135) );
  NAND2X1 U168 ( .A(n102), .B(n103), .Y(n100) );
  AOI21X1 U169 ( .A0(n108), .A1(n106), .B0(n109), .Y(n102) );
  INVX1 U170 ( .A(n110), .Y(n109) );
  XOR2X1 U171 ( .A(n149), .B(n150), .Y(SUM[17]) );
  NOR2BX1 U172 ( .AN(n138), .B(n136), .Y(n150) );
  NAND2X1 U173 ( .A(n66), .B(n67), .Y(n73) );
  XOR2X1 U174 ( .A(n146), .B(n147), .Y(SUM[18]) );
  NAND2X1 U175 ( .A(n80), .B(n91), .Y(n98) );
  NAND2X1 U176 ( .A(n78), .B(n79), .Y(n74) );
  AOI21X1 U177 ( .A0(n84), .A1(n82), .B0(n85), .Y(n78) );
  NAND4BXL U178 ( .AN(n80), .B(n81), .C(n82), .D(n83), .Y(n79) );
  INVX1 U179 ( .A(n86), .Y(n85) );
  XOR2X1 U180 ( .A(n151), .B(n153), .Y(SUM[16]) );
  NOR2BX1 U181 ( .AN(n137), .B(n154), .Y(n153) );
  INVX1 U182 ( .A(n152), .Y(n154) );
  XOR2X1 U183 ( .A(n98), .B(n99), .Y(n217) );
  NOR2BX1 U184 ( .AN(n92), .B(n90), .Y(n99) );
  NOR2X1 U185 ( .A(n18), .B(n170), .Y(n169) );
  INVX1 U186 ( .A(n105), .Y(n114) );
  NAND2X1 U187 ( .A(n111), .B(n112), .Y(n108) );
  NAND2X1 U188 ( .A(n107), .B(n113), .Y(n111) );
  OAI21XL U189 ( .A0(n114), .A1(n115), .B0(n116), .Y(n113) );
  NAND2X1 U190 ( .A(n60), .B(n61), .Y(n59) );
  INVX1 U191 ( .A(n81), .Y(n90) );
  NAND2X1 U192 ( .A(n87), .B(n88), .Y(n84) );
  NAND2X1 U193 ( .A(n83), .B(n89), .Y(n87) );
  OAI21XL U194 ( .A0(n90), .A1(n91), .B0(n92), .Y(n89) );
  XOR3X2 U195 ( .A(B[31]), .B(A[31]), .C(n59), .Y(SUM[31]) );
  OAI2BB1X1 U196 ( .A0N(B[0]), .A1N(A[0]), .B0(n71), .Y(n212) );
  NOR2X1 U197 ( .A(n55), .B(n57), .Y(n211) );
  OR2X2 U198 ( .A(A[3]), .B(B[3]), .Y(n213) );
  OR2X2 U199 ( .A(A[2]), .B(B[2]), .Y(n72) );
  NOR2X1 U200 ( .A(A[13]), .B(B[13]), .Y(n16) );
  AND2X2 U201 ( .A(n71), .B(n69), .Y(n56) );
  NAND3X1 U202 ( .A(A[0]), .B(B[0]), .C(n70), .Y(n69) );
  OR2X2 U203 ( .A(A[10]), .B(B[10]), .Y(n194) );
  NAND2X1 U204 ( .A(B[8]), .B(A[8]), .Y(n31) );
  OR2X2 U205 ( .A(A[11]), .B(B[11]), .Y(n193) );
  NAND2X1 U206 ( .A(B[10]), .B(A[10]), .Y(n197) );
  NAND2X1 U207 ( .A(B[3]), .B(A[3]), .Y(n54) );
  OR2X2 U208 ( .A(A[4]), .B(B[4]), .Y(n45) );
  XOR2X1 U209 ( .A(n24), .B(n142), .Y(SUM[1]) );
  NAND2X1 U210 ( .A(B[0]), .B(A[0]), .Y(n24) );
  OR2X2 U211 ( .A(A[9]), .B(B[9]), .Y(n198) );
  OR2X2 U212 ( .A(A[6]), .B(B[6]), .Y(n209) );
  OR2X2 U213 ( .A(A[7]), .B(B[7]), .Y(n208) );
  NOR2X1 U214 ( .A(A[15]), .B(B[15]), .Y(n18) );
  NOR2X1 U215 ( .A(A[19]), .B(B[19]), .Y(n20) );
  NAND2X1 U216 ( .A(B[16]), .B(A[16]), .Y(n137) );
  NAND2X1 U217 ( .A(B[12]), .B(A[12]), .Y(n165) );
  NAND2X1 U218 ( .A(B[17]), .B(A[17]), .Y(n138) );
  NAND2X1 U219 ( .A(B[14]), .B(A[14]), .Y(n164) );
  NOR2X1 U220 ( .A(n22), .B(n23), .Y(SUM[0]) );
  NOR2X1 U221 ( .A(A[0]), .B(B[0]), .Y(n22) );
  AND2X2 U222 ( .A(B[0]), .B(A[0]), .Y(n23) );
  OR2X2 U223 ( .A(A[14]), .B(B[14]), .Y(n161) );
  OR2X2 U224 ( .A(A[18]), .B(B[18]), .Y(n140) );
  OR2X2 U225 ( .A(A[22]), .B(B[22]), .Y(n107) );
  NAND2X1 U226 ( .A(B[22]), .B(A[22]), .Y(n112) );
  NAND2X1 U227 ( .A(B[20]), .B(A[20]), .Y(n115) );
  OR2X2 U228 ( .A(A[23]), .B(B[23]), .Y(n106) );
  NAND2X1 U229 ( .A(B[21]), .B(A[21]), .Y(n116) );
  OR2X2 U230 ( .A(A[21]), .B(B[21]), .Y(n105) );
  OR2X2 U231 ( .A(A[20]), .B(B[20]), .Y(n125) );
  OR2X2 U232 ( .A(A[26]), .B(B[26]), .Y(n83) );
  NAND2X1 U233 ( .A(B[24]), .B(A[24]), .Y(n91) );
  NAND2X1 U234 ( .A(B[26]), .B(A[26]), .Y(n88) );
  OR2X2 U235 ( .A(A[27]), .B(B[27]), .Y(n82) );
  NAND2X1 U236 ( .A(B[25]), .B(A[25]), .Y(n92) );
  OR2X2 U237 ( .A(A[25]), .B(B[25]), .Y(n81) );
  NAND2X1 U238 ( .A(B[23]), .B(A[23]), .Y(n110) );
  NAND2X1 U239 ( .A(B[27]), .B(A[27]), .Y(n86) );
  OR2X2 U240 ( .A(A[24]), .B(B[24]), .Y(n101) );
  NAND2X1 U241 ( .A(B[30]), .B(A[30]), .Y(n60) );
  NAND2X1 U242 ( .A(B[29]), .B(A[29]), .Y(n66) );
  NAND2X1 U243 ( .A(B[28]), .B(A[28]), .Y(n77) );
  OR2X2 U244 ( .A(A[28]), .B(B[28]), .Y(n75) );
  OR2X2 U245 ( .A(A[30]), .B(B[30]), .Y(n63) );
  OR2X2 U246 ( .A(A[29]), .B(B[29]), .Y(n67) );
endmodule


module hash_core_DW01_add_24 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n340, n341, n342, n343, n344, n345, n346, n1, n2, n3, n4, n5, n6, n8,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339;

  NAND2X2 U2 ( .A(n236), .B(n268), .Y(n64) );
  NAND3X1 U3 ( .A(n294), .B(n295), .C(n296), .Y(n282) );
  CLKINVX2 U4 ( .A(n285), .Y(n284) );
  NAND2X2 U5 ( .A(B[19]), .B(n16), .Y(n214) );
  INVX8 U6 ( .A(n216), .Y(n225) );
  NAND2X2 U7 ( .A(n178), .B(n191), .Y(n188) );
  NAND2X4 U8 ( .A(B[10]), .B(A[10]), .Y(n316) );
  NAND2BX4 U9 ( .AN(n106), .B(n94), .Y(n98) );
  OAI21X2 U10 ( .A0(n257), .A1(n258), .B0(n259), .Y(n256) );
  INVX4 U11 ( .A(n251), .Y(n260) );
  BUFX20 U12 ( .A(n341), .Y(SUM[21]) );
  NOR2X2 U13 ( .A(n225), .B(n226), .Y(n230) );
  INVX2 U14 ( .A(n179), .Y(n184) );
  NOR2X2 U15 ( .A(n232), .B(n233), .Y(n254) );
  OR2X1 U16 ( .A(A[9]), .B(B[9]), .Y(n1) );
  NAND2XL U17 ( .A(n1), .B(n295), .Y(n334) );
  OR2X4 U18 ( .A(n250), .B(n273), .Y(n2) );
  NAND2X4 U19 ( .A(n2), .B(n274), .Y(n231) );
  AND3X2 U20 ( .A(n263), .B(n270), .C(n269), .Y(n250) );
  XNOR2X2 U21 ( .A(n231), .B(n272), .Y(n13) );
  NAND2X2 U22 ( .A(n253), .B(n4), .Y(n5) );
  NAND2X4 U23 ( .A(n3), .B(n42), .Y(n6) );
  NAND2X4 U24 ( .A(n5), .B(n6), .Y(SUM[18]) );
  INVX4 U25 ( .A(n253), .Y(n3) );
  INVX2 U26 ( .A(n42), .Y(n4) );
  OAI2BB1X4 U27 ( .A0N(n254), .A1N(n255), .B0(n218), .Y(n253) );
  AND2X4 U28 ( .A(n215), .B(n244), .Y(n42) );
  OAI21X2 U29 ( .A0(A[11]), .A1(B[11]), .B0(n296), .Y(n320) );
  NAND2X1 U30 ( .A(B[18]), .B(A[18]), .Y(n244) );
  BUFX12 U31 ( .A(n342), .Y(SUM[14]) );
  NAND2X4 U32 ( .A(n136), .B(n240), .Y(n339) );
  NAND2X2 U33 ( .A(B[1]), .B(A[1]), .Y(n136) );
  INVX8 U34 ( .A(n295), .Y(n76) );
  AND3X2 U35 ( .A(n315), .B(n319), .C(n306), .Y(n51) );
  NAND2BX2 U36 ( .AN(n60), .B(n293), .Y(n319) );
  CLKINVX4 U37 ( .A(n108), .Y(n33) );
  AOI21X4 U38 ( .A0(n45), .A1(n95), .B0(n110), .Y(n108) );
  BUFX4 U39 ( .A(n325), .Y(n8) );
  NAND2X2 U40 ( .A(n218), .B(n236), .Y(n247) );
  NOR2X4 U41 ( .A(n260), .B(n261), .Y(n259) );
  AOI21X4 U42 ( .A0(n286), .A1(n287), .B0(n288), .Y(n283) );
  INVX2 U43 ( .A(n289), .Y(n288) );
  CLKINVX3 U44 ( .A(n291), .Y(n286) );
  NAND3BX2 U45 ( .AN(n250), .B(n251), .C(n252), .Y(n248) );
  AOI21X1 U46 ( .A0(B[11]), .A1(A[11]), .B0(n297), .Y(n325) );
  NOR2BX4 U47 ( .AN(n316), .B(n327), .Y(n329) );
  CLKINVX2 U48 ( .A(n296), .Y(n327) );
  INVX4 U49 ( .A(n290), .Y(n100) );
  NAND2BX4 U50 ( .AN(n117), .B(n114), .Y(n290) );
  OAI21X1 U51 ( .A0(A[13]), .A1(B[13]), .B0(n308), .Y(n307) );
  NOR2BX1 U52 ( .AN(n71), .B(n76), .Y(n82) );
  OAI2BB1X4 U53 ( .A0N(B[9]), .A1N(A[9]), .B0(n71), .Y(n323) );
  BUFX12 U54 ( .A(n340), .Y(SUM[27]) );
  NOR2XL U55 ( .A(A[3]), .B(B[3]), .Y(n338) );
  OR2X4 U56 ( .A(A[3]), .B(B[3]), .Y(n114) );
  BUFX12 U57 ( .A(n345), .Y(SUM[5]) );
  AND2X2 U58 ( .A(n216), .B(n214), .Y(n43) );
  INVX4 U59 ( .A(n118), .Y(n115) );
  CLKINVX3 U60 ( .A(n118), .Y(n47) );
  NAND2X2 U61 ( .A(n118), .B(n48), .Y(n49) );
  OAI2BB1X2 U62 ( .A0N(n134), .A1N(n135), .B0(n136), .Y(n118) );
  NAND2X4 U63 ( .A(B[21]), .B(A[21]), .Y(n175) );
  OR2X4 U64 ( .A(A[20]), .B(B[20]), .Y(n190) );
  NAND2X4 U65 ( .A(B[20]), .B(A[20]), .Y(n194) );
  NOR3X4 U66 ( .A(n195), .B(n202), .C(n203), .Y(n201) );
  INVX4 U67 ( .A(n178), .Y(n195) );
  AND2X1 U68 ( .A(n194), .B(n214), .Y(n213) );
  INVX4 U69 ( .A(n194), .Y(n200) );
  NAND2BX4 U70 ( .AN(n194), .B(n191), .Y(n174) );
  NOR2BX4 U71 ( .AN(n194), .B(n202), .Y(n227) );
  AOI21X4 U72 ( .A0(n222), .A1(n190), .B0(n200), .Y(n221) );
  NOR2X4 U73 ( .A(n203), .B(n202), .Y(n206) );
  CLKINVX4 U74 ( .A(n191), .Y(n203) );
  OAI21X1 U75 ( .A0(n149), .A1(n155), .B0(n156), .Y(n152) );
  INVX4 U76 ( .A(n162), .Y(n149) );
  OR2X4 U77 ( .A(A[1]), .B(B[1]), .Y(n134) );
  NAND2X4 U78 ( .A(B[2]), .B(A[2]), .Y(n117) );
  OR2X4 U79 ( .A(A[2]), .B(B[2]), .Y(n133) );
  NAND2X2 U80 ( .A(n124), .B(n122), .Y(n37) );
  CLKINVX3 U81 ( .A(n121), .Y(n36) );
  NOR2BX2 U82 ( .AN(n143), .B(n61), .Y(n158) );
  NAND2X2 U83 ( .A(n162), .B(n154), .Y(n160) );
  NOR2BX2 U84 ( .AN(n155), .B(n150), .Y(n185) );
  NAND3X2 U85 ( .A(n15), .B(n173), .C(n39), .Y(n182) );
  NAND3X2 U86 ( .A(n174), .B(n175), .C(n193), .Y(n183) );
  INVX1 U87 ( .A(n128), .Y(n131) );
  NAND2X1 U88 ( .A(B[13]), .B(A[13]), .Y(n263) );
  OAI21X2 U89 ( .A0(n151), .A1(n152), .B0(n153), .Y(n142) );
  INVX1 U90 ( .A(n161), .Y(n151) );
  NAND3X2 U91 ( .A(n145), .B(n146), .C(n147), .Y(n141) );
  NOR2X1 U92 ( .A(n297), .B(n280), .Y(n314) );
  OAI21X2 U93 ( .A0(n69), .A1(n71), .B0(n68), .Y(n335) );
  NAND2X2 U94 ( .A(n99), .B(n106), .Y(n333) );
  INVX2 U95 ( .A(n190), .Y(n202) );
  NOR2X2 U96 ( .A(n232), .B(n233), .Y(n229) );
  NAND2X2 U97 ( .A(B[16]), .B(A[16]), .Y(n236) );
  NAND2X2 U98 ( .A(B[24]), .B(A[24]), .Y(n155) );
  OR2X2 U99 ( .A(A[25]), .B(B[25]), .Y(n162) );
  NOR2X1 U100 ( .A(n149), .B(n150), .Y(n167) );
  OAI21X1 U101 ( .A0(n262), .A1(n305), .B0(n304), .Y(n303) );
  INVX1 U102 ( .A(n309), .Y(n22) );
  INVX1 U103 ( .A(n80), .Y(n337) );
  AOI21X2 U104 ( .A0(n95), .A1(n109), .B0(n97), .Y(n92) );
  NAND2X2 U105 ( .A(B[4]), .B(A[4]), .Y(n106) );
  INVX1 U106 ( .A(n240), .Y(n135) );
  BUFX12 U107 ( .A(n343), .Y(SUM[12]) );
  NAND2X1 U108 ( .A(n262), .B(n308), .Y(n318) );
  BUFX8 U109 ( .A(n344), .Y(SUM[9]) );
  XOR2X2 U110 ( .A(n119), .B(n120), .Y(SUM[31]) );
  AND2X2 U111 ( .A(n311), .B(n308), .Y(n31) );
  INVX1 U112 ( .A(n306), .Y(n311) );
  AOI31X1 U113 ( .A0(n269), .A1(n263), .A2(n270), .B0(n271), .Y(n267) );
  NAND2X2 U114 ( .A(n252), .B(n251), .Y(n271) );
  NOR2X4 U115 ( .A(n280), .B(n281), .Y(n279) );
  AND2X2 U116 ( .A(n89), .B(n80), .Y(n12) );
  INVX8 U117 ( .A(n62), .Y(n94) );
  NAND4BXL U118 ( .AN(n62), .B(n95), .C(n80), .D(n79), .Y(n291) );
  AND2X4 U119 ( .A(n17), .B(n229), .Y(n14) );
  OAI2BB1X2 U120 ( .A0N(n230), .A1N(n224), .B0(n214), .Y(n223) );
  NAND4BBX4 U121 ( .AN(n187), .BN(n188), .C(n189), .D(n190), .Y(n15) );
  NAND4BBX2 U122 ( .AN(n187), .BN(n188), .C(n189), .D(n190), .Y(n171) );
  NOR2X1 U123 ( .A(A[23]), .B(B[23]), .Y(n187) );
  NOR2X1 U124 ( .A(n130), .B(n131), .Y(n125) );
  AND2X2 U125 ( .A(n270), .B(n252), .Y(n41) );
  NAND3BX2 U126 ( .AN(n64), .B(n256), .C(n249), .Y(n255) );
  NAND3BX4 U127 ( .AN(n267), .B(n18), .C(n268), .Y(n265) );
  AND2X2 U128 ( .A(n317), .B(n316), .Y(n60) );
  BUFX3 U129 ( .A(A[19]), .Y(n16) );
  NAND2X4 U130 ( .A(n84), .B(n289), .Y(n321) );
  OAI21X4 U131 ( .A0(n282), .A1(n283), .B0(n284), .Y(n278) );
  AOI2BB1X4 U132 ( .A0N(n84), .A1N(n334), .B0(n335), .Y(n330) );
  NOR2X4 U133 ( .A(n225), .B(n226), .Y(n17) );
  INVX4 U134 ( .A(n215), .Y(n226) );
  NAND3BX4 U135 ( .AN(n277), .B(n278), .C(n279), .Y(n18) );
  CLKINVX3 U136 ( .A(n171), .Y(n19) );
  INVX4 U137 ( .A(n19), .Y(n20) );
  NOR2BX2 U138 ( .AN(n268), .B(n260), .Y(n299) );
  NAND3BX2 U139 ( .AN(n170), .B(n15), .C(n172), .Y(n168) );
  OAI21X4 U140 ( .A0(n115), .A1(n116), .B0(n117), .Y(n112) );
  CLKINVX3 U141 ( .A(n133), .Y(n116) );
  NOR2X1 U142 ( .A(n149), .B(n150), .Y(n145) );
  NAND2X1 U143 ( .A(n183), .B(n178), .Y(n39) );
  NAND2X1 U144 ( .A(n191), .B(n175), .Y(n220) );
  NAND2X2 U145 ( .A(n57), .B(n141), .Y(n139) );
  NAND3X1 U146 ( .A(n94), .B(n95), .C(n96), .Y(n105) );
  AOI21X4 U147 ( .A0(n245), .A1(n246), .B0(n247), .Y(n242) );
  INVX2 U148 ( .A(n252), .Y(n261) );
  NOR2X2 U149 ( .A(n61), .B(n148), .Y(n153) );
  NOR2X2 U150 ( .A(n148), .B(n61), .Y(n147) );
  NOR2X2 U151 ( .A(n75), .B(n76), .Y(n73) );
  NAND3X4 U152 ( .A(n292), .B(n252), .C(n293), .Y(n277) );
  NAND3X2 U153 ( .A(n268), .B(n248), .C(n249), .Y(n246) );
  BUFX4 U154 ( .A(n91), .Y(n21) );
  AOI21X4 U155 ( .A0(n139), .A1(n127), .B0(n140), .Y(n138) );
  NAND2X1 U156 ( .A(B[25]), .B(A[25]), .Y(n156) );
  NOR2BX4 U157 ( .AN(n106), .B(n78), .Y(n111) );
  NAND3X4 U158 ( .A(n129), .B(n128), .C(n127), .Y(n40) );
  NAND2X2 U159 ( .A(B[26]), .B(A[26]), .Y(n161) );
  NAND2X2 U160 ( .A(n73), .B(n74), .Y(n72) );
  NAND2X1 U161 ( .A(n154), .B(n161), .Y(n165) );
  NAND4BX2 U162 ( .AN(n332), .B(n295), .C(n79), .D(n74), .Y(n331) );
  NOR2X1 U163 ( .A(A[9]), .B(B[9]), .Y(n332) );
  NAND2X4 U164 ( .A(n309), .B(n23), .Y(n24) );
  NAND2X2 U165 ( .A(n22), .B(n310), .Y(n25) );
  NAND2X4 U166 ( .A(n24), .B(n25), .Y(SUM[13]) );
  INVX4 U167 ( .A(n310), .Y(n23) );
  NAND2X4 U168 ( .A(n316), .B(n315), .Y(n26) );
  NAND2X4 U169 ( .A(n27), .B(n317), .Y(n285) );
  INVX4 U170 ( .A(n26), .Y(n27) );
  NAND2X4 U171 ( .A(B[11]), .B(A[11]), .Y(n315) );
  NAND2X2 U172 ( .A(n314), .B(n285), .Y(n313) );
  NAND2X4 U173 ( .A(n14), .B(n231), .Y(n210) );
  NAND2BX2 U174 ( .AN(n209), .B(n210), .Y(n207) );
  NAND3X1 U175 ( .A(n53), .B(n109), .C(n77), .Y(n70) );
  INVX8 U176 ( .A(n13), .Y(SUM[16]) );
  NAND2X4 U177 ( .A(B[14]), .B(A[14]), .Y(n270) );
  NAND3X2 U178 ( .A(n142), .B(n143), .C(n141), .Y(n129) );
  INVX3 U179 ( .A(n18), .Y(n276) );
  BUFX3 U180 ( .A(n346), .Y(SUM[0]) );
  NAND2BX4 U181 ( .AN(n198), .B(n199), .Y(n196) );
  OAI21X2 U182 ( .A0(n200), .A1(n189), .B0(n201), .Y(n199) );
  NOR2X2 U183 ( .A(A[13]), .B(B[13]), .Y(n305) );
  NAND2X2 U184 ( .A(B[13]), .B(A[13]), .Y(n304) );
  XOR2X4 U185 ( .A(n81), .B(n82), .Y(SUM[8]) );
  NOR2X2 U186 ( .A(n306), .B(n307), .Y(n301) );
  AOI21X2 U187 ( .A0(n121), .A1(n122), .B0(n123), .Y(n120) );
  NAND2X2 U188 ( .A(n32), .B(n108), .Y(n35) );
  NAND2BX2 U189 ( .AN(n223), .B(n210), .Y(n222) );
  NOR2X2 U190 ( .A(n184), .B(n195), .Y(n192) );
  OAI21X1 U191 ( .A0(n195), .A1(n175), .B0(n204), .Y(n198) );
  AOI21X4 U192 ( .A0(n167), .A1(n168), .B0(n169), .Y(n166) );
  NOR3X2 U193 ( .A(n76), .B(n62), .C(n78), .Y(n77) );
  NAND2BX4 U194 ( .AN(n262), .B(n292), .Y(n269) );
  NAND2X2 U195 ( .A(n313), .B(n262), .Y(n312) );
  NAND2X4 U196 ( .A(B[12]), .B(A[12]), .Y(n262) );
  AOI31X1 U197 ( .A0(n174), .A1(n175), .A2(n176), .B0(n177), .Y(n170) );
  NAND2X2 U198 ( .A(n79), .B(n74), .Y(n289) );
  NOR2X2 U199 ( .A(n184), .B(n150), .Y(n181) );
  INVX4 U200 ( .A(n163), .Y(n150) );
  NAND2X2 U201 ( .A(B[8]), .B(A[8]), .Y(n71) );
  NOR2BX2 U202 ( .AN(n117), .B(n116), .Y(n132) );
  NOR2X2 U203 ( .A(n69), .B(n76), .Y(n322) );
  INVX4 U204 ( .A(n294), .Y(n69) );
  OR2X4 U205 ( .A(A[10]), .B(B[10]), .Y(n296) );
  NOR2X4 U206 ( .A(n31), .B(n312), .Y(n310) );
  INVX8 U207 ( .A(n58), .Y(SUM[17]) );
  NAND2X2 U208 ( .A(n107), .B(n33), .Y(n34) );
  NAND2X4 U209 ( .A(n34), .B(n35), .Y(n345) );
  INVXL U210 ( .A(n107), .Y(n32) );
  NAND2X1 U211 ( .A(n94), .B(n99), .Y(n107) );
  NAND3BX1 U212 ( .AN(n100), .B(n102), .C(n101), .Y(n96) );
  NAND3BX1 U213 ( .AN(n100), .B(n102), .C(n101), .Y(n45) );
  NAND3BX1 U214 ( .AN(n100), .B(n102), .C(n101), .Y(n46) );
  NAND4BX4 U215 ( .AN(n338), .B(n339), .C(n134), .D(n133), .Y(n101) );
  OR2X1 U216 ( .A(A[24]), .B(B[24]), .Y(n163) );
  INVX1 U217 ( .A(n132), .Y(n48) );
  INVX1 U218 ( .A(n124), .Y(n123) );
  XOR2X4 U219 ( .A(n46), .B(n111), .Y(SUM[4]) );
  NOR2BX2 U220 ( .AN(n173), .B(n184), .Y(n197) );
  INVX8 U221 ( .A(n55), .Y(SUM[24]) );
  INVXL U222 ( .A(n87), .Y(n86) );
  INVX2 U223 ( .A(n237), .Y(n232) );
  XNOR2X4 U224 ( .A(n146), .B(n185), .Y(n55) );
  NAND2XL U225 ( .A(n47), .B(n132), .Y(n50) );
  NAND2X4 U226 ( .A(n49), .B(n50), .Y(SUM[2]) );
  XOR2X4 U227 ( .A(n137), .B(n138), .Y(SUM[29]) );
  AND2X1 U228 ( .A(n102), .B(n114), .Y(n113) );
  NAND2X2 U229 ( .A(B[23]), .B(A[23]), .Y(n173) );
  NAND2X1 U230 ( .A(B[27]), .B(A[27]), .Y(n143) );
  OR2X2 U231 ( .A(A[28]), .B(B[28]), .Y(n127) );
  NAND2X1 U232 ( .A(B[28]), .B(A[28]), .Y(n130) );
  NOR2X2 U233 ( .A(n85), .B(n86), .Y(n83) );
  XOR2X4 U234 ( .A(n36), .B(n37), .Y(SUM[30]) );
  NAND2XL U235 ( .A(n126), .B(n128), .Y(n137) );
  AND2X1 U236 ( .A(n95), .B(n94), .Y(n56) );
  AND2X2 U237 ( .A(n162), .B(n156), .Y(n38) );
  NAND3BX4 U238 ( .AN(n125), .B(n126), .C(n40), .Y(n121) );
  XNOR2X4 U239 ( .A(n300), .B(n41), .Y(n342) );
  AND2X2 U240 ( .A(n130), .B(n127), .Y(n144) );
  XOR2X4 U241 ( .A(n241), .B(n43), .Y(SUM[19]) );
  AND3X4 U242 ( .A(n219), .B(n218), .C(n217), .Y(n211) );
  OR2X4 U243 ( .A(A[22]), .B(B[22]), .Y(n178) );
  OR2X4 U244 ( .A(A[8]), .B(B[8]), .Y(n295) );
  NAND3X2 U245 ( .A(n217), .B(n218), .C(n235), .Y(n224) );
  NAND2XL U246 ( .A(B[22]), .B(A[22]), .Y(n204) );
  NOR2BX1 U247 ( .AN(n240), .B(n44), .Y(n346) );
  NOR2XL U248 ( .A(A[0]), .B(B[0]), .Y(n44) );
  INVX1 U249 ( .A(n156), .Y(n169) );
  XOR2X4 U250 ( .A(n51), .B(n318), .Y(n343) );
  XNOR2X4 U251 ( .A(n52), .B(n205), .Y(SUM[22]) );
  AND2X2 U252 ( .A(n178), .B(n204), .Y(n52) );
  NAND2XL U253 ( .A(n292), .B(n304), .Y(n309) );
  INVX1 U254 ( .A(n130), .Y(n140) );
  INVXL U255 ( .A(n106), .Y(n110) );
  NAND2X1 U256 ( .A(n156), .B(n155), .Y(n164) );
  NOR2BX2 U257 ( .AN(n236), .B(n233), .Y(n272) );
  NAND2XL U258 ( .A(n252), .B(n251), .Y(n273) );
  INVX1 U259 ( .A(n268), .Y(n275) );
  NOR2X2 U260 ( .A(n225), .B(n226), .Y(n234) );
  OAI21XL U261 ( .A0(n305), .A1(n262), .B0(n263), .Y(n257) );
  AOI21X1 U262 ( .A0(n88), .A1(n89), .B0(n75), .Y(n85) );
  NAND3XL U263 ( .A(n102), .B(n290), .C(n101), .Y(n287) );
  AND2X1 U264 ( .A(n79), .B(n80), .Y(n53) );
  XNOR2X4 U265 ( .A(n298), .B(n299), .Y(n54) );
  INVX8 U266 ( .A(n54), .Y(SUM[15]) );
  NAND3X4 U267 ( .A(n56), .B(n109), .C(n336), .Y(n84) );
  OAI21X2 U268 ( .A0(n211), .A1(n212), .B0(n213), .Y(n209) );
  NAND2XL U269 ( .A(n215), .B(n216), .Y(n212) );
  AND2X2 U270 ( .A(n142), .B(n143), .Y(n57) );
  INVXL U271 ( .A(n236), .Y(n266) );
  NAND2XL U272 ( .A(n237), .B(n215), .Y(n243) );
  NAND2X1 U273 ( .A(n98), .B(n99), .Y(n97) );
  NOR2BX2 U274 ( .AN(n68), .B(n69), .Y(n67) );
  NAND3X2 U275 ( .A(n70), .B(n71), .C(n72), .Y(n66) );
  XOR2X4 U276 ( .A(n59), .B(n264), .Y(n58) );
  AND2X1 U277 ( .A(n237), .B(n218), .Y(n59) );
  INVX1 U278 ( .A(n270), .Y(n258) );
  NAND2XL U279 ( .A(n99), .B(n98), .Y(n104) );
  NAND2X2 U280 ( .A(B[17]), .B(A[17]), .Y(n218) );
  NAND2X2 U281 ( .A(B[3]), .B(A[3]), .Y(n102) );
  NAND2X2 U282 ( .A(B[15]), .B(A[15]), .Y(n268) );
  NOR2X4 U283 ( .A(A[27]), .B(B[27]), .Y(n61) );
  NAND2X2 U284 ( .A(B[6]), .B(A[6]), .Y(n89) );
  OR2X2 U285 ( .A(A[29]), .B(B[29]), .Y(n128) );
  NAND2XL U286 ( .A(B[22]), .B(A[22]), .Y(n193) );
  OR2X2 U287 ( .A(A[30]), .B(B[30]), .Y(n122) );
  NOR2X4 U288 ( .A(A[5]), .B(B[5]), .Y(n62) );
  XNOR2X4 U289 ( .A(n324), .B(n8), .Y(n63) );
  INVX8 U290 ( .A(n63), .Y(SUM[11]) );
  NAND2X1 U291 ( .A(B[29]), .B(A[29]), .Y(n126) );
  NAND2X1 U292 ( .A(B[30]), .B(A[30]), .Y(n124) );
  NAND2X1 U293 ( .A(B[0]), .B(A[0]), .Y(n240) );
  XNOR2X1 U294 ( .A(B[31]), .B(A[31]), .Y(n119) );
  NAND3BX4 U295 ( .AN(n100), .B(n102), .C(n101), .Y(n109) );
  NAND2X1 U296 ( .A(B[7]), .B(A[7]), .Y(n87) );
  AOI21X1 U297 ( .A0(B[7]), .A1(A[7]), .B0(n75), .Y(n91) );
  INVX8 U298 ( .A(n293), .Y(n297) );
  NAND2XL U299 ( .A(n178), .B(n179), .Y(n177) );
  NOR2X2 U300 ( .A(A[15]), .B(B[15]), .Y(n281) );
  NAND2X1 U301 ( .A(n83), .B(n84), .Y(n81) );
  OAI21X2 U302 ( .A0(n300), .A1(n261), .B0(n270), .Y(n298) );
  NAND2XL U303 ( .A(B[18]), .B(A[18]), .Y(n235) );
  NAND2XL U304 ( .A(B[18]), .B(A[18]), .Y(n219) );
  NAND2X1 U305 ( .A(B[22]), .B(A[22]), .Y(n176) );
  AOI21X2 U306 ( .A0(n163), .A1(n146), .B0(n164), .Y(n159) );
  INVX4 U307 ( .A(n328), .Y(n326) );
  NAND2XL U308 ( .A(B[9]), .B(A[9]), .Y(n68) );
  NOR2X4 U309 ( .A(n275), .B(n276), .Y(n274) );
  INVX8 U310 ( .A(n308), .Y(n280) );
  NAND2XL U311 ( .A(n94), .B(n80), .Y(n93) );
  INVX8 U312 ( .A(n79), .Y(n75) );
  XOR2X4 U313 ( .A(n66), .B(n67), .Y(n344) );
  XOR2X4 U314 ( .A(n90), .B(n21), .Y(SUM[7]) );
  OAI21X4 U315 ( .A0(n92), .A1(n93), .B0(n89), .Y(n90) );
  XOR2X4 U316 ( .A(n103), .B(n12), .Y(SUM[6]) );
  NAND2BX4 U317 ( .AN(n104), .B(n105), .Y(n103) );
  CLKINVX3 U318 ( .A(n95), .Y(n78) );
  XOR2X4 U319 ( .A(n112), .B(n113), .Y(SUM[3]) );
  XOR2X4 U320 ( .A(n129), .B(n144), .Y(SUM[28]) );
  CLKINVX3 U321 ( .A(n154), .Y(n148) );
  XOR2X4 U322 ( .A(n157), .B(n158), .Y(n340) );
  OAI21X4 U323 ( .A0(n159), .A1(n160), .B0(n161), .Y(n157) );
  XOR2X4 U324 ( .A(n165), .B(n166), .Y(SUM[26]) );
  AND2X2 U325 ( .A(n155), .B(n173), .Y(n172) );
  OR2X4 U326 ( .A(A[26]), .B(B[26]), .Y(n154) );
  XOR2X4 U327 ( .A(n180), .B(n38), .Y(SUM[25]) );
  OAI2BB1X4 U328 ( .A0N(n181), .A1N(n182), .B0(n155), .Y(n180) );
  NAND2BX4 U329 ( .AN(n186), .B(n20), .Y(n146) );
  OAI2BB1X4 U330 ( .A0N(n192), .A1N(n183), .B0(n173), .Y(n186) );
  XOR2X4 U331 ( .A(n196), .B(n197), .Y(SUM[23]) );
  OR2X4 U332 ( .A(A[23]), .B(B[23]), .Y(n179) );
  AOI21X4 U333 ( .A0(n206), .A1(n207), .B0(n208), .Y(n205) );
  CLKINVX3 U334 ( .A(n175), .Y(n208) );
  XOR2X4 U335 ( .A(n221), .B(n220), .Y(n341) );
  OR2X4 U336 ( .A(A[21]), .B(B[21]), .Y(n191) );
  XOR2X4 U337 ( .A(n189), .B(n227), .Y(SUM[20]) );
  NAND2BX4 U338 ( .AN(n228), .B(n210), .Y(n189) );
  OAI2BB1X4 U339 ( .A0N(n234), .A1N(n224), .B0(n214), .Y(n228) );
  NAND2BX4 U340 ( .AN(n236), .B(n237), .Y(n217) );
  XOR2X4 U341 ( .A(n135), .B(n238), .Y(SUM[1]) );
  NOR2BX4 U342 ( .AN(n136), .B(n239), .Y(n238) );
  CLKINVX3 U343 ( .A(n134), .Y(n239) );
  OR2X4 U344 ( .A(n16), .B(B[19]), .Y(n216) );
  OAI21X4 U345 ( .A0(n242), .A1(n243), .B0(n244), .Y(n241) );
  OR2X4 U346 ( .A(A[18]), .B(B[18]), .Y(n215) );
  AOI21X4 U347 ( .A0(n245), .A1(n265), .B0(n266), .Y(n264) );
  OR2X4 U348 ( .A(A[17]), .B(B[17]), .Y(n237) );
  CLKINVX3 U349 ( .A(n245), .Y(n233) );
  OR2X4 U350 ( .A(A[16]), .B(B[16]), .Y(n245) );
  NAND3BX4 U351 ( .AN(n277), .B(n278), .C(n279), .Y(n249) );
  OR2X4 U352 ( .A(A[15]), .B(B[15]), .Y(n251) );
  NOR3X4 U353 ( .A(n301), .B(n302), .C(n303), .Y(n300) );
  NOR4BX4 U354 ( .AN(n285), .B(n305), .C(n280), .D(n297), .Y(n302) );
  OR2X4 U355 ( .A(A[14]), .B(B[14]), .Y(n252) );
  OR2X4 U356 ( .A(A[13]), .B(B[13]), .Y(n292) );
  OR2X4 U357 ( .A(A[12]), .B(B[12]), .Y(n308) );
  NAND3BX4 U358 ( .AN(n320), .B(n321), .C(n322), .Y(n306) );
  NAND3X4 U359 ( .A(n296), .B(n294), .C(n323), .Y(n317) );
  OR2X4 U360 ( .A(A[11]), .B(B[11]), .Y(n293) );
  OAI21X4 U361 ( .A0(n326), .A1(n327), .B0(n316), .Y(n324) );
  XOR2X4 U362 ( .A(n328), .B(n329), .Y(SUM[10]) );
  NAND2X4 U363 ( .A(n330), .B(n331), .Y(n328) );
  NAND3X4 U364 ( .A(n87), .B(n89), .C(n88), .Y(n74) );
  NAND3X4 U365 ( .A(n94), .B(n80), .C(n333), .Y(n88) );
  NAND2X4 U366 ( .A(B[5]), .B(A[5]), .Y(n99) );
  OR2X4 U367 ( .A(A[9]), .B(B[9]), .Y(n294) );
  NOR2X4 U368 ( .A(n337), .B(n75), .Y(n336) );
  OR2X4 U369 ( .A(A[7]), .B(B[7]), .Y(n79) );
  OR2X4 U370 ( .A(A[6]), .B(B[6]), .Y(n80) );
  OR2X4 U371 ( .A(A[4]), .B(B[4]), .Y(n95) );
endmodule


module hash_core_DW01_add_38 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n259, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258;

  INVX8 U2 ( .A(n177), .Y(n173) );
  NAND4BX4 U3 ( .AN(n176), .B(n177), .C(n178), .D(n179), .Y(n166) );
  NAND2X2 U4 ( .A(B[18]), .B(A[18]), .Y(n184) );
  NAND2X2 U5 ( .A(n144), .B(n2), .Y(n3) );
  NAND2X4 U6 ( .A(n1), .B(n145), .Y(n4) );
  NAND2X4 U7 ( .A(n3), .B(n4), .Y(SUM[25]) );
  INVX4 U8 ( .A(n144), .Y(n1) );
  INVX1 U9 ( .A(n145), .Y(n2) );
  OAI2BB1X4 U10 ( .A0N(n113), .A1N(n114), .B0(n140), .Y(n144) );
  AND2X2 U11 ( .A(n117), .B(n112), .Y(n145) );
  NAND2X2 U12 ( .A(n153), .B(n6), .Y(n7) );
  NAND2X4 U13 ( .A(n5), .B(n154), .Y(n8) );
  NAND2X4 U14 ( .A(n7), .B(n8), .Y(SUM[23]) );
  CLKINVX4 U15 ( .A(n153), .Y(n5) );
  CLKINVX4 U16 ( .A(n154), .Y(n6) );
  OAI2BB1X4 U17 ( .A0N(n155), .A1N(n129), .B0(n152), .Y(n153) );
  NOR2BX4 U18 ( .AN(n127), .B(n132), .Y(n154) );
  NOR2BX4 U19 ( .AN(n240), .B(n241), .Y(n234) );
  NAND2X2 U20 ( .A(B[10]), .B(A[10]), .Y(n240) );
  INVX1 U21 ( .A(n180), .Y(n199) );
  NAND2X2 U22 ( .A(n180), .B(n181), .Y(n176) );
  OR2X4 U23 ( .A(A[16]), .B(B[16]), .Y(n180) );
  NAND3BX4 U24 ( .AN(n219), .B(n220), .C(n221), .Y(n211) );
  AOI21X4 U25 ( .A0(n182), .A1(n177), .B0(n183), .Y(n165) );
  NOR2BX2 U26 ( .AN(n152), .B(n21), .Y(n156) );
  NOR2X4 U27 ( .A(n172), .B(n185), .Y(n182) );
  BUFX8 U28 ( .A(n208), .Y(n9) );
  NAND3BX4 U29 ( .AN(n23), .B(B[20]), .C(n150), .Y(n149) );
  INVX4 U30 ( .A(n238), .Y(n45) );
  BUFX4 U31 ( .A(n184), .Y(n10) );
  NAND2X4 U32 ( .A(n44), .B(n48), .Y(n239) );
  NAND2X4 U33 ( .A(B[9]), .B(A[9]), .Y(n44) );
  AOI21X4 U34 ( .A0(n191), .A1(n177), .B0(n192), .Y(n190) );
  INVX4 U35 ( .A(n218), .Y(n210) );
  NAND4BBX2 U36 ( .AN(n37), .BN(n39), .C(n58), .D(n252), .Y(n218) );
  BUFX4 U37 ( .A(n259), .Y(SUM[12]) );
  NOR2X4 U38 ( .A(n257), .B(n258), .Y(n255) );
  OAI21X2 U39 ( .A0(n187), .A1(n188), .B0(n103), .Y(n258) );
  NOR2BX1 U40 ( .AN(n62), .B(n39), .Y(n64) );
  NOR2X2 U41 ( .A(A[4]), .B(B[4]), .Y(n39) );
  AOI21X2 U42 ( .A0(n210), .A1(n215), .B0(n216), .Y(n213) );
  CLKINVX2 U43 ( .A(n217), .Y(n216) );
  CLKINVX4 U44 ( .A(n71), .Y(n257) );
  OAI2BB1X4 U45 ( .A0N(n60), .A1N(n26), .B0(n59), .Y(n56) );
  AND2X4 U46 ( .A(n59), .B(n62), .Y(n32) );
  NAND2X4 U47 ( .A(B[4]), .B(A[4]), .Y(n62) );
  CLKINVX8 U48 ( .A(n215), .Y(n253) );
  OAI21X4 U49 ( .A0(n255), .A1(n256), .B0(n67), .Y(n215) );
  INVX3 U50 ( .A(n98), .Y(n86) );
  NOR2BX2 U51 ( .AN(n117), .B(n15), .Y(n116) );
  INVX1 U52 ( .A(A[20]), .Y(n23) );
  NOR2BX2 U53 ( .AN(n175), .B(n199), .Y(n198) );
  INVXL U54 ( .A(n37), .Y(n26) );
  NAND2X2 U55 ( .A(n12), .B(n87), .Y(n134) );
  CLKINVX3 U56 ( .A(n152), .Y(n151) );
  NOR2X2 U57 ( .A(n174), .B(n175), .Y(n168) );
  INVX1 U58 ( .A(n171), .Y(n170) );
  NOR2X2 U59 ( .A(n172), .B(n10), .Y(n183) );
  NAND3X2 U60 ( .A(n38), .B(n87), .C(n88), .Y(n97) );
  NAND3BX2 U61 ( .AN(n21), .B(n147), .C(n128), .Y(n20) );
  OR2X2 U62 ( .A(A[12]), .B(B[12]), .Y(n220) );
  NAND2X1 U63 ( .A(n100), .B(n254), .Y(n256) );
  OR2X2 U64 ( .A(A[1]), .B(B[1]), .Y(n101) );
  INVX1 U65 ( .A(n88), .Y(n84) );
  NOR2X1 U66 ( .A(n79), .B(n13), .Y(n78) );
  OAI2BB1X1 U67 ( .A0N(B[28]), .A1N(A[28]), .B0(n80), .Y(n77) );
  NAND2BX1 U68 ( .AN(n13), .B(n75), .Y(n89) );
  OAI21X1 U69 ( .A0(n79), .A1(n92), .B0(n80), .Y(n91) );
  INVX4 U70 ( .A(n195), .Y(n194) );
  NAND3X1 U71 ( .A(n17), .B(n126), .C(n127), .Y(n123) );
  NAND2X1 U72 ( .A(B[26]), .B(A[26]), .Y(n12) );
  INVX1 U73 ( .A(A[13]), .Y(n18) );
  INVX1 U74 ( .A(n220), .Y(n229) );
  OR2X2 U75 ( .A(A[3]), .B(B[3]), .Y(n254) );
  NAND2X1 U76 ( .A(B[2]), .B(A[2]), .Y(n71) );
  INVX1 U77 ( .A(n101), .Y(n187) );
  NAND2X1 U78 ( .A(B[0]), .B(A[0]), .Y(n188) );
  XOR2X2 U79 ( .A(n195), .B(n196), .Y(SUM[17]) );
  NOR2BX1 U80 ( .AN(n27), .B(n174), .Y(n196) );
  XOR2X2 U81 ( .A(n157), .B(n159), .Y(SUM[21]) );
  NOR2BX1 U82 ( .AN(n140), .B(n138), .Y(n146) );
  XOR2X2 U83 ( .A(n50), .B(n51), .Y(SUM[7]) );
  NOR2X4 U84 ( .A(n19), .B(n142), .Y(n139) );
  NAND2X2 U85 ( .A(n20), .B(n127), .Y(n142) );
  NOR2BX1 U86 ( .AN(n9), .B(n40), .Y(n226) );
  NOR2BX1 U87 ( .AN(n48), .B(n49), .Y(n47) );
  INVX2 U88 ( .A(n46), .Y(n233) );
  XOR2X1 U89 ( .A(n46), .B(n47), .Y(SUM[8]) );
  INVX2 U90 ( .A(n129), .Y(n21) );
  OR2X2 U91 ( .A(A[26]), .B(B[26]), .Y(n87) );
  NOR2X1 U92 ( .A(A[26]), .B(B[26]), .Y(n111) );
  CLKINVX3 U93 ( .A(n113), .Y(n138) );
  INVX1 U94 ( .A(n253), .Y(n63) );
  NOR2X2 U95 ( .A(B[30]), .B(A[30]), .Y(n13) );
  AND2X2 U96 ( .A(n98), .B(n97), .Y(n14) );
  AND2X2 U97 ( .A(B[26]), .B(A[26]), .Y(n15) );
  NAND2X2 U98 ( .A(B[8]), .B(A[8]), .Y(n48) );
  OR2X2 U99 ( .A(n130), .B(n131), .Y(n17) );
  DLY1X1 U100 ( .A(n40), .Y(n16) );
  INVX4 U101 ( .A(n231), .Y(n230) );
  NOR2X2 U102 ( .A(n219), .B(n40), .Y(n202) );
  NAND2X2 U103 ( .A(n150), .B(n129), .Y(n130) );
  XOR2X2 U104 ( .A(n227), .B(n228), .Y(SUM[13]) );
  NOR2X2 U105 ( .A(B[27]), .B(A[27]), .Y(n120) );
  OR2X2 U106 ( .A(B[27]), .B(A[27]), .Y(n38) );
  OAI21XL U107 ( .A0(B[27]), .A1(A[27]), .B0(n87), .Y(n85) );
  NAND2X4 U108 ( .A(n14), .B(n82), .Y(n24) );
  XOR2X2 U109 ( .A(n161), .B(n163), .Y(SUM[20]) );
  NOR2X2 U110 ( .A(n132), .B(n133), .Y(n122) );
  OAI2BB1X2 U111 ( .A0N(n94), .A1N(n82), .B0(n35), .Y(n34) );
  NAND2X1 U112 ( .A(B[6]), .B(A[6]), .Y(n55) );
  NAND2X1 U113 ( .A(B[21]), .B(A[21]), .Y(n158) );
  NOR2BX1 U114 ( .AN(n10), .B(n173), .Y(n193) );
  OAI21X4 U115 ( .A0(n213), .A1(n209), .B0(n214), .Y(n212) );
  OAI2BB1X4 U116 ( .A0N(n234), .A1N(n235), .B0(n236), .Y(n214) );
  INVX4 U117 ( .A(n225), .Y(n224) );
  XOR2X4 U118 ( .A(n225), .B(n226), .Y(SUM[14]) );
  OAI2BB1X4 U119 ( .A0N(n227), .A1N(n36), .B0(n207), .Y(n225) );
  NAND2X4 U120 ( .A(n46), .B(n243), .Y(n30) );
  OAI21X2 U121 ( .A0(n54), .A1(n31), .B0(n55), .Y(n50) );
  INVXL U122 ( .A(n56), .Y(n54) );
  NOR2BX4 U123 ( .AN(n18), .B(B[13]), .Y(n41) );
  NOR3BX2 U124 ( .AN(n147), .B(n131), .C(n130), .Y(n19) );
  NOR3BX2 U125 ( .AN(n147), .B(n131), .C(n130), .Y(n141) );
  AOI21X2 U126 ( .A0(n81), .A1(n82), .B0(n83), .Y(n76) );
  NAND2X1 U127 ( .A(B[3]), .B(A[3]), .Y(n67) );
  NAND3BX2 U128 ( .AN(n21), .B(n147), .C(n128), .Y(n143) );
  NAND2X2 U129 ( .A(n179), .B(n180), .Y(n197) );
  AOI21X4 U130 ( .A0(n22), .A1(A[21]), .B0(n151), .Y(n148) );
  BUFX1 U131 ( .A(B[21]), .Y(n22) );
  OAI21X4 U132 ( .A0(n138), .A1(n139), .B0(n140), .Y(n136) );
  NAND2X4 U133 ( .A(n197), .B(n175), .Y(n195) );
  XOR2X4 U134 ( .A(n191), .B(n193), .Y(SUM[18]) );
  OAI21X2 U135 ( .A0(n76), .A1(n77), .B0(n78), .Y(n74) );
  NAND2X4 U136 ( .A(B[27]), .B(A[27]), .Y(n98) );
  XOR2X2 U137 ( .A(n42), .B(n43), .Y(SUM[9]) );
  NOR2X4 U138 ( .A(n41), .B(n40), .Y(n221) );
  OR2X2 U139 ( .A(A[8]), .B(B[8]), .Y(n243) );
  NAND2X1 U140 ( .A(B[15]), .B(A[15]), .Y(n205) );
  NAND2X2 U141 ( .A(n117), .B(n125), .Y(n124) );
  NOR2X4 U142 ( .A(A[15]), .B(B[15]), .Y(n219) );
  NOR2X4 U143 ( .A(A[14]), .B(B[14]), .Y(n40) );
  AOI21X4 U144 ( .A0(n202), .A1(n203), .B0(n204), .Y(n201) );
  OAI211X2 U145 ( .A0(n41), .A1(n206), .B0(n207), .C0(n9), .Y(n203) );
  NAND2BX4 U146 ( .AN(n211), .B(n212), .Y(n200) );
  XNOR2X4 U147 ( .A(n25), .B(n73), .Y(SUM[31]) );
  AND2X2 U148 ( .A(n74), .B(n75), .Y(n25) );
  NAND2XL U149 ( .A(B[17]), .B(A[17]), .Y(n27) );
  NAND2X4 U150 ( .A(B[5]), .B(A[5]), .Y(n59) );
  NOR2X4 U151 ( .A(A[5]), .B(B[5]), .Y(n37) );
  OR2X4 U152 ( .A(n249), .B(n45), .Y(n28) );
  NAND2X4 U153 ( .A(n28), .B(n44), .Y(n246) );
  INVXL U154 ( .A(n42), .Y(n249) );
  AOI21X4 U155 ( .A0(n237), .A1(n246), .B0(n247), .Y(n245) );
  NAND2X1 U156 ( .A(B[7]), .B(A[7]), .Y(n52) );
  NAND2X2 U157 ( .A(B[29]), .B(A[29]), .Y(n80) );
  NAND2X1 U158 ( .A(B[19]), .B(A[19]), .Y(n171) );
  AND2X1 U159 ( .A(n158), .B(n150), .Y(n159) );
  NOR2BXL U160 ( .AN(n205), .B(n219), .Y(n223) );
  OR2X2 U161 ( .A(A[2]), .B(B[2]), .Y(n100) );
  INVX2 U162 ( .A(n205), .Y(n204) );
  INVX4 U163 ( .A(n58), .Y(n31) );
  AOI21X4 U164 ( .A0(n112), .A1(n136), .B0(n137), .Y(n135) );
  AND2X2 U165 ( .A(n93), .B(n95), .Y(n35) );
  NOR2BX1 U166 ( .AN(n71), .B(n70), .Y(n99) );
  NOR2X2 U167 ( .A(n111), .B(n120), .Y(n110) );
  NAND2X1 U168 ( .A(B[1]), .B(A[1]), .Y(n103) );
  OAI21X4 U169 ( .A0(n39), .A1(n253), .B0(n62), .Y(n60) );
  XOR2X4 U170 ( .A(n89), .B(n29), .Y(SUM[30]) );
  NOR2X4 U171 ( .A(n90), .B(n91), .Y(n29) );
  NAND3BX4 U172 ( .AN(n141), .B(n127), .C(n143), .Y(n114) );
  CLKINVX3 U173 ( .A(n34), .Y(n90) );
  INVXL U174 ( .A(n117), .Y(n137) );
  AND2X1 U175 ( .A(n240), .B(n237), .Y(n248) );
  INVXL U176 ( .A(n240), .Y(n247) );
  NAND2X4 U177 ( .A(n30), .B(n48), .Y(n42) );
  OR3X4 U178 ( .A(n37), .B(n32), .C(n31), .Y(n251) );
  NOR2BXL U179 ( .AN(n207), .B(n41), .Y(n228) );
  INVXL U180 ( .A(n10), .Y(n192) );
  INVXL U181 ( .A(n254), .Y(n68) );
  INVXL U182 ( .A(n41), .Y(n36) );
  NAND2XL U183 ( .A(B[30]), .B(A[30]), .Y(n75) );
  AOI2BB1X2 U184 ( .A0N(n84), .A1N(n85), .B0(n86), .Y(n81) );
  NAND2XL U185 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NAND2XL U186 ( .A(B[20]), .B(A[20]), .Y(n160) );
  NOR2BX1 U187 ( .AN(n188), .B(n33), .Y(SUM[0]) );
  NOR2XL U188 ( .A(A[0]), .B(B[0]), .Y(n33) );
  NOR2BX1 U189 ( .AN(n206), .B(n229), .Y(n232) );
  XOR2X1 U190 ( .A(n56), .B(n57), .Y(SUM[6]) );
  NOR2BX1 U191 ( .AN(n55), .B(n31), .Y(n57) );
  XOR2X1 U192 ( .A(n60), .B(n61), .Y(SUM[5]) );
  NOR2BX1 U193 ( .AN(n59), .B(n37), .Y(n61) );
  NOR2BXL U194 ( .AN(n52), .B(n53), .Y(n51) );
  NOR2BX1 U195 ( .AN(n44), .B(n45), .Y(n43) );
  NAND2XL U196 ( .A(n171), .B(n178), .Y(n189) );
  NAND2XL U197 ( .A(n93), .B(n80), .Y(n104) );
  INVX1 U198 ( .A(n107), .Y(n106) );
  NAND3X2 U199 ( .A(n237), .B(n238), .C(n239), .Y(n235) );
  INVXL U200 ( .A(n147), .Y(n132) );
  XOR2X1 U201 ( .A(n65), .B(n66), .Y(SUM[3]) );
  OAI21XL U202 ( .A0(n69), .A1(n70), .B0(n71), .Y(n65) );
  NOR2BX1 U203 ( .AN(n67), .B(n68), .Y(n66) );
  INVX1 U204 ( .A(n72), .Y(n69) );
  XOR2X1 U205 ( .A(n72), .B(n99), .Y(SUM[2]) );
  XOR2X1 U206 ( .A(n63), .B(n64), .Y(SUM[4]) );
  XOR2X1 U207 ( .A(n102), .B(n186), .Y(SUM[1]) );
  NOR2BXL U208 ( .AN(n103), .B(n187), .Y(n186) );
  INVX1 U209 ( .A(n100), .Y(n70) );
  OAI2BB1X1 U210 ( .A0N(n101), .A1N(n102), .B0(n103), .Y(n72) );
  INVX1 U211 ( .A(n188), .Y(n102) );
  XOR2X1 U212 ( .A(B[31]), .B(A[31]), .Y(n73) );
  NAND2X2 U213 ( .A(B[13]), .B(A[13]), .Y(n207) );
  NAND2XL U214 ( .A(B[28]), .B(A[28]), .Y(n107) );
  NAND2XL U215 ( .A(A[28]), .B(B[28]), .Y(n92) );
  NAND2X4 U216 ( .A(n200), .B(n201), .Y(n179) );
  XOR2X1 U217 ( .A(n179), .B(n198), .Y(SUM[16]) );
  NAND2X2 U218 ( .A(B[23]), .B(A[23]), .Y(n127) );
  NAND2X1 U219 ( .A(n128), .B(n129), .Y(n126) );
  OR2X4 U220 ( .A(A[22]), .B(B[22]), .Y(n129) );
  NAND2X2 U221 ( .A(B[24]), .B(A[24]), .Y(n140) );
  OAI2BB1X2 U222 ( .A0N(n115), .A1N(n112), .B0(n116), .Y(n88) );
  XOR2X2 U223 ( .A(n114), .B(n146), .Y(SUM[24]) );
  NAND2X2 U224 ( .A(B[25]), .B(A[25]), .Y(n117) );
  NAND2X2 U225 ( .A(B[14]), .B(A[14]), .Y(n208) );
  INVX8 U226 ( .A(n181), .Y(n174) );
  NAND3X1 U227 ( .A(n112), .B(n113), .C(n114), .Y(n109) );
  NAND2X2 U228 ( .A(B[16]), .B(A[16]), .Y(n175) );
  XOR2X1 U229 ( .A(n231), .B(n232), .Y(n259) );
  NAND2XL U230 ( .A(n236), .B(n242), .Y(n244) );
  NAND2X1 U231 ( .A(n113), .B(n112), .Y(n133) );
  INVX8 U232 ( .A(n178), .Y(n172) );
  AND2X1 U233 ( .A(A[24]), .B(B[24]), .Y(n115) );
  NAND3X1 U234 ( .A(A[24]), .B(B[24]), .C(n112), .Y(n125) );
  CLKINVX3 U235 ( .A(n93), .Y(n79) );
  NOR2X4 U236 ( .A(n86), .B(n96), .Y(n94) );
  CLKINVX3 U237 ( .A(n97), .Y(n96) );
  XOR2X4 U238 ( .A(n104), .B(n105), .Y(SUM[29]) );
  AOI21X4 U239 ( .A0(n24), .A1(n95), .B0(n106), .Y(n105) );
  OR2X4 U240 ( .A(A[29]), .B(B[29]), .Y(n93) );
  XOR2X4 U241 ( .A(n24), .B(n108), .Y(SUM[28]) );
  NOR2BX4 U242 ( .AN(n107), .B(n83), .Y(n108) );
  CLKINVX3 U243 ( .A(n95), .Y(n83) );
  OR2X4 U244 ( .A(A[28]), .B(B[28]), .Y(n95) );
  NAND2BX4 U245 ( .AN(n109), .B(n110), .Y(n82) );
  XOR2X4 U246 ( .A(n118), .B(n119), .Y(SUM[27]) );
  NOR2BX4 U247 ( .AN(n98), .B(n120), .Y(n119) );
  OAI21X4 U248 ( .A0(n121), .A1(n111), .B0(n12), .Y(n118) );
  AOI21X4 U249 ( .A0(n122), .A1(n123), .B0(n124), .Y(n121) );
  XOR2X4 U250 ( .A(n135), .B(n134), .Y(SUM[26]) );
  OR2X4 U251 ( .A(B[25]), .B(A[25]), .Y(n112) );
  OR2X4 U252 ( .A(A[24]), .B(B[24]), .Y(n113) );
  NAND2X4 U253 ( .A(n148), .B(n149), .Y(n128) );
  OR2X4 U254 ( .A(A[23]), .B(B[23]), .Y(n147) );
  XOR2X4 U255 ( .A(n155), .B(n156), .Y(SUM[22]) );
  NAND2X4 U256 ( .A(B[22]), .B(A[22]), .Y(n152) );
  OAI2BB1X4 U257 ( .A0N(n150), .A1N(n157), .B0(n158), .Y(n155) );
  OR2X4 U258 ( .A(A[21]), .B(B[21]), .Y(n150) );
  NAND2X4 U259 ( .A(n131), .B(n160), .Y(n157) );
  NAND2X4 U260 ( .A(n161), .B(n162), .Y(n131) );
  NOR2BX4 U261 ( .AN(n160), .B(n164), .Y(n163) );
  CLKINVX3 U262 ( .A(n162), .Y(n164) );
  OR2X4 U263 ( .A(A[20]), .B(B[20]), .Y(n162) );
  NAND3X4 U264 ( .A(n165), .B(n166), .C(n167), .Y(n161) );
  AOI21X4 U265 ( .A0(n169), .A1(n168), .B0(n170), .Y(n167) );
  NOR2X4 U266 ( .A(n172), .B(n173), .Y(n169) );
  XOR2X4 U267 ( .A(n189), .B(n190), .Y(SUM[19]) );
  OR2X4 U268 ( .A(A[19]), .B(B[19]), .Y(n178) );
  OR2X4 U269 ( .A(A[18]), .B(B[18]), .Y(n177) );
  OAI21X4 U270 ( .A0(n194), .A1(n174), .B0(n27), .Y(n191) );
  OR2X4 U271 ( .A(A[17]), .B(B[17]), .Y(n181) );
  XOR2X4 U272 ( .A(n222), .B(n223), .Y(SUM[15]) );
  OAI21X4 U273 ( .A0(n224), .A1(n16), .B0(n9), .Y(n222) );
  OAI21X4 U274 ( .A0(n229), .A1(n230), .B0(n206), .Y(n227) );
  NAND2X4 U275 ( .A(B[12]), .B(A[12]), .Y(n206) );
  OAI21X4 U276 ( .A0(n233), .A1(n209), .B0(n214), .Y(n231) );
  CLKINVX3 U277 ( .A(n242), .Y(n241) );
  NAND4BBX4 U278 ( .AN(n49), .BN(n45), .C(n237), .D(n236), .Y(n209) );
  CLKINVX3 U279 ( .A(n243), .Y(n49) );
  XOR2X4 U280 ( .A(n244), .B(n245), .Y(SUM[11]) );
  NAND2X4 U281 ( .A(B[11]), .B(A[11]), .Y(n242) );
  OR2X4 U282 ( .A(A[11]), .B(B[11]), .Y(n236) );
  XOR2X4 U283 ( .A(n246), .B(n248), .Y(SUM[10]) );
  OR2X4 U284 ( .A(A[10]), .B(B[10]), .Y(n237) );
  OR2X4 U285 ( .A(A[9]), .B(B[9]), .Y(n238) );
  OAI21X4 U286 ( .A0(n253), .A1(n218), .B0(n217), .Y(n46) );
  NAND2BX4 U287 ( .AN(n53), .B(n250), .Y(n217) );
  NAND3X4 U288 ( .A(n251), .B(n55), .C(n52), .Y(n250) );
  CLKINVX3 U289 ( .A(n252), .Y(n53) );
  OR2X4 U290 ( .A(A[7]), .B(B[7]), .Y(n252) );
  OR2X4 U291 ( .A(A[6]), .B(B[6]), .Y(n58) );
endmodule


module hash_core_DW01_add_40 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n274, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273;

  INVX2 U2 ( .A(n257), .Y(n256) );
  NAND2X2 U3 ( .A(n142), .B(n158), .Y(n157) );
  AOI21X4 U4 ( .A0(n218), .A1(n219), .B0(n220), .Y(n217) );
  CLKINVX8 U5 ( .A(n211), .Y(n210) );
  NAND2X2 U6 ( .A(n29), .B(n127), .Y(n30) );
  NOR2X4 U7 ( .A(n24), .B(n138), .Y(n134) );
  NAND2X4 U8 ( .A(B[13]), .B(A[13]), .Y(n223) );
  NAND2X1 U9 ( .A(A[24]), .B(B[24]), .Y(n1) );
  NAND2X2 U10 ( .A(n2), .B(n125), .Y(n139) );
  CLKINVX3 U11 ( .A(n1), .Y(n2) );
  NAND2X4 U12 ( .A(n37), .B(n4), .Y(n5) );
  NAND2X2 U13 ( .A(n3), .B(n206), .Y(n6) );
  NAND2X4 U14 ( .A(n5), .B(n6), .Y(SUM[19]) );
  CLKINVX2 U15 ( .A(n37), .Y(n3) );
  INVX4 U16 ( .A(n206), .Y(n4) );
  NAND2X2 U17 ( .A(n261), .B(n8), .Y(n9) );
  NAND2X2 U18 ( .A(n7), .B(n263), .Y(n10) );
  NAND2X4 U19 ( .A(n9), .B(n10), .Y(SUM[10]) );
  INVX2 U20 ( .A(n261), .Y(n7) );
  INVX1 U21 ( .A(n263), .Y(n8) );
  NAND2X1 U22 ( .A(A[18]), .B(B[18]), .Y(n201) );
  NAND2X2 U23 ( .A(n132), .B(n12), .Y(n13) );
  NAND2X4 U24 ( .A(n11), .B(n133), .Y(n14) );
  NAND2X4 U25 ( .A(n13), .B(n14), .Y(SUM[27]) );
  CLKINVX8 U26 ( .A(n132), .Y(n11) );
  INVX2 U27 ( .A(n133), .Y(n12) );
  CLKINVX3 U28 ( .A(n221), .Y(n220) );
  NAND2X2 U29 ( .A(B[15]), .B(A[15]), .Y(n221) );
  OAI21X4 U30 ( .A0(n153), .A1(n154), .B0(n155), .Y(n151) );
  OAI2BB1XL U31 ( .A0N(n112), .A1N(n113), .B0(n114), .Y(n82) );
  OAI21X2 U32 ( .A0(n204), .A1(n205), .B0(n114), .Y(n273) );
  NAND2X2 U33 ( .A(B[26]), .B(A[26]), .Y(n135) );
  BUFX4 U34 ( .A(n73), .Y(n15) );
  OR2X4 U35 ( .A(B[27]), .B(A[27]), .Y(n46) );
  NOR2X4 U36 ( .A(B[27]), .B(A[27]), .Y(n124) );
  NAND2X4 U37 ( .A(B[27]), .B(A[27]), .Y(n109) );
  NOR2X2 U38 ( .A(n123), .B(n124), .Y(n122) );
  NAND3X1 U39 ( .A(n125), .B(n126), .C(n127), .Y(n121) );
  CLKINVX3 U40 ( .A(n198), .Y(n192) );
  BUFX4 U41 ( .A(n201), .Y(n34) );
  NAND3X2 U42 ( .A(n51), .B(n235), .C(n236), .Y(n227) );
  NAND2BX2 U43 ( .AN(n48), .B(n84), .Y(n98) );
  NAND2X2 U44 ( .A(n30), .B(n155), .Y(n159) );
  NOR2X2 U45 ( .A(n190), .B(n34), .Y(n200) );
  INVX1 U46 ( .A(A[20]), .Y(n18) );
  NAND3X1 U47 ( .A(n252), .B(n253), .C(n254), .Y(n250) );
  NOR2BX2 U48 ( .AN(n255), .B(n256), .Y(n249) );
  NAND2X1 U49 ( .A(n130), .B(n139), .Y(n138) );
  INVX1 U50 ( .A(n171), .Y(n17) );
  CLKINVX3 U51 ( .A(n237), .Y(n25) );
  NAND2X2 U52 ( .A(n196), .B(n197), .Y(n213) );
  INVX1 U53 ( .A(n20), .Y(n21) );
  NAND2X2 U54 ( .A(n36), .B(n58), .Y(n52) );
  OAI2BB1X1 U55 ( .A0N(B[28]), .A1N(A[28]), .B0(n89), .Y(n86) );
  NAND2X1 U56 ( .A(n111), .B(n269), .Y(n271) );
  NOR2X1 U57 ( .A(n272), .B(n273), .Y(n270) );
  INVX1 U58 ( .A(n103), .Y(n88) );
  NOR2X1 U59 ( .A(n95), .B(n107), .Y(n104) );
  OR2X2 U60 ( .A(A[29]), .B(B[29]), .Y(n103) );
  INVX1 U61 ( .A(n153), .Y(n29) );
  NOR2BX1 U62 ( .AN(n168), .B(n171), .Y(n173) );
  NOR2BX1 U63 ( .AN(n114), .B(n204), .Y(n203) );
  NOR2BX1 U64 ( .AN(n224), .B(n49), .Y(n240) );
  BUFX3 U65 ( .A(n274), .Y(SUM[13]) );
  NOR2BX1 U66 ( .AN(n155), .B(n153), .Y(n162) );
  INVX1 U67 ( .A(n34), .Y(n208) );
  NOR2BX1 U68 ( .AN(n34), .B(n191), .Y(n209) );
  INVX1 U69 ( .A(n255), .Y(n262) );
  XOR2X2 U70 ( .A(n174), .B(n176), .Y(SUM[21]) );
  NOR2BX2 U71 ( .AN(n175), .B(n177), .Y(n176) );
  XOR2X1 U72 ( .A(n70), .B(n71), .Y(SUM[5]) );
  XOR2X1 U73 ( .A(n75), .B(n76), .Y(SUM[3]) );
  NAND2X1 U74 ( .A(n135), .B(n96), .Y(n149) );
  NOR2BX1 U75 ( .AN(n193), .B(n215), .Y(n214) );
  INVX1 U76 ( .A(n197), .Y(n215) );
  XOR2X2 U77 ( .A(n60), .B(n61), .Y(SUM[7]) );
  NOR2BX1 U78 ( .AN(n65), .B(n64), .Y(n67) );
  NAND2X2 U79 ( .A(B[14]), .B(A[14]), .Y(n224) );
  OR2X2 U80 ( .A(A[26]), .B(B[26]), .Y(n96) );
  NOR2X1 U81 ( .A(A[26]), .B(B[26]), .Y(n123) );
  AND2X2 U82 ( .A(n109), .B(n108), .Y(n16) );
  AOI21X4 U83 ( .A0(B[21]), .A1(A[21]), .B0(n167), .Y(n164) );
  INVX2 U84 ( .A(n168), .Y(n167) );
  NOR2BX2 U85 ( .AN(n119), .B(n92), .Y(n120) );
  NAND2X1 U86 ( .A(B[28]), .B(A[28]), .Y(n119) );
  INVX1 U87 ( .A(n144), .Y(n19) );
  OR2X2 U88 ( .A(A[15]), .B(B[15]), .Y(n51) );
  AOI21X4 U89 ( .A0(n199), .A1(n194), .B0(n200), .Y(n183) );
  NOR2BX4 U90 ( .AN(n109), .B(n124), .Y(n133) );
  OAI2BB1X4 U91 ( .A0N(n172), .A1N(n17), .B0(n168), .Y(n169) );
  INVX2 U92 ( .A(n97), .Y(n93) );
  NOR2BX4 U93 ( .AN(n163), .B(n148), .Y(n136) );
  INVXL U94 ( .A(n166), .Y(n177) );
  NAND3BX4 U95 ( .AN(n18), .B(B[20]), .C(n166), .Y(n165) );
  NOR2X2 U96 ( .A(n145), .B(n146), .Y(n140) );
  NOR2BX1 U97 ( .AN(n178), .B(n182), .Y(n181) );
  NAND2X1 U98 ( .A(B[20]), .B(A[20]), .Y(n178) );
  NAND2X4 U99 ( .A(n16), .B(n91), .Y(n117) );
  NAND2X4 U100 ( .A(n126), .B(n125), .Y(n148) );
  NOR2X4 U101 ( .A(n190), .B(n202), .Y(n199) );
  NAND2X1 U102 ( .A(n143), .B(n144), .Y(n141) );
  NOR2X1 U103 ( .A(A[4]), .B(B[4]), .Y(n45) );
  NAND3X4 U104 ( .A(n266), .B(n65), .C(n62), .Y(n265) );
  NAND2X1 U105 ( .A(B[7]), .B(A[7]), .Y(n62) );
  NAND3BX4 U106 ( .AN(n19), .B(n163), .C(n143), .Y(n158) );
  INVX1 U107 ( .A(n144), .Y(n171) );
  INVXL U108 ( .A(n179), .Y(n20) );
  INVX2 U109 ( .A(n109), .Y(n95) );
  INVX4 U110 ( .A(n126), .Y(n153) );
  OR2X4 U111 ( .A(A[24]), .B(B[24]), .Y(n126) );
  NAND4X2 U112 ( .A(n196), .B(n194), .C(n195), .D(n22), .Y(n184) );
  AND2X2 U113 ( .A(n197), .B(n198), .Y(n22) );
  XOR2X2 U114 ( .A(n172), .B(n173), .Y(SUM[22]) );
  CLKBUFX4 U115 ( .A(n50), .Y(n23) );
  INVX4 U116 ( .A(n268), .Y(n63) );
  OR2X4 U117 ( .A(A[7]), .B(B[7]), .Y(n268) );
  NOR2BXL U118 ( .AN(n62), .B(n63), .Y(n61) );
  OR2X4 U119 ( .A(A[12]), .B(B[12]), .Y(n235) );
  OR2X4 U120 ( .A(A[11]), .B(B[11]), .Y(n251) );
  OAI2BB1X4 U121 ( .A0N(n249), .A1N(n250), .B0(n251), .Y(n230) );
  NOR2BX1 U122 ( .AN(n202), .B(n192), .Y(n212) );
  NAND2X2 U123 ( .A(B[17]), .B(A[17]), .Y(n202) );
  NOR2BX2 U124 ( .AN(n54), .B(n55), .Y(n53) );
  INVX3 U125 ( .A(n253), .Y(n55) );
  NAND2X1 U126 ( .A(n103), .B(n89), .Y(n115) );
  XOR2X2 U127 ( .A(n239), .B(n240), .Y(SUM[14]) );
  OAI21X2 U128 ( .A0(n85), .A1(n86), .B0(n87), .Y(n83) );
  NOR2X4 U129 ( .A(n31), .B(n92), .Y(n85) );
  NOR2BX1 U130 ( .AN(n221), .B(n47), .Y(n238) );
  AND2X4 U131 ( .A(n136), .B(n137), .Y(n24) );
  NAND2X4 U132 ( .A(n237), .B(n26), .Y(n27) );
  NAND2X4 U133 ( .A(n25), .B(n238), .Y(n28) );
  NAND2X4 U134 ( .A(n27), .B(n28), .Y(SUM[15]) );
  INVX2 U135 ( .A(n238), .Y(n26) );
  NAND2X4 U136 ( .A(B[24]), .B(A[24]), .Y(n155) );
  AND2X4 U137 ( .A(n90), .B(n91), .Y(n31) );
  AOI2BB1X2 U138 ( .A0N(n93), .A1N(n94), .B0(n95), .Y(n90) );
  INVX4 U139 ( .A(n106), .Y(n92) );
  NAND2X4 U140 ( .A(n239), .B(n32), .Y(n33) );
  NAND2X4 U141 ( .A(n33), .B(n224), .Y(n237) );
  INVX12 U142 ( .A(n49), .Y(n32) );
  NOR2X2 U143 ( .A(A[15]), .B(B[15]), .Y(n47) );
  NAND2BX4 U144 ( .AN(n227), .B(n228), .Y(n216) );
  OAI21X2 U145 ( .A0(n229), .A1(n225), .B0(n230), .Y(n228) );
  OAI21X2 U146 ( .A0(n45), .A1(n72), .B0(n15), .Y(n70) );
  INVX3 U147 ( .A(n111), .Y(n80) );
  OR2X2 U148 ( .A(A[2]), .B(B[2]), .Y(n111) );
  OR2X4 U149 ( .A(A[8]), .B(B[8]), .Y(n258) );
  NOR2X4 U150 ( .A(A[14]), .B(B[14]), .Y(n49) );
  OAI21X2 U151 ( .A0(n88), .A1(n102), .B0(n89), .Y(n101) );
  NAND2X1 U152 ( .A(B[29]), .B(A[29]), .Y(n89) );
  OAI211X2 U153 ( .A0(n50), .A1(n222), .B0(n223), .C0(n224), .Y(n219) );
  XOR2X2 U154 ( .A(n127), .B(n162), .Y(SUM[24]) );
  OAI21X2 U155 ( .A0(n41), .A1(n64), .B0(n65), .Y(n60) );
  NAND2X1 U156 ( .A(B[6]), .B(A[6]), .Y(n65) );
  NAND3BX2 U157 ( .AN(n140), .B(n141), .C(n142), .Y(n137) );
  NOR2X1 U158 ( .A(n88), .B(n48), .Y(n87) );
  NOR2X2 U159 ( .A(A[30]), .B(B[30]), .Y(n48) );
  OAI21X4 U160 ( .A0(n264), .A1(n55), .B0(n54), .Y(n261) );
  NAND2X2 U161 ( .A(B[9]), .B(A[9]), .Y(n54) );
  NOR2X2 U162 ( .A(n47), .B(n49), .Y(n218) );
  NAND2X2 U163 ( .A(n69), .B(n15), .Y(n267) );
  XOR2X2 U164 ( .A(n66), .B(n67), .Y(SUM[6]) );
  NOR2X4 U165 ( .A(n192), .B(n193), .Y(n186) );
  NAND2X4 U166 ( .A(B[22]), .B(A[22]), .Y(n168) );
  AOI21X2 U167 ( .A0(n104), .A1(n91), .B0(n105), .Y(n100) );
  NAND2X4 U168 ( .A(B[5]), .B(A[5]), .Y(n69) );
  NOR2X4 U169 ( .A(A[5]), .B(B[5]), .Y(n44) );
  INVX4 U170 ( .A(n235), .Y(n244) );
  NAND2X2 U171 ( .A(n54), .B(n58), .Y(n254) );
  INVXL U172 ( .A(n233), .Y(n232) );
  INVXL U173 ( .A(n234), .Y(n226) );
  INVXL U174 ( .A(n69), .Y(n43) );
  NOR2BX1 U175 ( .AN(n77), .B(n78), .Y(n76) );
  NAND2X2 U176 ( .A(B[25]), .B(A[25]), .Y(n130) );
  AOI21X2 U177 ( .A0(n70), .A1(n42), .B0(n43), .Y(n41) );
  INVX2 U178 ( .A(n44), .Y(n42) );
  NOR2BXL U179 ( .AN(n69), .B(n44), .Y(n71) );
  AND2X1 U180 ( .A(n255), .B(n252), .Y(n263) );
  INVX1 U181 ( .A(n130), .Y(n152) );
  NOR2BX1 U182 ( .AN(n81), .B(n80), .Y(n110) );
  OAI21XL U183 ( .A0(n79), .A1(n80), .B0(n81), .Y(n75) );
  NAND3X4 U184 ( .A(n46), .B(n96), .C(n97), .Y(n108) );
  NAND2X2 U185 ( .A(B[16]), .B(A[16]), .Y(n193) );
  NAND2XL U186 ( .A(B[3]), .B(A[3]), .Y(n77) );
  NAND2XL U187 ( .A(B[1]), .B(A[1]), .Y(n114) );
  INVX4 U188 ( .A(n231), .Y(n72) );
  OAI21X4 U189 ( .A0(n270), .A1(n271), .B0(n77), .Y(n231) );
  XOR2X4 U190 ( .A(n150), .B(n149), .Y(SUM[26]) );
  NAND2X4 U191 ( .A(n56), .B(n258), .Y(n36) );
  NOR2BXL U192 ( .AN(n223), .B(n23), .Y(n243) );
  NAND2XL U193 ( .A(n189), .B(n195), .Y(n37) );
  INVX1 U194 ( .A(n41), .Y(n66) );
  NAND2XL U195 ( .A(B[4]), .B(A[4]), .Y(n73) );
  OR2X4 U196 ( .A(A[3]), .B(B[3]), .Y(n269) );
  OR2X4 U197 ( .A(A[17]), .B(B[17]), .Y(n198) );
  NAND2X1 U198 ( .A(B[19]), .B(A[19]), .Y(n189) );
  NAND2X4 U199 ( .A(B[11]), .B(A[11]), .Y(n257) );
  NAND2X4 U200 ( .A(B[12]), .B(A[12]), .Y(n222) );
  NAND2X2 U201 ( .A(B[2]), .B(A[2]), .Y(n81) );
  NAND2X2 U202 ( .A(B[0]), .B(A[0]), .Y(n205) );
  OR2X4 U203 ( .A(A[1]), .B(B[1]), .Y(n112) );
  NOR2BX1 U204 ( .AN(n205), .B(n38), .Y(SUM[0]) );
  NOR2XL U205 ( .A(A[0]), .B(B[0]), .Y(n38) );
  XOR2X4 U206 ( .A(n39), .B(n40), .Y(SUM[31]) );
  AND2X2 U207 ( .A(n83), .B(n84), .Y(n39) );
  XNOR2X1 U208 ( .A(B[31]), .B(A[31]), .Y(n40) );
  AOI21X1 U209 ( .A0(n226), .A1(n231), .B0(n232), .Y(n229) );
  NOR2BX1 U210 ( .AN(n222), .B(n244), .Y(n247) );
  INVX1 U211 ( .A(n52), .Y(n264) );
  INVX1 U212 ( .A(n81), .Y(n272) );
  XOR2X1 U213 ( .A(n56), .B(n57), .Y(SUM[8]) );
  NOR2BX1 U214 ( .AN(n58), .B(n59), .Y(n57) );
  XOR2X1 U215 ( .A(n242), .B(n243), .Y(n274) );
  XOR2X2 U216 ( .A(n211), .B(n212), .Y(SUM[17]) );
  XOR2X1 U217 ( .A(n52), .B(n53), .Y(SUM[9]) );
  XOR2X1 U218 ( .A(n231), .B(n74), .Y(SUM[4]) );
  NOR2BX1 U219 ( .AN(n15), .B(n45), .Y(n74) );
  INVX1 U220 ( .A(n119), .Y(n118) );
  NAND4BBX2 U221 ( .AN(n44), .BN(n45), .C(n68), .D(n268), .Y(n234) );
  INVXL U222 ( .A(n68), .Y(n64) );
  INVXL U223 ( .A(n163), .Y(n147) );
  INVXL U224 ( .A(n125), .Y(n161) );
  NOR2BX2 U225 ( .AN(n142), .B(n147), .Y(n170) );
  NAND2XL U226 ( .A(n103), .B(n106), .Y(n105) );
  INVX1 U227 ( .A(n108), .Y(n107) );
  INVX1 U228 ( .A(n258), .Y(n59) );
  INVX1 U229 ( .A(n189), .Y(n188) );
  INVX1 U230 ( .A(n82), .Y(n79) );
  XOR2X1 U231 ( .A(n82), .B(n110), .Y(SUM[2]) );
  INVX1 U232 ( .A(n269), .Y(n78) );
  NAND2XL U233 ( .A(B[21]), .B(A[21]), .Y(n175) );
  NAND2X2 U234 ( .A(B[8]), .B(A[8]), .Y(n58) );
  INVX1 U235 ( .A(n112), .Y(n204) );
  NAND2X2 U236 ( .A(B[10]), .B(A[10]), .Y(n255) );
  NAND2XL U237 ( .A(B[30]), .B(A[30]), .Y(n84) );
  AND2X2 U238 ( .A(n130), .B(n131), .Y(n129) );
  NOR2X4 U239 ( .A(A[13]), .B(B[13]), .Y(n50) );
  NAND2XL U240 ( .A(A[28]), .B(B[28]), .Y(n102) );
  XOR2X1 U241 ( .A(n113), .B(n203), .Y(SUM[1]) );
  INVX1 U242 ( .A(n205), .Y(n113) );
  NAND2X4 U243 ( .A(n217), .B(n216), .Y(n196) );
  XOR2X1 U244 ( .A(n246), .B(n247), .Y(SUM[12]) );
  NAND2X2 U245 ( .A(B[23]), .B(A[23]), .Y(n142) );
  NAND2X1 U246 ( .A(B[26]), .B(A[26]), .Y(n131) );
  OAI21XL U247 ( .A0(B[27]), .A1(A[27]), .B0(n96), .Y(n94) );
  NAND2X2 U248 ( .A(n166), .B(n144), .Y(n145) );
  NAND2XL U249 ( .A(n251), .B(n257), .Y(n259) );
  XOR2X1 U250 ( .A(n21), .B(n181), .Y(SUM[20]) );
  NOR2X2 U251 ( .A(n156), .B(n157), .Y(n154) );
  INVX4 U252 ( .A(n246), .Y(n245) );
  XOR2X1 U253 ( .A(n196), .B(n214), .Y(SUM[16]) );
  AND2X1 U254 ( .A(A[24]), .B(B[24]), .Y(n128) );
  INVX8 U255 ( .A(n194), .Y(n191) );
  INVX4 U256 ( .A(n242), .Y(n241) );
  INVX8 U257 ( .A(n195), .Y(n190) );
  XOR2X4 U258 ( .A(n98), .B(n99), .Y(SUM[30]) );
  NOR2X4 U259 ( .A(n100), .B(n101), .Y(n99) );
  XOR2X4 U260 ( .A(n115), .B(n116), .Y(SUM[29]) );
  AOI21X4 U261 ( .A0(n117), .A1(n106), .B0(n118), .Y(n116) );
  XOR2X4 U262 ( .A(n117), .B(n120), .Y(SUM[28]) );
  OR2X4 U263 ( .A(A[28]), .B(B[28]), .Y(n106) );
  NAND2BX4 U264 ( .AN(n121), .B(n122), .Y(n91) );
  OAI2BB1X4 U265 ( .A0N(n128), .A1N(n125), .B0(n129), .Y(n97) );
  OAI21X4 U266 ( .A0(n134), .A1(n123), .B0(n135), .Y(n132) );
  AOI21X4 U267 ( .A0(n125), .A1(n151), .B0(n152), .Y(n150) );
  XOR2X4 U268 ( .A(n159), .B(n160), .Y(SUM[25]) );
  NOR2BX4 U269 ( .AN(n130), .B(n161), .Y(n160) );
  OR2X4 U270 ( .A(B[25]), .B(A[25]), .Y(n125) );
  NAND3BX4 U271 ( .AN(n156), .B(n158), .C(n142), .Y(n127) );
  NAND2X4 U272 ( .A(n164), .B(n165), .Y(n143) );
  NOR3BX4 U273 ( .AN(n163), .B(n146), .C(n145), .Y(n156) );
  XOR2X4 U274 ( .A(n169), .B(n170), .Y(SUM[23]) );
  OR2X4 U275 ( .A(A[23]), .B(B[23]), .Y(n163) );
  OR2X4 U276 ( .A(A[22]), .B(B[22]), .Y(n144) );
  OAI2BB1X4 U277 ( .A0N(n166), .A1N(n174), .B0(n175), .Y(n172) );
  OR2X4 U278 ( .A(A[21]), .B(B[21]), .Y(n166) );
  NAND2X4 U279 ( .A(n146), .B(n178), .Y(n174) );
  NAND2X4 U280 ( .A(n179), .B(n180), .Y(n146) );
  CLKINVX3 U281 ( .A(n180), .Y(n182) );
  OR2X4 U282 ( .A(A[20]), .B(B[20]), .Y(n180) );
  NAND3X4 U283 ( .A(n184), .B(n183), .C(n185), .Y(n179) );
  AOI21X4 U284 ( .A0(n186), .A1(n187), .B0(n188), .Y(n185) );
  NOR2X4 U285 ( .A(n190), .B(n191), .Y(n187) );
  AOI21X4 U286 ( .A0(n194), .A1(n207), .B0(n208), .Y(n206) );
  OR2X4 U287 ( .A(A[19]), .B(B[19]), .Y(n195) );
  XOR2X4 U288 ( .A(n207), .B(n209), .Y(SUM[18]) );
  OR2X4 U289 ( .A(B[18]), .B(A[18]), .Y(n194) );
  OAI21X4 U290 ( .A0(n210), .A1(n192), .B0(n202), .Y(n207) );
  NAND2X4 U291 ( .A(n213), .B(n193), .Y(n211) );
  OR2X4 U292 ( .A(A[16]), .B(B[16]), .Y(n197) );
  NOR2X4 U293 ( .A(n49), .B(n50), .Y(n236) );
  OAI21X4 U294 ( .A0(n241), .A1(n23), .B0(n223), .Y(n239) );
  OAI21X4 U295 ( .A0(n244), .A1(n245), .B0(n222), .Y(n242) );
  OAI21X4 U296 ( .A0(n248), .A1(n225), .B0(n230), .Y(n246) );
  NAND4BBX4 U297 ( .AN(n59), .BN(n55), .C(n252), .D(n251), .Y(n225) );
  CLKINVX3 U298 ( .A(n56), .Y(n248) );
  XOR2X4 U299 ( .A(n259), .B(n260), .Y(SUM[11]) );
  AOI21X4 U300 ( .A0(n252), .A1(n261), .B0(n262), .Y(n260) );
  OR2X4 U301 ( .A(A[10]), .B(B[10]), .Y(n252) );
  OR2X4 U302 ( .A(A[9]), .B(B[9]), .Y(n253) );
  OAI21X4 U303 ( .A0(n72), .A1(n234), .B0(n233), .Y(n56) );
  NAND2BX4 U304 ( .AN(n63), .B(n265), .Y(n233) );
  NAND3BX4 U305 ( .AN(n44), .B(n267), .C(n68), .Y(n266) );
  OR2X4 U306 ( .A(A[6]), .B(B[6]), .Y(n68) );
endmodule


module hash_core_DW01_add_46 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n234, n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233;

  OAI21X1 U2 ( .A0(n184), .A1(n182), .B0(n185), .Y(n167) );
  NAND2X1 U3 ( .A(B[13]), .B(A[13]), .Y(n191) );
  OAI21X1 U4 ( .A0(n105), .A1(n95), .B0(n94), .Y(n103) );
  NAND2X2 U5 ( .A(n1), .B(n2), .Y(n3) );
  NAND2X4 U6 ( .A(n3), .B(n45), .Y(n40) );
  CLKINVX1 U7 ( .A(n43), .Y(n1) );
  INVX12 U8 ( .A(n44), .Y(n2) );
  NAND2XL U9 ( .A(n50), .B(n51), .Y(n44) );
  AOI2BB1X4 U10 ( .A0N(n46), .A1N(n47), .B0(n48), .Y(n45) );
  NAND2X2 U11 ( .A(n176), .B(n175), .Y(n4) );
  NAND2X4 U12 ( .A(n5), .B(n177), .Y(n168) );
  CLKINVX3 U13 ( .A(n4), .Y(n5) );
  NAND3BX4 U14 ( .AN(n167), .B(n169), .C(n168), .Y(n143) );
  OAI21X2 U15 ( .A0(n22), .A1(n154), .B0(n155), .Y(n153) );
  NOR2X2 U16 ( .A(A[17]), .B(B[17]), .Y(n22) );
  XOR2X2 U17 ( .A(n67), .B(n78), .Y(SUM[2]) );
  BUFX4 U18 ( .A(n234), .Y(SUM[14]) );
  OAI21X4 U19 ( .A0(n163), .A1(n22), .B0(n155), .Y(n161) );
  AOI21X2 U20 ( .A0(n28), .A1(n212), .B0(n217), .Y(n219) );
  OAI2BB1X2 U21 ( .A0N(n220), .A1N(n36), .B0(n221), .Y(n28) );
  INVX4 U22 ( .A(n67), .Y(n65) );
  XOR2X4 U23 ( .A(n40), .B(n41), .Y(SUM[7]) );
  AOI2BB2X2 U24 ( .B0(n170), .B1(n38), .A0N(n171), .A1N(n172), .Y(n169) );
  NOR2X2 U25 ( .A(n172), .B(n174), .Y(n175) );
  NOR2X2 U26 ( .A(n174), .B(n172), .Y(n170) );
  NAND2X2 U27 ( .A(n180), .B(n181), .Y(n172) );
  NOR2BXL U28 ( .AN(n34), .B(n35), .Y(n33) );
  NAND2X4 U29 ( .A(n30), .B(n34), .Y(n206) );
  NAND2X2 U30 ( .A(B[8]), .B(A[8]), .Y(n34) );
  NAND2X2 U31 ( .A(B[11]), .B(A[11]), .Y(n204) );
  NOR2X4 U32 ( .A(A[11]), .B(B[11]), .Y(n21) );
  NOR2X2 U33 ( .A(n31), .B(n209), .Y(n205) );
  NOR2X4 U34 ( .A(n35), .B(n31), .Y(n211) );
  INVX8 U35 ( .A(n212), .Y(n31) );
  NOR2X1 U36 ( .A(A[0]), .B(B[0]), .Y(n15) );
  NAND2X4 U37 ( .A(B[0]), .B(A[0]), .Y(n158) );
  NAND2X2 U38 ( .A(n210), .B(n211), .Y(n174) );
  INVX1 U39 ( .A(n24), .Y(n13) );
  INVX1 U40 ( .A(n127), .Y(n119) );
  INVXL U41 ( .A(n23), .Y(n8) );
  INVXL U42 ( .A(n130), .Y(n9) );
  INVXL U43 ( .A(n17), .Y(n12) );
  CLKINVX2 U44 ( .A(n158), .Y(n80) );
  NAND2X2 U45 ( .A(n10), .B(n50), .Y(n11) );
  OAI21XL U46 ( .A0(n23), .A1(n129), .B0(n130), .Y(n128) );
  CLKINVX3 U47 ( .A(n50), .Y(n54) );
  NOR2X1 U48 ( .A(A[21]), .B(B[21]), .Y(n23) );
  NAND2X1 U49 ( .A(B[16]), .B(A[16]), .Y(n154) );
  NAND2X1 U50 ( .A(B[12]), .B(A[12]), .Y(n190) );
  NOR2X2 U51 ( .A(A[12]), .B(B[12]), .Y(n19) );
  OR2X2 U52 ( .A(A[10]), .B(B[10]), .Y(n216) );
  NAND2X1 U53 ( .A(B[4]), .B(A[4]), .Y(n57) );
  NAND2X1 U54 ( .A(n83), .B(n84), .Y(n77) );
  INVX1 U55 ( .A(n7), .Y(n133) );
  XNOR2X2 U56 ( .A(n14), .B(n192), .Y(SUM[15]) );
  XOR2X1 U57 ( .A(n193), .B(n195), .Y(n234) );
  CLKINVX3 U58 ( .A(n216), .Y(n209) );
  NOR2X1 U59 ( .A(n39), .B(n35), .Y(n220) );
  OR2X2 U60 ( .A(A[9]), .B(B[9]), .Y(n212) );
  NOR2BX1 U61 ( .AN(n42), .B(n18), .Y(n41) );
  NOR2BX1 U62 ( .AN(n63), .B(n64), .Y(n62) );
  NOR2BX1 U63 ( .AN(n81), .B(n157), .Y(n156) );
  NOR2X2 U64 ( .A(n54), .B(n60), .Y(n232) );
  CLKINVX3 U65 ( .A(n55), .Y(n60) );
  CLKINVX3 U66 ( .A(n43), .Y(n10) );
  XOR2X2 U67 ( .A(n58), .B(n43), .Y(SUM[5]) );
  NAND2X2 U68 ( .A(n232), .B(n233), .Y(n39) );
  XOR2X2 U69 ( .A(n159), .B(n160), .Y(SUM[19]) );
  OAI2BB1X4 U70 ( .A0N(n196), .A1N(n12), .B0(n191), .Y(n193) );
  OAI2BB1X4 U71 ( .A0N(n16), .A1N(n198), .B0(n190), .Y(n196) );
  AOI21X1 U72 ( .A0(n187), .A1(n193), .B0(n189), .Y(n192) );
  NAND2BX4 U73 ( .AN(n66), .B(n231), .Y(n178) );
  CLKINVX3 U74 ( .A(n222), .Y(n35) );
  AOI21X1 U75 ( .A0(n28), .A1(n212), .B0(n217), .Y(n215) );
  XOR2X2 U76 ( .A(n196), .B(n197), .Y(SUM[13]) );
  AOI21X4 U77 ( .A0(n36), .A1(n55), .B0(n56), .Y(n43) );
  OR2X4 U78 ( .A(A[8]), .B(B[8]), .Y(n222) );
  NAND2X2 U79 ( .A(B[7]), .B(A[7]), .Y(n42) );
  AOI21X4 U80 ( .A0(n135), .A1(n8), .B0(n9), .Y(n7) );
  OAI21X4 U81 ( .A0(n25), .A1(n137), .B0(n129), .Y(n135) );
  OR2X4 U82 ( .A(A[14]), .B(B[14]), .Y(n187) );
  NAND2X4 U83 ( .A(n11), .B(n47), .Y(n52) );
  NAND2X4 U84 ( .A(B[2]), .B(A[2]), .Y(n66) );
  OAI2BB1X1 U85 ( .A0N(n13), .A1N(n143), .B0(n154), .Y(n164) );
  NAND2X4 U86 ( .A(B[5]), .B(A[5]), .Y(n47) );
  NOR2X4 U87 ( .A(A[7]), .B(B[7]), .Y(n18) );
  NAND2XL U88 ( .A(B[17]), .B(A[17]), .Y(n155) );
  NAND2XL U89 ( .A(B[21]), .B(A[21]), .Y(n130) );
  XOR2X2 U90 ( .A(n28), .B(n29), .Y(SUM[9]) );
  OAI21X1 U91 ( .A0(n65), .A1(n20), .B0(n66), .Y(n61) );
  OAI2BB1X4 U92 ( .A0N(n79), .A1N(n80), .B0(n81), .Y(n67) );
  NAND2X2 U93 ( .A(B[3]), .B(A[3]), .Y(n63) );
  NAND2XL U94 ( .A(B[14]), .B(A[14]), .Y(n194) );
  NOR2X1 U95 ( .A(n144), .B(n145), .Y(n141) );
  OAI21X2 U96 ( .A0(n215), .A1(n209), .B0(n208), .Y(n213) );
  NAND2X4 U97 ( .A(n139), .B(n140), .Y(n118) );
  AOI21X2 U98 ( .A0(n47), .A1(n57), .B0(n54), .Y(n224) );
  NAND2X2 U99 ( .A(n89), .B(n98), .Y(n108) );
  NOR2BXL U100 ( .AN(n57), .B(n60), .Y(n59) );
  NOR2BXL U101 ( .AN(n30), .B(n31), .Y(n29) );
  NAND2X1 U102 ( .A(n152), .B(n153), .Y(n150) );
  NOR2BX1 U103 ( .AN(n154), .B(n24), .Y(n166) );
  INVX1 U104 ( .A(n152), .Y(n144) );
  NOR2X4 U105 ( .A(A[2]), .B(B[2]), .Y(n20) );
  NOR2X1 U106 ( .A(A[20]), .B(B[20]), .Y(n25) );
  NOR2XL U107 ( .A(n174), .B(n39), .Y(n200) );
  AOI21XL U108 ( .A0(n202), .A1(n38), .B0(n173), .Y(n201) );
  INVXL U109 ( .A(n174), .Y(n202) );
  INVX1 U110 ( .A(n173), .Y(n171) );
  XOR2X2 U111 ( .A(n36), .B(n59), .Y(SUM[4]) );
  AND2X1 U112 ( .A(n185), .B(n186), .Y(n14) );
  CLKINVX4 U113 ( .A(n208), .Y(n207) );
  NOR2X1 U114 ( .A(n18), .B(n46), .Y(n233) );
  NAND2X2 U115 ( .A(n110), .B(n111), .Y(n89) );
  NAND3X2 U116 ( .A(n141), .B(n142), .C(n143), .Y(n140) );
  INVX1 U117 ( .A(n19), .Y(n16) );
  AOI2BB1X2 U118 ( .A0N(n18), .A1N(n49), .B0(n227), .Y(n226) );
  NOR2X1 U119 ( .A(n209), .B(n21), .Y(n210) );
  NOR2BX1 U120 ( .AN(n100), .B(n92), .Y(n91) );
  INVX8 U121 ( .A(n51), .Y(n46) );
  NOR2BXL U122 ( .AN(n99), .B(n97), .Y(n109) );
  AOI21XL U123 ( .A0(n38), .A1(n222), .B0(n223), .Y(n221) );
  NOR2BXL U124 ( .AN(n194), .B(n183), .Y(n195) );
  NOR2BXL U125 ( .AN(n49), .B(n46), .Y(n53) );
  NAND2XL U126 ( .A(n71), .B(n72), .Y(n70) );
  OR2X4 U127 ( .A(A[4]), .B(B[4]), .Y(n55) );
  OR2X4 U128 ( .A(A[5]), .B(B[5]), .Y(n50) );
  NOR2BX1 U129 ( .AN(n158), .B(n15), .Y(SUM[0]) );
  NOR2X2 U130 ( .A(A[13]), .B(B[13]), .Y(n17) );
  NAND2X1 U131 ( .A(B[9]), .B(A[9]), .Y(n30) );
  NAND2XL U132 ( .A(B[6]), .B(A[6]), .Y(n49) );
  NAND2XL U133 ( .A(B[15]), .B(A[15]), .Y(n185) );
  NAND2XL U134 ( .A(B[18]), .B(A[18]), .Y(n151) );
  NAND2XL U135 ( .A(B[19]), .B(A[19]), .Y(n149) );
  NAND2XL U136 ( .A(B[22]), .B(A[22]), .Y(n126) );
  NAND2XL U137 ( .A(B[23]), .B(A[23]), .Y(n124) );
  OR2XL U138 ( .A(A[24]), .B(B[24]), .Y(n111) );
  OAI2BB1X1 U139 ( .A0N(n200), .A1N(n36), .B0(n201), .Y(n198) );
  INVXL U140 ( .A(n38), .Y(n37) );
  INVX1 U141 ( .A(n39), .Y(n177) );
  NOR2X1 U142 ( .A(n119), .B(n120), .Y(n116) );
  INVX1 U143 ( .A(n178), .Y(n228) );
  NOR2BX1 U144 ( .AN(n191), .B(n17), .Y(n197) );
  NOR2BX1 U145 ( .AN(n204), .B(n21), .Y(n214) );
  NOR2X1 U146 ( .A(n18), .B(n46), .Y(n225) );
  INVX1 U147 ( .A(n57), .Y(n56) );
  INVX1 U148 ( .A(n118), .Y(n137) );
  INVX1 U149 ( .A(n164), .Y(n163) );
  XOR2X2 U150 ( .A(n61), .B(n62), .Y(SUM[3]) );
  XOR2X1 U151 ( .A(n131), .B(n132), .Y(SUM[23]) );
  NOR2BX1 U152 ( .AN(n124), .B(n120), .Y(n132) );
  OAI21XL U153 ( .A0(n7), .A1(n119), .B0(n126), .Y(n131) );
  XOR2X1 U154 ( .A(n133), .B(n134), .Y(SUM[22]) );
  NOR2BX1 U155 ( .AN(n126), .B(n119), .Y(n134) );
  INVX1 U156 ( .A(n34), .Y(n223) );
  NOR2X1 U157 ( .A(n182), .B(n183), .Y(n181) );
  NOR2X1 U158 ( .A(n17), .B(n19), .Y(n180) );
  AOI21X1 U159 ( .A0(n146), .A1(n147), .B0(n148), .Y(n139) );
  INVX1 U160 ( .A(n149), .Y(n148) );
  XOR2X2 U161 ( .A(n218), .B(n219), .Y(SUM[10]) );
  NAND2X1 U162 ( .A(n208), .B(n216), .Y(n218) );
  XOR2X1 U163 ( .A(n161), .B(n162), .Y(SUM[18]) );
  NOR2BX1 U164 ( .AN(n151), .B(n144), .Y(n162) );
  INVX1 U165 ( .A(n186), .Y(n182) );
  INVX1 U166 ( .A(n187), .Y(n183) );
  AOI21X1 U167 ( .A0(n187), .A1(n188), .B0(n189), .Y(n184) );
  OAI21XL U168 ( .A0(n17), .A1(n190), .B0(n191), .Y(n188) );
  XOR2X1 U169 ( .A(n143), .B(n166), .Y(SUM[16]) );
  XOR2X1 U170 ( .A(n164), .B(n165), .Y(SUM[17]) );
  NOR2BX1 U171 ( .AN(n155), .B(n22), .Y(n165) );
  XOR2X1 U172 ( .A(n135), .B(n136), .Y(SUM[21]) );
  NOR2BX1 U173 ( .AN(n130), .B(n23), .Y(n136) );
  XOR2X1 U174 ( .A(n103), .B(n104), .Y(SUM[27]) );
  NOR2BX1 U175 ( .AN(n100), .B(n26), .Y(n104) );
  INVX1 U176 ( .A(n106), .Y(n105) );
  NAND2X1 U177 ( .A(n50), .B(n47), .Y(n58) );
  XOR2X2 U178 ( .A(n32), .B(n33), .Y(SUM[8]) );
  OAI2BB1X1 U179 ( .A0N(n177), .A1N(n36), .B0(n37), .Y(n32) );
  XOR2X1 U180 ( .A(n198), .B(n199), .Y(SUM[12]) );
  NOR2BX1 U181 ( .AN(n190), .B(n19), .Y(n199) );
  XOR2X1 U182 ( .A(n80), .B(n156), .Y(SUM[1]) );
  NOR2BX1 U183 ( .AN(n66), .B(n20), .Y(n78) );
  NOR2BX1 U184 ( .AN(n149), .B(n145), .Y(n160) );
  OAI2BB1X1 U185 ( .A0N(n152), .A1N(n161), .B0(n151), .Y(n159) );
  NAND2X1 U186 ( .A(n114), .B(n115), .Y(n110) );
  AOI21X1 U187 ( .A0(n121), .A1(n122), .B0(n123), .Y(n114) );
  NAND3X1 U188 ( .A(n116), .B(n117), .C(n118), .Y(n115) );
  INVX1 U189 ( .A(n124), .Y(n123) );
  OAI2BB1X1 U190 ( .A0N(n102), .A1N(n108), .B0(n99), .Y(n106) );
  NAND3XL U191 ( .A(n63), .B(n178), .C(n179), .Y(n176) );
  INVX1 U192 ( .A(n49), .Y(n48) );
  INVX1 U193 ( .A(n42), .Y(n227) );
  OAI21XL U194 ( .A0(n27), .A1(n75), .B0(n76), .Y(n71) );
  INVX1 U195 ( .A(n77), .Y(n75) );
  OAI21XL U196 ( .A0(n89), .A1(n90), .B0(n91), .Y(n85) );
  NAND3BX1 U197 ( .AN(n26), .B(n101), .C(n102), .Y(n90) );
  XOR2X1 U198 ( .A(n106), .B(n107), .Y(SUM[26]) );
  NOR2BX1 U199 ( .AN(n94), .B(n95), .Y(n107) );
  NAND2X1 U200 ( .A(n125), .B(n126), .Y(n121) );
  NAND2X1 U201 ( .A(n127), .B(n128), .Y(n125) );
  INVX1 U202 ( .A(n30), .Y(n217) );
  INVX1 U203 ( .A(n147), .Y(n145) );
  INVX1 U204 ( .A(n194), .Y(n189) );
  XOR2X1 U205 ( .A(n71), .B(n73), .Y(SUM[30]) );
  NOR2BX1 U206 ( .AN(n69), .B(n74), .Y(n73) );
  INVX1 U207 ( .A(n72), .Y(n74) );
  XOR2X1 U208 ( .A(n85), .B(n87), .Y(SUM[28]) );
  NOR2BX1 U209 ( .AN(n84), .B(n88), .Y(n87) );
  INVX1 U210 ( .A(n86), .Y(n88) );
  XOR2X1 U211 ( .A(n118), .B(n138), .Y(SUM[20]) );
  NOR2BX1 U212 ( .AN(n129), .B(n25), .Y(n138) );
  XOR2X1 U213 ( .A(n110), .B(n112), .Y(SUM[24]) );
  NOR2BX1 U214 ( .AN(n98), .B(n113), .Y(n112) );
  INVX1 U215 ( .A(n111), .Y(n113) );
  XOR2X1 U216 ( .A(n77), .B(n82), .Y(SUM[29]) );
  NOR2BX1 U217 ( .AN(n76), .B(n27), .Y(n82) );
  XOR2X1 U218 ( .A(n108), .B(n109), .Y(SUM[25]) );
  NOR2X1 U219 ( .A(n22), .B(n24), .Y(n142) );
  NAND2X1 U220 ( .A(n85), .B(n86), .Y(n83) );
  NAND2X1 U221 ( .A(n150), .B(n151), .Y(n146) );
  INVX1 U222 ( .A(n122), .Y(n120) );
  NOR2X1 U223 ( .A(n23), .B(n25), .Y(n117) );
  NAND2X1 U224 ( .A(n69), .B(n70), .Y(n68) );
  INVX1 U225 ( .A(n101), .Y(n95) );
  INVX1 U226 ( .A(n102), .Y(n97) );
  AOI21X1 U227 ( .A0(n93), .A1(n94), .B0(n26), .Y(n92) );
  NAND2BX1 U228 ( .AN(n95), .B(n96), .Y(n93) );
  OAI21XL U229 ( .A0(n97), .A1(n98), .B0(n99), .Y(n96) );
  XOR3X2 U230 ( .A(B[31]), .B(A[31]), .C(n68), .Y(SUM[31]) );
  NAND2X1 U231 ( .A(B[10]), .B(A[10]), .Y(n208) );
  NAND2X2 U232 ( .A(B[1]), .B(A[1]), .Y(n81) );
  OR2X2 U233 ( .A(A[15]), .B(B[15]), .Y(n186) );
  NOR2X1 U234 ( .A(A[16]), .B(B[16]), .Y(n24) );
  OR2X2 U235 ( .A(A[18]), .B(B[18]), .Y(n152) );
  OR2X2 U236 ( .A(A[19]), .B(B[19]), .Y(n147) );
  NAND2X1 U237 ( .A(B[20]), .B(A[20]), .Y(n129) );
  OR2X2 U238 ( .A(A[23]), .B(B[23]), .Y(n122) );
  OR2X2 U239 ( .A(A[22]), .B(B[22]), .Y(n127) );
  NOR2X1 U240 ( .A(A[27]), .B(B[27]), .Y(n26) );
  NAND2X1 U241 ( .A(B[24]), .B(A[24]), .Y(n98) );
  NAND2X1 U242 ( .A(B[26]), .B(A[26]), .Y(n94) );
  NAND2X1 U243 ( .A(B[25]), .B(A[25]), .Y(n99) );
  OR2X2 U244 ( .A(A[25]), .B(B[25]), .Y(n102) );
  NAND2X1 U245 ( .A(B[27]), .B(A[27]), .Y(n100) );
  OR2X2 U246 ( .A(A[28]), .B(B[28]), .Y(n86) );
  NOR2X1 U247 ( .A(A[29]), .B(B[29]), .Y(n27) );
  OR2X2 U248 ( .A(A[26]), .B(B[26]), .Y(n101) );
  NAND2X1 U249 ( .A(B[30]), .B(A[30]), .Y(n69) );
  NAND2X1 U250 ( .A(B[28]), .B(A[28]), .Y(n84) );
  OR2X2 U251 ( .A(A[30]), .B(B[30]), .Y(n72) );
  NAND3BX4 U252 ( .AN(n228), .B(n63), .C(n179), .Y(n36) );
  NAND2X1 U253 ( .A(B[29]), .B(A[29]), .Y(n76) );
  XOR2X4 U254 ( .A(n52), .B(n53), .Y(SUM[6]) );
  OAI21X4 U255 ( .A0(n203), .A1(n21), .B0(n204), .Y(n173) );
  AOI21X4 U256 ( .A0(n205), .A1(n206), .B0(n207), .Y(n203) );
  XOR2X4 U257 ( .A(n213), .B(n214), .Y(SUM[11]) );
  OAI2BB1X4 U258 ( .A0N(n224), .A1N(n225), .B0(n226), .Y(n38) );
  NAND2X4 U259 ( .A(n229), .B(n230), .Y(n179) );
  NOR2X4 U260 ( .A(n64), .B(n20), .Y(n230) );
  CLKINVX3 U261 ( .A(n231), .Y(n64) );
  AOI21X4 U262 ( .A0(n81), .A1(n158), .B0(n157), .Y(n229) );
  CLKINVX3 U263 ( .A(n79), .Y(n157) );
  OR2X4 U264 ( .A(A[1]), .B(B[1]), .Y(n79) );
  OR2X4 U265 ( .A(A[3]), .B(B[3]), .Y(n231) );
  OR2X4 U266 ( .A(A[6]), .B(B[6]), .Y(n51) );
endmodule


module hash_core_DW01_add_50 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273;

  NOR2X2 U2 ( .A(n49), .B(n41), .Y(n250) );
  NOR2X2 U3 ( .A(n41), .B(n248), .Y(n242) );
  CLKINVX3 U4 ( .A(n215), .Y(n213) );
  INVX2 U5 ( .A(n251), .Y(n41) );
  OR2X4 U6 ( .A(A[0]), .B(B[0]), .Y(n34) );
  AND2X2 U7 ( .A(n56), .B(n55), .Y(n1) );
  AND2X4 U8 ( .A(n57), .B(n1), .Y(n27) );
  OR2X2 U9 ( .A(n58), .B(n61), .Y(n56) );
  NAND2XL U10 ( .A(n125), .B(n3), .Y(n4) );
  NAND2X2 U11 ( .A(n2), .B(n31), .Y(n5) );
  NAND2X2 U12 ( .A(n4), .B(n5), .Y(SUM[26]) );
  INVX1 U13 ( .A(n125), .Y(n2) );
  INVX1 U14 ( .A(n31), .Y(n3) );
  NAND2X4 U15 ( .A(n127), .B(n122), .Y(n125) );
  XOR2X2 U16 ( .A(n123), .B(n124), .Y(SUM[27]) );
  CLKINVX1 U17 ( .A(n102), .Y(n173) );
  AND2X1 U18 ( .A(n102), .B(n34), .Y(SUM[0]) );
  CLKINVX8 U19 ( .A(n102), .Y(n88) );
  NAND2X4 U20 ( .A(B[0]), .B(A[0]), .Y(n102) );
  AOI21X4 U21 ( .A0(n199), .A1(n200), .B0(n201), .Y(n188) );
  NOR2X2 U22 ( .A(n194), .B(n193), .Y(n199) );
  OAI21X4 U23 ( .A0(n260), .A1(n259), .B0(n261), .Y(n256) );
  INVX2 U24 ( .A(n45), .Y(n260) );
  INVX4 U25 ( .A(n51), .Y(n231) );
  AOI21X2 U26 ( .A0(n50), .A1(n60), .B0(n45), .Y(n264) );
  NAND2X4 U27 ( .A(n11), .B(n12), .Y(n13) );
  INVX4 U28 ( .A(n194), .Y(n12) );
  CLKINVX2 U29 ( .A(n45), .Y(n252) );
  OAI2BB1X4 U30 ( .A0N(n242), .A1N(n243), .B0(n244), .Y(n238) );
  OAI21X4 U31 ( .A0(n42), .A1(n43), .B0(n44), .Y(n38) );
  AOI21X2 U32 ( .A0(n45), .A1(n46), .B0(n47), .Y(n44) );
  NAND2BX4 U33 ( .AN(n220), .B(n12), .Y(n232) );
  NAND2X4 U34 ( .A(n16), .B(n17), .Y(SUM[16]) );
  BUFX4 U35 ( .A(n245), .Y(n6) );
  BUFX4 U36 ( .A(n40), .Y(n7) );
  XOR2X4 U37 ( .A(n181), .B(n182), .Y(SUM[17]) );
  NOR2BX1 U38 ( .AN(n7), .B(n41), .Y(n39) );
  NAND2X2 U39 ( .A(n7), .B(n48), .Y(n243) );
  NOR2BX4 U40 ( .AN(n6), .B(n246), .Y(n244) );
  NAND2X2 U41 ( .A(n213), .B(n214), .Y(n187) );
  INVX1 U42 ( .A(n155), .Y(n29) );
  NOR2BXL U43 ( .AN(n144), .B(n142), .Y(n155) );
  NAND2X2 U44 ( .A(n10), .B(n261), .Y(n262) );
  NOR2BX1 U45 ( .AN(n48), .B(n49), .Y(n52) );
  NOR2X2 U46 ( .A(n203), .B(n218), .Y(n217) );
  INVX1 U47 ( .A(n247), .Y(n246) );
  AOI21X2 U48 ( .A0(n205), .A1(n206), .B0(n207), .Y(n202) );
  INVX1 U49 ( .A(n77), .Y(n196) );
  OAI21XL U50 ( .A0(n142), .A1(n143), .B0(n144), .Y(n141) );
  NOR2X2 U51 ( .A(n248), .B(n241), .Y(n249) );
  INVX1 U52 ( .A(n236), .Y(n241) );
  INVX4 U53 ( .A(n63), .Y(n66) );
  INVX2 U54 ( .A(n198), .Y(n74) );
  INVX4 U55 ( .A(n62), .Y(n72) );
  CLKINVX3 U56 ( .A(n90), .Y(n89) );
  NAND3BX1 U57 ( .AN(n35), .B(n171), .C(n172), .Y(n160) );
  INVX1 U58 ( .A(n170), .Y(n161) );
  NOR2X1 U59 ( .A(A[23]), .B(B[23]), .Y(n36) );
  NAND2X2 U60 ( .A(n153), .B(n144), .Y(n151) );
  INVX1 U61 ( .A(n146), .Y(n140) );
  NAND2BX2 U62 ( .AN(n241), .B(n238), .Y(n215) );
  OAI2BB1X1 U63 ( .A0N(n7), .A1N(n48), .B0(n251), .Y(n261) );
  NAND2X1 U64 ( .A(n251), .B(n46), .Y(n259) );
  NAND2X1 U65 ( .A(B[8]), .B(A[8]), .Y(n48) );
  NOR2X1 U66 ( .A(n72), .B(n73), .Y(n71) );
  NAND2X2 U67 ( .A(B[2]), .B(A[2]), .Y(n85) );
  CLKINVX3 U68 ( .A(n89), .Y(n9) );
  INVX1 U69 ( .A(n180), .Y(n30) );
  NAND2X1 U70 ( .A(n14), .B(n185), .Y(n17) );
  NAND2X1 U71 ( .A(n204), .B(n219), .Y(n221) );
  AOI21X2 U72 ( .A0(n228), .A1(n224), .B0(n229), .Y(n227) );
  OR2X2 U73 ( .A(A[11]), .B(B[11]), .Y(n236) );
  INVX1 U74 ( .A(n48), .Y(n47) );
  NAND2X2 U75 ( .A(n37), .B(n59), .Y(n79) );
  XOR2X1 U76 ( .A(n94), .B(n33), .Y(SUM[30]) );
  NAND2X2 U77 ( .A(n101), .B(n9), .Y(n100) );
  OAI21X1 U78 ( .A0(n209), .A1(n210), .B0(n211), .Y(n206) );
  NOR2BX1 U79 ( .AN(n211), .B(n209), .Y(n230) );
  NOR2X2 U80 ( .A(n209), .B(n220), .Y(n216) );
  INVX2 U81 ( .A(n228), .Y(n209) );
  OAI21X4 U82 ( .A0(n178), .A1(n165), .B0(n164), .Y(n176) );
  CLKINVX2 U83 ( .A(n231), .Y(n11) );
  INVX1 U84 ( .A(n86), .Y(n84) );
  INVXL U85 ( .A(n271), .Y(n8) );
  XOR2X2 U86 ( .A(n37), .B(n28), .Y(SUM[4]) );
  NOR3X2 U87 ( .A(n192), .B(n193), .C(n194), .Y(n191) );
  INVX1 U88 ( .A(n208), .Y(n207) );
  NAND2X1 U89 ( .A(n208), .B(n205), .Y(n226) );
  INVX1 U90 ( .A(n87), .Y(n175) );
  NAND2XL U91 ( .A(n212), .B(n54), .Y(n200) );
  NAND2BX2 U92 ( .AN(n165), .B(n166), .Y(n163) );
  NOR2BX1 U93 ( .AN(n164), .B(n165), .Y(n180) );
  OR2X4 U94 ( .A(n264), .B(n259), .Y(n10) );
  NAND2X4 U95 ( .A(n13), .B(n215), .Y(n239) );
  NAND2XL U96 ( .A(n183), .B(n15), .Y(n16) );
  INVXL U97 ( .A(n183), .Y(n14) );
  INVXL U98 ( .A(n185), .Y(n15) );
  NOR2BX2 U99 ( .AN(n168), .B(n186), .Y(n185) );
  NAND2X2 U100 ( .A(B[6]), .B(A[6]), .Y(n64) );
  INVX4 U101 ( .A(n60), .Y(n42) );
  NAND3BX1 U102 ( .AN(n58), .B(n59), .C(n60), .Y(n57) );
  NAND2BX2 U103 ( .AN(n49), .B(n50), .Y(n43) );
  CLKINVX4 U104 ( .A(n192), .Y(n50) );
  XOR2X2 U105 ( .A(n128), .B(n129), .Y(SUM[25]) );
  OAI2BB1X4 U106 ( .A0N(B[0]), .A1N(A[0]), .B0(n90), .Y(n198) );
  OAI21X2 U107 ( .A0(n70), .A1(n69), .B0(n71), .Y(n68) );
  OAI21X1 U108 ( .A0(n74), .A1(n75), .B0(n76), .Y(n70) );
  OAI21X4 U109 ( .A0(n83), .A1(n84), .B0(n85), .Y(n80) );
  AOI21X2 U110 ( .A0(n87), .A1(n88), .B0(n89), .Y(n83) );
  OAI21XL U111 ( .A0(n218), .A1(n211), .B0(n208), .Y(n225) );
  INVX1 U112 ( .A(n211), .Y(n229) );
  NAND2X2 U113 ( .A(B[13]), .B(A[13]), .Y(n211) );
  NAND2X4 U114 ( .A(n130), .B(n131), .Y(n110) );
  OAI21X4 U115 ( .A0(n134), .A1(n135), .B0(n136), .Y(n130) );
  NAND3BX4 U116 ( .AN(n197), .B(n77), .C(n269), .Y(n37) );
  INVX2 U117 ( .A(n151), .Y(n150) );
  OAI21XL U118 ( .A0(n74), .A1(n8), .B0(n195), .Y(n190) );
  NOR2XL U119 ( .A(n196), .B(n197), .Y(n195) );
  CLKINVX2 U120 ( .A(n179), .Y(n178) );
  OAI21X4 U121 ( .A0(n159), .A1(n160), .B0(n21), .Y(n20) );
  XOR2XL U122 ( .A(n103), .B(n97), .Y(SUM[29]) );
  NOR2BXL U123 ( .AN(n170), .B(n35), .Y(n177) );
  NAND2X2 U124 ( .A(B[16]), .B(A[16]), .Y(n168) );
  NAND2X1 U125 ( .A(B[21]), .B(A[21]), .Y(n144) );
  OR2XL U126 ( .A(A[16]), .B(B[16]), .Y(n184) );
  AND2X2 U127 ( .A(n86), .B(n85), .Y(n19) );
  NAND2X2 U128 ( .A(n79), .B(n61), .Y(n78) );
  NAND3BXL U129 ( .AN(n36), .B(n146), .C(n147), .Y(n135) );
  AOI21X1 U130 ( .A0(n113), .A1(n125), .B0(n126), .Y(n124) );
  NOR2BX1 U131 ( .AN(n210), .B(n220), .Y(n240) );
  NOR2BXL U132 ( .AN(n145), .B(n36), .Y(n149) );
  NAND3XL U133 ( .A(n34), .B(n88), .C(n87), .Y(n101) );
  NOR2X1 U134 ( .A(A[19]), .B(B[19]), .Y(n35) );
  NAND2XL U135 ( .A(B[18]), .B(A[18]), .Y(n164) );
  NAND2X1 U136 ( .A(B[17]), .B(A[17]), .Y(n169) );
  NAND2X1 U137 ( .A(B[24]), .B(A[24]), .Y(n121) );
  NAND2X1 U138 ( .A(B[25]), .B(A[25]), .Y(n122) );
  OR2X2 U139 ( .A(A[25]), .B(B[25]), .Y(n111) );
  INVXL U140 ( .A(n193), .Y(n214) );
  NAND2X2 U141 ( .A(n190), .B(n191), .Y(n189) );
  AOI2BB1X4 U142 ( .A0N(n233), .A1N(n234), .B0(n235), .Y(n18) );
  NOR2BX4 U143 ( .AN(n9), .B(n175), .Y(n174) );
  INVX1 U144 ( .A(n270), .Y(n82) );
  XOR2X4 U145 ( .A(n100), .B(n19), .Y(SUM[2]) );
  NOR2BX1 U146 ( .AN(n145), .B(n137), .Y(n136) );
  INVXL U147 ( .A(n118), .Y(n126) );
  NOR2X2 U148 ( .A(n161), .B(n162), .Y(n21) );
  NAND2X2 U149 ( .A(n111), .B(n128), .Y(n127) );
  OAI21X1 U150 ( .A0(n167), .A1(n168), .B0(n169), .Y(n166) );
  INVXL U151 ( .A(n131), .Y(n133) );
  XNOR2X1 U152 ( .A(n104), .B(n22), .Y(SUM[28]) );
  NAND2X1 U153 ( .A(n107), .B(n105), .Y(n22) );
  AND2X1 U154 ( .A(n62), .B(n65), .Y(n23) );
  NOR2BXL U155 ( .AN(n169), .B(n167), .Y(n182) );
  XNOR2X4 U156 ( .A(n27), .B(n24), .Y(SUM[7]) );
  AND2X1 U157 ( .A(n53), .B(n54), .Y(n24) );
  NAND2XL U158 ( .A(n61), .B(n77), .Y(n69) );
  NOR2BXL U159 ( .AN(n139), .B(n140), .Y(n152) );
  AND2X1 U160 ( .A(n64), .B(n63), .Y(n25) );
  INVXL U161 ( .A(n210), .Y(n235) );
  INVXL U162 ( .A(n6), .Y(n254) );
  AND2X1 U163 ( .A(n247), .B(n236), .Y(n26) );
  NAND2XL U164 ( .A(n94), .B(n95), .Y(n93) );
  OR2X4 U165 ( .A(A[17]), .B(B[17]), .Y(n172) );
  OR2X4 U166 ( .A(A[18]), .B(B[18]), .Y(n171) );
  NAND2XL U167 ( .A(B[22]), .B(A[22]), .Y(n139) );
  NAND2X2 U168 ( .A(B[20]), .B(A[20]), .Y(n143) );
  NAND2XL U169 ( .A(B[19]), .B(A[19]), .Y(n170) );
  OR2X4 U170 ( .A(A[21]), .B(B[21]), .Y(n147) );
  NAND2XL U171 ( .A(B[23]), .B(A[23]), .Y(n145) );
  OR2XL U172 ( .A(A[20]), .B(B[20]), .Y(n156) );
  NOR2XL U173 ( .A(n209), .B(n218), .Y(n223) );
  INVXL U174 ( .A(n238), .Y(n233) );
  INVX1 U175 ( .A(n171), .Y(n165) );
  AND2X1 U176 ( .A(n61), .B(n59), .Y(n28) );
  INVX1 U177 ( .A(n172), .Y(n167) );
  XOR2X1 U178 ( .A(n130), .B(n132), .Y(SUM[24]) );
  NOR2BX1 U179 ( .AN(n121), .B(n133), .Y(n132) );
  XOR2X1 U180 ( .A(n20), .B(n157), .Y(SUM[20]) );
  NOR2BX1 U181 ( .AN(n143), .B(n158), .Y(n157) );
  INVX1 U182 ( .A(n156), .Y(n158) );
  INVX1 U183 ( .A(n184), .Y(n186) );
  NOR2BXL U184 ( .AN(n6), .B(n248), .Y(n263) );
  XNOR2X4 U185 ( .A(n154), .B(n29), .Y(SUM[21]) );
  NOR2BX1 U186 ( .AN(n122), .B(n120), .Y(n129) );
  NAND2X1 U187 ( .A(n116), .B(n112), .Y(n123) );
  XNOR2X4 U188 ( .A(n179), .B(n30), .Y(SUM[18]) );
  AND2X2 U189 ( .A(n118), .B(n113), .Y(n31) );
  NAND2X1 U190 ( .A(n110), .B(n121), .Y(n128) );
  AOI21X1 U191 ( .A0(n163), .A1(n164), .B0(n35), .Y(n162) );
  AND2X2 U192 ( .A(n64), .B(n32), .Y(n55) );
  OR2XL U193 ( .A(n65), .B(n66), .Y(n32) );
  NAND2XL U194 ( .A(n62), .B(n63), .Y(n58) );
  NAND2XL U195 ( .A(n236), .B(n237), .Y(n234) );
  AOI21X1 U196 ( .A0(n104), .A1(n105), .B0(n106), .Y(n97) );
  INVX1 U197 ( .A(n107), .Y(n106) );
  OAI21XL U198 ( .A0(n96), .A1(n97), .B0(n98), .Y(n94) );
  INVX1 U199 ( .A(n99), .Y(n96) );
  INVX1 U200 ( .A(n147), .Y(n142) );
  NAND2X1 U201 ( .A(n98), .B(n99), .Y(n103) );
  NAND2X1 U202 ( .A(n108), .B(n109), .Y(n104) );
  AOI21X1 U203 ( .A0(n114), .A1(n112), .B0(n115), .Y(n108) );
  NAND4BXL U204 ( .AN(n110), .B(n111), .C(n112), .D(n113), .Y(n109) );
  INVX1 U205 ( .A(n116), .Y(n115) );
  AOI21X1 U206 ( .A0(n138), .A1(n139), .B0(n36), .Y(n137) );
  NAND2BX1 U207 ( .AN(n140), .B(n141), .Y(n138) );
  AND2X2 U208 ( .A(n92), .B(n95), .Y(n33) );
  INVX1 U209 ( .A(n111), .Y(n120) );
  NAND2X1 U210 ( .A(n92), .B(n93), .Y(n91) );
  NAND2X1 U211 ( .A(n117), .B(n118), .Y(n114) );
  NAND2X1 U212 ( .A(n113), .B(n119), .Y(n117) );
  OAI21XL U213 ( .A0(n120), .A1(n121), .B0(n122), .Y(n119) );
  NAND2XL U214 ( .A(B[7]), .B(A[7]), .Y(n54) );
  NAND2XL U215 ( .A(B[14]), .B(A[14]), .Y(n208) );
  NAND2XL U216 ( .A(B[12]), .B(A[12]), .Y(n210) );
  NAND2XL U217 ( .A(B[9]), .B(A[9]), .Y(n40) );
  NAND2XL U218 ( .A(B[10]), .B(A[10]), .Y(n245) );
  NAND2XL U219 ( .A(B[15]), .B(A[15]), .Y(n204) );
  NAND2XL U220 ( .A(B[11]), .B(A[11]), .Y(n247) );
  XOR3X2 U221 ( .A(B[31]), .B(A[31]), .C(n91), .Y(SUM[31]) );
  OR2X2 U222 ( .A(A[22]), .B(B[22]), .Y(n146) );
  OR2X2 U223 ( .A(A[24]), .B(B[24]), .Y(n131) );
  OR2X2 U224 ( .A(A[26]), .B(B[26]), .Y(n113) );
  NAND2X1 U225 ( .A(B[26]), .B(A[26]), .Y(n118) );
  OR2X2 U226 ( .A(A[27]), .B(B[27]), .Y(n112) );
  NAND2X1 U227 ( .A(B[27]), .B(A[27]), .Y(n116) );
  NAND2X1 U228 ( .A(B[28]), .B(A[28]), .Y(n107) );
  OR2X2 U229 ( .A(A[28]), .B(B[28]), .Y(n105) );
  NAND2X1 U230 ( .A(B[30]), .B(A[30]), .Y(n92) );
  NAND2X1 U231 ( .A(B[29]), .B(A[29]), .Y(n98) );
  OR2X2 U232 ( .A(A[30]), .B(B[30]), .Y(n95) );
  OR2X2 U233 ( .A(A[29]), .B(B[29]), .Y(n99) );
  NAND2X2 U234 ( .A(B[3]), .B(A[3]), .Y(n77) );
  NAND3BX4 U235 ( .AN(n197), .B(n77), .C(n269), .Y(n60) );
  NAND3X4 U236 ( .A(n188), .B(n189), .C(n187), .Y(n183) );
  NOR2X2 U237 ( .A(n268), .B(n66), .Y(n273) );
  NAND2X4 U238 ( .A(n271), .B(n198), .Y(n269) );
  INVX4 U239 ( .A(n75), .Y(n271) );
  NAND2X2 U240 ( .A(B[1]), .B(A[1]), .Y(n90) );
  XOR2X2 U241 ( .A(n51), .B(n52), .Y(SUM[8]) );
  XOR2X4 U242 ( .A(n38), .B(n39), .Y(SUM[9]) );
  XOR2X4 U243 ( .A(n67), .B(n25), .Y(SUM[6]) );
  NAND2X4 U244 ( .A(n68), .B(n65), .Y(n67) );
  XOR2X4 U245 ( .A(n78), .B(n23), .Y(SUM[5]) );
  XOR2X4 U246 ( .A(n80), .B(n81), .Y(SUM[3]) );
  NOR2BX4 U247 ( .AN(n77), .B(n82), .Y(n81) );
  XOR2X4 U248 ( .A(n148), .B(n149), .Y(SUM[23]) );
  OAI21X4 U249 ( .A0(n150), .A1(n140), .B0(n139), .Y(n148) );
  XOR2X4 U250 ( .A(n151), .B(n152), .Y(SUM[22]) );
  NAND2X4 U251 ( .A(n147), .B(n154), .Y(n153) );
  NAND2X4 U252 ( .A(n134), .B(n143), .Y(n154) );
  NAND2X4 U253 ( .A(n20), .B(n156), .Y(n134) );
  XOR2X4 U254 ( .A(n173), .B(n174), .Y(SUM[1]) );
  XOR2X4 U255 ( .A(n176), .B(n177), .Y(SUM[19]) );
  OAI2BB1X4 U256 ( .A0N(n172), .A1N(n181), .B0(n169), .Y(n179) );
  NAND2X4 U257 ( .A(n159), .B(n168), .Y(n181) );
  NAND2X4 U258 ( .A(n183), .B(n184), .Y(n159) );
  OAI21X4 U259 ( .A0(n202), .A1(n203), .B0(n204), .Y(n201) );
  NAND2X4 U260 ( .A(n216), .B(n217), .Y(n193) );
  CLKINVX3 U261 ( .A(n219), .Y(n203) );
  XOR2X4 U262 ( .A(n221), .B(n222), .Y(SUM[15]) );
  AOI21X4 U263 ( .A0(n223), .A1(n224), .B0(n225), .Y(n222) );
  CLKINVX3 U264 ( .A(n205), .Y(n218) );
  OR2X4 U265 ( .A(A[15]), .B(B[15]), .Y(n219) );
  XOR2X4 U266 ( .A(n227), .B(n226), .Y(SUM[14]) );
  OR2X4 U267 ( .A(A[14]), .B(B[14]), .Y(n205) );
  XOR2X4 U268 ( .A(n224), .B(n230), .Y(SUM[13]) );
  OR2X4 U269 ( .A(A[13]), .B(B[13]), .Y(n228) );
  OAI21X4 U270 ( .A0(n231), .A1(n232), .B0(n18), .Y(n224) );
  XOR2X4 U271 ( .A(n239), .B(n240), .Y(SUM[12]) );
  CLKINVX3 U272 ( .A(n237), .Y(n220) );
  OR2X4 U273 ( .A(A[12]), .B(B[12]), .Y(n237) );
  NAND2X4 U274 ( .A(n249), .B(n250), .Y(n194) );
  CLKINVX3 U275 ( .A(n46), .Y(n49) );
  OAI21X4 U276 ( .A0(n42), .A1(n192), .B0(n252), .Y(n51) );
  XOR2X4 U277 ( .A(n253), .B(n26), .Y(SUM[11]) );
  NAND2BX4 U278 ( .AN(n254), .B(n255), .Y(n253) );
  OAI21X4 U279 ( .A0(n256), .A1(n257), .B0(n258), .Y(n255) );
  NOR3BX4 U280 ( .AN(n37), .B(n259), .C(n192), .Y(n257) );
  XOR2X4 U281 ( .A(n262), .B(n263), .Y(SUM[10]) );
  CLKINVX3 U282 ( .A(n258), .Y(n248) );
  OR2X4 U283 ( .A(A[10]), .B(B[10]), .Y(n258) );
  OR2X4 U284 ( .A(A[8]), .B(B[8]), .Y(n46) );
  OR2X4 U285 ( .A(A[9]), .B(B[9]), .Y(n251) );
  NAND2X4 U286 ( .A(n212), .B(n54), .Y(n45) );
  NAND3X4 U287 ( .A(n265), .B(n266), .C(n267), .Y(n212) );
  NAND3X4 U288 ( .A(n65), .B(n64), .C(n61), .Y(n267) );
  NAND2X4 U289 ( .A(B[4]), .B(A[4]), .Y(n61) );
  NAND2X4 U290 ( .A(B[5]), .B(A[5]), .Y(n65) );
  NOR2X4 U291 ( .A(n268), .B(n66), .Y(n266) );
  NAND2X4 U292 ( .A(n72), .B(n64), .Y(n265) );
  NAND3X4 U293 ( .A(n86), .B(n270), .C(n87), .Y(n75) );
  OR2X4 U294 ( .A(B[1]), .B(A[1]), .Y(n87) );
  OR2X4 U295 ( .A(A[2]), .B(B[2]), .Y(n86) );
  CLKINVX3 U296 ( .A(n76), .Y(n197) );
  NAND2BX4 U297 ( .AN(n85), .B(n270), .Y(n76) );
  OR2X4 U298 ( .A(A[3]), .B(B[3]), .Y(n270) );
  NAND2X4 U299 ( .A(n272), .B(n273), .Y(n192) );
  OR2X4 U300 ( .A(A[6]), .B(B[6]), .Y(n63) );
  CLKINVX3 U301 ( .A(n53), .Y(n268) );
  OR2X4 U302 ( .A(A[7]), .B(B[7]), .Y(n53) );
  NOR2X4 U303 ( .A(n72), .B(n73), .Y(n272) );
  CLKINVX3 U304 ( .A(n59), .Y(n73) );
  OR2X4 U305 ( .A(A[4]), .B(B[4]), .Y(n59) );
  OR2X4 U306 ( .A(A[5]), .B(B[5]), .Y(n62) );
endmodule


module hash_core_DW01_add_56 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n264, n265, n266, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263;

  NAND2X2 U2 ( .A(n50), .B(n195), .Y(n255) );
  NAND3BX2 U3 ( .AN(n172), .B(n162), .C(n173), .Y(n170) );
  NAND2X1 U4 ( .A(n57), .B(n58), .Y(n55) );
  NAND3BX4 U5 ( .AN(n196), .B(n190), .C(n191), .Y(n192) );
  AOI21X1 U6 ( .A0(n47), .A1(n48), .B0(n196), .Y(n228) );
  CLKINVX3 U7 ( .A(n235), .Y(n234) );
  NOR2BX4 U8 ( .AN(n191), .B(n196), .Y(n221) );
  CLKINVX8 U9 ( .A(n16), .Y(n169) );
  NAND3X4 U10 ( .A(n189), .B(n194), .C(n195), .Y(n193) );
  NAND2X2 U11 ( .A(n83), .B(n2), .Y(n3) );
  NAND2X2 U12 ( .A(n1), .B(n85), .Y(n4) );
  NAND2X4 U13 ( .A(n3), .B(n4), .Y(SUM[30]) );
  INVX1 U14 ( .A(n83), .Y(n1) );
  INVX2 U15 ( .A(n85), .Y(n2) );
  OR2X4 U16 ( .A(n38), .B(n87), .Y(n5) );
  NAND2X4 U17 ( .A(n5), .B(n88), .Y(n83) );
  CLKINVX3 U18 ( .A(n89), .Y(n87) );
  NAND2X2 U19 ( .A(n83), .B(n84), .Y(n82) );
  OR2X2 U20 ( .A(A[26]), .B(B[26]), .Y(n115) );
  NAND2XL U21 ( .A(n174), .B(n175), .Y(n6) );
  NAND2X4 U22 ( .A(n7), .B(n153), .Y(n173) );
  INVX1 U23 ( .A(n6), .Y(n7) );
  OR2X2 U24 ( .A(n33), .B(n136), .Y(n8) );
  NAND2X1 U25 ( .A(n8), .B(n137), .Y(n135) );
  NOR2X2 U26 ( .A(A[21]), .B(B[21]), .Y(n33) );
  NAND2X2 U27 ( .A(B[20]), .B(A[20]), .Y(n136) );
  NAND2X1 U28 ( .A(B[21]), .B(A[21]), .Y(n137) );
  NAND2BX4 U29 ( .AN(n134), .B(n135), .Y(n131) );
  NAND2XL U30 ( .A(n181), .B(n180), .Y(n9) );
  AND2X2 U31 ( .A(n182), .B(n10), .Y(n21) );
  INVX2 U32 ( .A(n9), .Y(n10) );
  NAND3X4 U33 ( .A(n199), .B(n198), .C(n197), .Y(n181) );
  NOR4X4 U34 ( .A(n35), .B(n34), .C(n155), .D(n156), .Y(n154) );
  INVX2 U35 ( .A(n195), .Y(n53) );
  INVX4 U36 ( .A(n91), .Y(n165) );
  AOI21X4 U37 ( .A0(n59), .A1(n41), .B0(n61), .Y(n54) );
  OAI21X4 U38 ( .A0(n169), .A1(n34), .B0(n159), .Y(n167) );
  NAND2BX4 U39 ( .AN(n34), .B(n160), .Y(n158) );
  OAI21X4 U40 ( .A0(n155), .A1(n161), .B0(n162), .Y(n160) );
  INVX2 U41 ( .A(n190), .Y(n218) );
  NAND2X2 U42 ( .A(n153), .B(n154), .Y(n152) );
  NAND2XL U43 ( .A(n153), .B(n22), .Y(n23) );
  OAI21X4 U44 ( .A0(n101), .A1(n102), .B0(n103), .Y(n97) );
  NOR2X2 U45 ( .A(n104), .B(n105), .Y(n103) );
  XOR2X4 U46 ( .A(n97), .B(n99), .Y(SUM[28]) );
  XOR2X4 U47 ( .A(n74), .B(n75), .Y(SUM[3]) );
  NOR2BX1 U48 ( .AN(n138), .B(n133), .Y(n143) );
  INVX4 U49 ( .A(n141), .Y(n133) );
  BUFX4 U50 ( .A(n266), .Y(SUM[20]) );
  CLKINVX8 U51 ( .A(n39), .Y(SUM[21]) );
  XOR2X4 U52 ( .A(n79), .B(n90), .Y(SUM[2]) );
  NOR2BX2 U53 ( .AN(n78), .B(n37), .Y(n90) );
  NOR2BX4 U54 ( .AN(n166), .B(n30), .Y(SUM[0]) );
  NAND2X4 U55 ( .A(B[0]), .B(A[0]), .Y(n166) );
  OR2X4 U56 ( .A(A[16]), .B(B[16]), .Y(n175) );
  XOR2X2 U57 ( .A(n92), .B(n164), .Y(SUM[1]) );
  NAND2X2 U58 ( .A(B[17]), .B(A[17]), .Y(n162) );
  NOR2BX4 U59 ( .AN(n132), .B(n134), .Y(n146) );
  INVX12 U60 ( .A(n140), .Y(n134) );
  INVX4 U61 ( .A(n161), .Y(n178) );
  NOR2BX4 U62 ( .AN(n161), .B(n156), .Y(n179) );
  NOR2X4 U63 ( .A(n161), .B(n155), .Y(n172) );
  NAND2X2 U64 ( .A(B[16]), .B(A[16]), .Y(n161) );
  NAND2X2 U65 ( .A(n47), .B(n48), .Y(n46) );
  CLKINVX2 U66 ( .A(n166), .Y(n92) );
  CLKINVX3 U67 ( .A(n174), .Y(n155) );
  INVX1 U68 ( .A(n175), .Y(n156) );
  OR2X2 U69 ( .A(A[23]), .B(B[23]), .Y(n141) );
  OR2X2 U70 ( .A(A[22]), .B(B[22]), .Y(n140) );
  INVX4 U71 ( .A(n239), .Y(n45) );
  CLKBUFX3 U72 ( .A(B[7]), .Y(n19) );
  BUFX12 U73 ( .A(n60), .Y(n41) );
  INVX1 U74 ( .A(n201), .Y(n250) );
  CLKINVX3 U75 ( .A(n265), .Y(n39) );
  XOR2X2 U76 ( .A(n89), .B(n94), .Y(SUM[29]) );
  OAI21X2 U77 ( .A0(n119), .A1(n109), .B0(n107), .Y(n117) );
  XOR2X2 U78 ( .A(n123), .B(n124), .Y(SUM[25]) );
  NAND2BX2 U79 ( .AN(n243), .B(n244), .Y(n242) );
  INVX1 U80 ( .A(n44), .Y(n248) );
  NOR2BX1 U81 ( .AN(n93), .B(n165), .Y(n164) );
  AND2X2 U82 ( .A(n50), .B(n41), .Y(n12) );
  NOR2BX1 U83 ( .AN(n44), .B(n45), .Y(n43) );
  NAND2X1 U84 ( .A(B[6]), .B(A[6]), .Y(n56) );
  INVX1 U85 ( .A(B[5]), .Y(n261) );
  AND3X2 U86 ( .A(n139), .B(n140), .C(n141), .Y(n13) );
  INVX4 U87 ( .A(n189), .Y(n203) );
  OAI21X2 U88 ( .A0(n77), .A1(n37), .B0(n78), .Y(n74) );
  OAI2BB1X4 U89 ( .A0N(n229), .A1N(n230), .B0(n231), .Y(n14) );
  OAI2BB1X2 U90 ( .A0N(n229), .A1N(n230), .B0(n231), .Y(n186) );
  CLKBUFX3 U91 ( .A(n233), .Y(n15) );
  NAND3X2 U92 ( .A(A[12]), .B(B[12]), .C(n190), .Y(n210) );
  NOR2X4 U93 ( .A(n236), .B(n232), .Y(n229) );
  INVX1 U94 ( .A(n225), .Y(n224) );
  NAND2X1 U95 ( .A(B[12]), .B(A[12]), .Y(n225) );
  INVX2 U96 ( .A(n149), .Y(n128) );
  AOI21X2 U97 ( .A0(n44), .A1(n49), .B0(n45), .Y(n230) );
  NAND3BX4 U98 ( .AN(n172), .B(n162), .C(n173), .Y(n16) );
  NOR2BX4 U99 ( .AN(n63), .B(n41), .Y(n67) );
  NAND3X1 U100 ( .A(n49), .B(n245), .C(n246), .Y(n244) );
  BUFX2 U101 ( .A(B[14]), .Y(n17) );
  OAI2BB1X2 U102 ( .A0N(A[7]), .A1N(B[7]), .B0(n263), .Y(n256) );
  NAND2BX4 U103 ( .AN(n256), .B(n257), .Y(n18) );
  NAND2X1 U104 ( .A(B[19]), .B(A[19]), .Y(n163) );
  OAI2BB1X4 U105 ( .A0N(n59), .A1N(n41), .B0(n63), .Y(n69) );
  AOI21X4 U106 ( .A0(n183), .A1(n18), .B0(n185), .Y(n182) );
  INVX4 U107 ( .A(n219), .Y(n217) );
  NAND2X4 U108 ( .A(n95), .B(n96), .Y(n89) );
  NAND2X4 U109 ( .A(n97), .B(n98), .Y(n95) );
  AOI21X4 U110 ( .A0(n194), .A1(n213), .B0(n214), .Y(n212) );
  NOR3BX4 U111 ( .AN(n186), .B(n187), .C(n188), .Y(n185) );
  OAI21X2 U112 ( .A0(n17), .A1(A[14]), .B0(n191), .Y(n187) );
  XOR2X4 U113 ( .A(n226), .B(n227), .Y(SUM[12]) );
  NAND2BX2 U114 ( .AN(n53), .B(n18), .Y(n47) );
  NOR2BX4 U115 ( .AN(n208), .B(n218), .Y(n220) );
  OAI21X2 U116 ( .A0(n54), .A1(n55), .B0(n56), .Y(n51) );
  NAND4BX4 U117 ( .AN(n254), .B(n57), .C(n58), .D(n59), .Y(n200) );
  NAND3X4 U118 ( .A(n245), .B(n49), .C(n246), .Y(n20) );
  INVX4 U119 ( .A(n57), .Y(n71) );
  NAND2X4 U120 ( .A(B[8]), .B(A[8]), .Y(n49) );
  NAND3X2 U121 ( .A(n245), .B(n49), .C(n246), .Y(n42) );
  NOR3BX2 U122 ( .AN(n191), .B(n196), .C(n200), .Y(n199) );
  NAND2X2 U123 ( .A(n21), .B(n179), .Y(n24) );
  NAND2X4 U124 ( .A(n23), .B(n24), .Y(SUM[16]) );
  INVXL U125 ( .A(n179), .Y(n22) );
  AOI21X2 U126 ( .A0(n93), .A1(n166), .B0(n165), .Y(n251) );
  NOR2X2 U127 ( .A(B[7]), .B(A[7]), .Y(n254) );
  NAND2BX2 U128 ( .AN(A[5]), .B(n261), .Y(n259) );
  BUFX4 U129 ( .A(n264), .Y(SUM[24]) );
  NAND2X4 U130 ( .A(n251), .B(n252), .Y(n202) );
  NOR2BX2 U131 ( .AN(n253), .B(n37), .Y(n252) );
  INVX4 U132 ( .A(n79), .Y(n77) );
  NAND2X4 U133 ( .A(B[25]), .B(A[25]), .Y(n113) );
  NOR2X2 U134 ( .A(n14), .B(n228), .Y(n227) );
  NAND2X2 U135 ( .A(n27), .B(n125), .Y(n101) );
  NAND2X4 U136 ( .A(n12), .B(n249), .Y(n246) );
  INVX2 U137 ( .A(n200), .Y(n249) );
  OR2XL U138 ( .A(A[24]), .B(B[24]), .Y(n125) );
  INVX4 U139 ( .A(n145), .Y(n144) );
  NAND2X1 U140 ( .A(B[18]), .B(A[18]), .Y(n159) );
  NOR2X4 U141 ( .A(A[18]), .B(B[18]), .Y(n34) );
  NOR2BX1 U142 ( .AN(n163), .B(n35), .Y(n168) );
  NOR2BXL U143 ( .AN(n114), .B(n108), .Y(n118) );
  INVX1 U144 ( .A(n120), .Y(n119) );
  NAND2X2 U145 ( .A(B[24]), .B(A[24]), .Y(n112) );
  NAND2X1 U146 ( .A(B[13]), .B(A[13]), .Y(n208) );
  NAND2X1 U147 ( .A(B[10]), .B(A[10]), .Y(n233) );
  AOI21X2 U148 ( .A0(n158), .A1(n159), .B0(n35), .Y(n157) );
  NAND2XL U149 ( .A(n49), .B(n50), .Y(n26) );
  NOR2BX1 U150 ( .AN(n88), .B(n38), .Y(n94) );
  NAND3BXL U151 ( .AN(n111), .B(n115), .C(n116), .Y(n102) );
  INVXL U152 ( .A(n215), .Y(n214) );
  INVX1 U153 ( .A(n116), .Y(n108) );
  NOR2X4 U154 ( .A(A[2]), .B(B[2]), .Y(n37) );
  NAND2X2 U155 ( .A(B[3]), .B(A[3]), .Y(n76) );
  OAI2BB1X4 U156 ( .A0N(n91), .A1N(n92), .B0(n93), .Y(n79) );
  INVX4 U157 ( .A(n115), .Y(n109) );
  INVX2 U158 ( .A(n122), .Y(n111) );
  NOR2BXL U159 ( .AN(n107), .B(n109), .Y(n121) );
  XOR2X4 U160 ( .A(n145), .B(n146), .Y(SUM[22]) );
  INVX1 U161 ( .A(n33), .Y(n31) );
  XNOR2X4 U162 ( .A(n26), .B(n46), .Y(SUM[8]) );
  NOR2BX2 U163 ( .AN(n163), .B(n157), .Y(n151) );
  OAI2BB1X4 U164 ( .A0N(n13), .A1N(n149), .B0(n28), .Y(n27) );
  NOR2X4 U165 ( .A(n129), .B(n130), .Y(n28) );
  CLKINVX3 U166 ( .A(n207), .Y(n206) );
  AND2X1 U167 ( .A(n215), .B(n194), .Y(n216) );
  XOR2X4 U168 ( .A(n240), .B(n29), .Y(SUM[11]) );
  AND2X1 U169 ( .A(n235), .B(n237), .Y(n29) );
  NOR2XL U170 ( .A(A[0]), .B(B[0]), .Y(n30) );
  NAND2XL U171 ( .A(B[26]), .B(A[26]), .Y(n107) );
  NAND2XL U172 ( .A(B[27]), .B(A[27]), .Y(n114) );
  NOR2X2 U173 ( .A(A[20]), .B(B[20]), .Y(n36) );
  NAND2XL U174 ( .A(B[30]), .B(A[30]), .Y(n81) );
  NAND2XL U175 ( .A(B[28]), .B(A[28]), .Y(n96) );
  OR2X4 U176 ( .A(A[17]), .B(B[17]), .Y(n174) );
  INVX4 U177 ( .A(n56), .Y(n260) );
  NAND2XL U178 ( .A(n225), .B(n191), .Y(n226) );
  INVX1 U179 ( .A(n114), .Y(n104) );
  OAI2BB1X4 U180 ( .A0N(n147), .A1N(n31), .B0(n137), .Y(n145) );
  XOR2X2 U181 ( .A(n120), .B(n121), .Y(SUM[26]) );
  NOR2BX1 U182 ( .AN(n159), .B(n34), .Y(n171) );
  XOR2X1 U183 ( .A(n27), .B(n126), .Y(n264) );
  NOR2BX1 U184 ( .AN(n112), .B(n127), .Y(n126) );
  INVX1 U185 ( .A(n125), .Y(n127) );
  NOR2BX1 U186 ( .AN(n81), .B(n86), .Y(n85) );
  INVX1 U187 ( .A(n84), .Y(n86) );
  NOR2BX1 U188 ( .AN(n96), .B(n100), .Y(n99) );
  INVX1 U189 ( .A(n98), .Y(n100) );
  NAND2X1 U190 ( .A(n162), .B(n174), .Y(n176) );
  XOR2X1 U191 ( .A(n149), .B(n150), .Y(n266) );
  NOR2BX1 U192 ( .AN(n136), .B(n36), .Y(n150) );
  NOR2BX1 U193 ( .AN(n113), .B(n111), .Y(n124) );
  AOI21X1 U194 ( .A0(n106), .A1(n107), .B0(n108), .Y(n105) );
  NAND2BX1 U195 ( .AN(n109), .B(n110), .Y(n106) );
  OAI21XL U196 ( .A0(n111), .A1(n112), .B0(n113), .Y(n110) );
  XNOR2X4 U197 ( .A(n32), .B(n247), .Y(SUM[10]) );
  AND2X1 U198 ( .A(n15), .B(n238), .Y(n32) );
  OAI21XL U199 ( .A0(n236), .A1(n44), .B0(n15), .Y(n241) );
  INVX1 U200 ( .A(n138), .Y(n129) );
  NAND2XL U201 ( .A(n238), .B(n239), .Y(n243) );
  AND2X2 U202 ( .A(n194), .B(n190), .Y(n198) );
  NOR2BX1 U203 ( .AN(n137), .B(n33), .Y(n148) );
  NOR2X4 U204 ( .A(A[19]), .B(B[19]), .Y(n35) );
  NAND2X2 U205 ( .A(B[9]), .B(A[9]), .Y(n44) );
  NAND2X2 U206 ( .A(B[4]), .B(A[4]), .Y(n63) );
  AND2X2 U207 ( .A(n189), .B(n194), .Y(n204) );
  NAND2X1 U208 ( .A(B[22]), .B(A[22]), .Y(n132) );
  NAND2X2 U209 ( .A(B[1]), .B(A[1]), .Y(n93) );
  NAND2XL U210 ( .A(B[4]), .B(A[4]), .Y(n262) );
  NAND2XL U211 ( .A(B[15]), .B(A[15]), .Y(n207) );
  OR2X2 U212 ( .A(A[27]), .B(B[27]), .Y(n116) );
  OR2X2 U213 ( .A(A[25]), .B(B[25]), .Y(n122) );
  NOR2X1 U214 ( .A(A[29]), .B(B[29]), .Y(n38) );
  NAND2X1 U215 ( .A(B[29]), .B(A[29]), .Y(n88) );
  OR2X2 U216 ( .A(A[28]), .B(B[28]), .Y(n98) );
  OR2X2 U217 ( .A(A[30]), .B(B[30]), .Y(n84) );
  XOR3X2 U218 ( .A(B[31]), .B(A[31]), .C(n80), .Y(SUM[31]) );
  NAND2X1 U219 ( .A(n81), .B(n82), .Y(n80) );
  NAND3BX4 U220 ( .AN(n250), .B(n76), .C(n202), .Y(n60) );
  NAND3X4 U221 ( .A(n181), .B(n182), .C(n180), .Y(n153) );
  NAND2XL U222 ( .A(n17), .B(A[14]), .Y(n215) );
  NAND2XL U223 ( .A(B[14]), .B(A[14]), .Y(n209) );
  NAND3X2 U224 ( .A(n208), .B(n209), .C(n210), .Y(n205) );
  OAI2BB1X1 U225 ( .A0N(n195), .A1N(n184), .B0(n48), .Y(n222) );
  AOI21X2 U226 ( .A0(n175), .A1(n153), .B0(n178), .Y(n177) );
  XOR2X4 U227 ( .A(n219), .B(n220), .Y(SUM[13]) );
  CLKINVX8 U228 ( .A(n58), .Y(n66) );
  NAND3X4 U229 ( .A(A[5]), .B(n58), .C(B[5]), .Y(n263) );
  AND2X1 U230 ( .A(n76), .B(n253), .Y(n75) );
  NAND2X1 U231 ( .A(B[23]), .B(A[23]), .Y(n138) );
  INVX4 U232 ( .A(n238), .Y(n236) );
  NAND2X2 U233 ( .A(B[5]), .B(A[5]), .Y(n62) );
  NAND2X1 U234 ( .A(B[11]), .B(A[11]), .Y(n235) );
  XOR2X4 U235 ( .A(n211), .B(n212), .Y(SUM[15]) );
  INVX4 U236 ( .A(n237), .Y(n232) );
  AOI21X2 U237 ( .A0(n19), .A1(A[7]), .B0(n53), .Y(n52) );
  XOR2X1 U238 ( .A(n147), .B(n148), .Y(n265) );
  NAND2XL U239 ( .A(n207), .B(n189), .Y(n211) );
  XOR2X4 U240 ( .A(n42), .B(n43), .Y(SUM[9]) );
  XOR2X4 U241 ( .A(n51), .B(n52), .Y(SUM[7]) );
  NAND2X4 U242 ( .A(n62), .B(n63), .Y(n61) );
  XOR2X4 U243 ( .A(n64), .B(n65), .Y(SUM[6]) );
  NOR2BX4 U244 ( .AN(n56), .B(n66), .Y(n65) );
  OAI21X4 U245 ( .A0(n67), .A1(n68), .B0(n62), .Y(n64) );
  NAND2X4 U246 ( .A(n59), .B(n57), .Y(n68) );
  XOR2X4 U247 ( .A(n69), .B(n70), .Y(SUM[5]) );
  NOR2BX4 U248 ( .AN(n62), .B(n71), .Y(n70) );
  OR2X4 U249 ( .A(A[5]), .B(B[5]), .Y(n57) );
  XOR2X4 U250 ( .A(n41), .B(n72), .Y(SUM[4]) );
  NOR2BX4 U251 ( .AN(n63), .B(n73), .Y(n72) );
  CLKINVX3 U252 ( .A(n59), .Y(n73) );
  XOR2X4 U253 ( .A(n117), .B(n118), .Y(SUM[27]) );
  OAI2BB1X4 U254 ( .A0N(n122), .A1N(n123), .B0(n113), .Y(n120) );
  NAND2X4 U255 ( .A(n101), .B(n112), .Y(n123) );
  AOI21X4 U256 ( .A0(n131), .A1(n132), .B0(n133), .Y(n130) );
  NOR2X4 U257 ( .A(n33), .B(n36), .Y(n139) );
  XOR2X4 U258 ( .A(n142), .B(n143), .Y(SUM[23]) );
  OAI21X4 U259 ( .A0(n144), .A1(n134), .B0(n132), .Y(n142) );
  OAI21X4 U260 ( .A0(n36), .A1(n128), .B0(n136), .Y(n147) );
  NAND2X4 U261 ( .A(n151), .B(n152), .Y(n149) );
  XOR2X4 U262 ( .A(n167), .B(n168), .Y(SUM[19]) );
  XOR2X4 U263 ( .A(n170), .B(n171), .Y(SUM[18]) );
  XOR2X4 U264 ( .A(n176), .B(n177), .Y(SUM[17]) );
  NAND2X4 U265 ( .A(n189), .B(n190), .Y(n188) );
  NOR2X4 U266 ( .A(n192), .B(n193), .Y(n183) );
  AOI31X2 U267 ( .A0(n76), .A1(n201), .A2(n202), .B0(n203), .Y(n197) );
  AOI21X4 U268 ( .A0(n204), .A1(n205), .B0(n206), .Y(n180) );
  OR2X4 U269 ( .A(A[15]), .B(B[15]), .Y(n189) );
  XOR2X4 U270 ( .A(n213), .B(n216), .Y(SUM[14]) );
  OR2X4 U271 ( .A(B[14]), .B(A[14]), .Y(n194) );
  OAI21X4 U272 ( .A0(n217), .A1(n218), .B0(n208), .Y(n213) );
  OR2X4 U273 ( .A(A[13]), .B(B[13]), .Y(n190) );
  OAI2BB1X4 U274 ( .A0N(n221), .A1N(n222), .B0(n223), .Y(n219) );
  AOI21X4 U275 ( .A0(n14), .A1(n191), .B0(n224), .Y(n223) );
  AOI2BB1X4 U276 ( .A0N(n232), .A1N(n233), .B0(n234), .Y(n231) );
  NAND4BX4 U277 ( .AN(n45), .B(n50), .C(n237), .D(n238), .Y(n196) );
  NAND2BX4 U278 ( .AN(n200), .B(n41), .Y(n48) );
  OR2X4 U279 ( .A(A[12]), .B(B[12]), .Y(n191) );
  OR2X4 U280 ( .A(A[11]), .B(B[11]), .Y(n237) );
  NAND2BX4 U281 ( .AN(n241), .B(n242), .Y(n240) );
  AOI21X4 U282 ( .A0(n239), .A1(n20), .B0(n248), .Y(n247) );
  OR2X4 U283 ( .A(A[1]), .B(B[1]), .Y(n91) );
  NAND2BX4 U284 ( .AN(n78), .B(n253), .Y(n201) );
  OR2X4 U285 ( .A(A[3]), .B(B[3]), .Y(n253) );
  NAND2X4 U286 ( .A(B[2]), .B(A[2]), .Y(n78) );
  OR2X4 U287 ( .A(A[4]), .B(B[4]), .Y(n59) );
  NAND2BX4 U288 ( .AN(n255), .B(n184), .Y(n245) );
  NAND2BX4 U289 ( .AN(n256), .B(n257), .Y(n184) );
  AOI21X4 U290 ( .A0(n258), .A1(n259), .B0(n260), .Y(n257) );
  NOR2X4 U291 ( .A(n262), .B(n66), .Y(n258) );
  OR2X4 U292 ( .A(A[6]), .B(B[6]), .Y(n58) );
  OR2X4 U293 ( .A(B[7]), .B(A[7]), .Y(n195) );
  OR2X4 U294 ( .A(A[8]), .B(B[8]), .Y(n50) );
  OR2X4 U295 ( .A(A[9]), .B(B[9]), .Y(n239) );
  OR2X4 U296 ( .A(A[10]), .B(B[10]), .Y(n238) );
endmodule


module hash_core ( clk, reset, Wt, inner_busy, first_block, output_enable, 
        digest );
  input [31:0] Wt;
  output [31:0] digest;
  input clk, reset, inner_busy, first_block, output_enable;
  wire   N121, N122, N123, N124, N125, N126, N127, N795, N796, N797, N798,
         N799, N800, N801, N802, N803, N804, N805, N806, N807, N808, N809,
         N810, N811, N812, N813, N814, N815, N816, N817, N818, N819, N820,
         N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831,
         N832, N833, N834, N835, N836, N837, N838, N839, N840, N841, N842,
         N843, N844, N845, N846, N847, N848, N849, N850, N851, N852, N853,
         N854, N855, N856, N857, N858, N859, N860, N861, N862, N863, N864,
         N865, N866, N867, N868, N869, N870, N871, N872, N873, N874, N875,
         N876, N877, N878, N879, N880, N881, N882, N883, N884, N885, N886,
         N887, N888, N889, N890, N891, N892, N893, N894, N895, N896, N897,
         N898, N899, N900, N901, N902, N903, N904, N905, N906, N907, N908,
         N909, N910, N911, N912, N913, N914, N915, N916, N917, N918, N919,
         N920, N921, N922, N923, N924, N925, N926, N927, N928, N929, N930,
         N931, N932, N933, N934, N935, N936, N937, N938, N939, N940, N941,
         N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952,
         N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963,
         N964, N965, N966, N967, N968, N969, N970, N971, N972, N973, N974,
         N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985,
         N986, N987, N988, N989, N990, N991, N992, N993, N994, N995, N996,
         N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006,
         N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016,
         N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026,
         N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036,
         N1037, N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046,
         N1047, N1048, N1049, N1050, N2946, N2947, N2948, N2949, N2950, N2951,
         N2952, N2953, N2954, N2955, N2956, N2957, N2958, N2959, N2960, N2961,
         N2962, N2963, N2964, N2965, N2966, N2967, N2968, N2969, N2970, N2971,
         N2972, N2973, N2974, N2975, N2976, N2977, N3047, N3048, N3049, N3050,
         N3051, N3052, N3053, N3054, N3055, N3056, N3057, N3058, N3059, N3060,
         N3061, N3062, N3063, N3064, N3065, N3066, N3067, N3068, N3069, N3070,
         N3071, N3072, N3073, N3074, N3075, N3076, N3077, N3078, N3079, N3080,
         N3081, n1140, n1141, n1142, n1143, n1144, n1145, n1151, n1152, n1153,
         n1154, n1156, n1157, n1160, n1161, n1163, n1165, n1167, n1168, n1370,
         n1383, n1388, n1393, n1396, n1434, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1456, n1457, n1458, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1487, n1488, n1489, n1490, n1491, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1611, n1612, n1615,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1631, n1632, n1633, n1635, n1636, n1640, n1641,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1720, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1755, n1756,
         n1757, n1758, n1759, n1760, n1763, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1785, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1849, n1859, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1878, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1984, n1985, n1986, n1990, n1991, n1992, n1994, n1995, n1996, n1998,
         n1999, n2000, n2002, n2003, n2004, n2006, n2007, n2008, n2010, n2011,
         n2012, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2070, n2071, n2072, n2074,
         n2075, n2076, n2078, n2079, n2080, n2082, n2083, n2084, n2086, n2087,
         n2088, n2090, n2091, n2092, n2094, n2095, n2096, n2098, n2099, n2100,
         n2102, n2103, n2104, n2106, n2107, n2108, n2110, n2111, n2112, n2114,
         n2116, n2117, n2118, n2119, n2121, n2122, n2124, n2125, n2126, n2127,
         n2128, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, T2_32_9_, T2_32_8_, T2_32_7_,
         T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_, T2_32_31_, T2_32_30_,
         T2_32_2_, T2_32_29_, T2_32_28_, T2_32_27_, T2_32_26_, T2_32_25_,
         T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_, T2_32_20_, T2_32_1_,
         T2_32_19_, T2_32_18_, T2_32_17_, T2_32_16_, T2_32_15_, T2_32_14_,
         T2_32_13_, T2_32_12_, T2_32_11_, T2_32_10_, T2_32_0_, N99, N98, N97,
         N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83,
         N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69,
         N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55,
         N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41,
         N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27,
         N26, N25, N24, N119, N118, N117, N116, N115, N114, N113, N112, N111,
         N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973;
  wire   [31:0] f1_EFG_32;
  wire   [31:0] f2_ABC_32;
  wire   [31:0] f3_A_32;
  wire   [31:0] f4_E_32;
  wire   [31:0] Kt;
  wire   [31:0] T1_32;
  wire   [31:0] next_E;
  wire   [31:0] next_A;
  wire   [255:0] SHA256_result;
  wire   [6:1] round;
  wire   [31:0] H0;
  wire   [31:0] H1;
  wire   [31:1] H2;
  wire   [31:0] H3;
  wire   [31:0] H4;
  wire   [31:0] H5;
  wire   [31:0] H6;
  wire   [31:0] H7;
  wire   [2:0] read_counter;

  DFFHQX4 C_reg_0_ ( .D(n2798), .CK(clk), .Q(SHA256_result[160]) );
  DFFHQX4 E_reg_0_ ( .D(n2734), .CK(clk), .Q(SHA256_result[96]) );
  DFFHQX4 E_reg_1_ ( .D(n2733), .CK(clk), .Q(SHA256_result[97]) );
  DFFHQX4 E_reg_2_ ( .D(n2732), .CK(clk), .Q(SHA256_result[98]) );
  DFFHQX4 E_reg_4_ ( .D(n2730), .CK(clk), .Q(SHA256_result[100]) );
  DFFHQX4 E_reg_6_ ( .D(n2728), .CK(clk), .Q(SHA256_result[102]) );
  DFFHQX4 E_reg_8_ ( .D(n2726), .CK(clk), .Q(SHA256_result[104]) );
  DFFHQX4 E_reg_9_ ( .D(n2725), .CK(clk), .Q(SHA256_result[105]) );
  DFFHQX4 E_reg_10_ ( .D(n2724), .CK(clk), .Q(SHA256_result[106]) );
  DFFHQX4 E_reg_11_ ( .D(n2723), .CK(clk), .Q(SHA256_result[107]) );
  DFFHQX4 E_reg_12_ ( .D(n2722), .CK(clk), .Q(SHA256_result[108]) );
  DFFHQX4 E_reg_13_ ( .D(n2721), .CK(clk), .Q(SHA256_result[109]) );
  DFFHQX4 E_reg_14_ ( .D(n2720), .CK(clk), .Q(SHA256_result[110]) );
  DFFHQX4 E_reg_15_ ( .D(n2719), .CK(clk), .Q(SHA256_result[111]) );
  DFFX4 F_reg_1_ ( .D(n2701), .CK(clk), .Q(SHA256_result[65]), .QN(n1167) );
  DFFHQX4 G_reg_1_ ( .D(n2510), .CK(clk), .Q(SHA256_result[33]) );
  DFFHQX4 G_reg_5_ ( .D(n2506), .CK(clk), .Q(SHA256_result[37]) );
  DFFHQX4 Kt_reg_13_ ( .D(N2959), .CK(clk), .Q(Kt[13]) );
  DFFHQX4 Kt_reg_8_ ( .D(N2954), .CK(clk), .Q(Kt[8]) );
  DFFHQX4 Kt_reg_6_ ( .D(N2952), .CK(clk), .Q(Kt[6]) );
  DFFHQX4 Kt_reg_4_ ( .D(N2950), .CK(clk), .Q(Kt[4]) );
  DFFHQX4 Kt_reg_3_ ( .D(N2949), .CK(clk), .Q(Kt[3]) );
  DFFHQX4 Kt_reg_2_ ( .D(N2948), .CK(clk), .Q(Kt[2]) );
  DFFHQX4 Kt_reg_1_ ( .D(N2947), .CK(clk), .Q(Kt[1]) );
  DFFHQX4 Kt_reg_0_ ( .D(N2946), .CK(clk), .Q(Kt[0]) );
  AND2X2 U1425 ( .A(n2232), .B(n1393), .Y(n2171) );
  CLKINVX4 U2005 ( .A(reset), .Y(n1434) );
  hash_core_DW01_add_0 add_317 ( .A({SHA256_result[63:39], n50, 
        SHA256_result[37:33], n82}), .B(H7), .SUM({N1050, N1049, N1048, N1047, 
        N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, 
        N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, 
        N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019}) );
  hash_core_DW01_add_1 add_316 ( .A(SHA256_result[95:64]), .B({H6[31:2], n96, 
        H6[0]}), .SUM({N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, 
        N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, 
        N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, 
        N989, N988, N987}) );
  hash_core_DW01_add_2 add_315 ( .A({SHA256_result[127:126], n51, 
        SHA256_result[124:98], n69, SHA256_result[96]}), .B(H5), .SUM({N986, 
        N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, 
        N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, 
        N961, N960, N959, N958, N957, N956, N955}) );
  hash_core_DW01_add_4 add_313 ( .A(SHA256_result[191:160]), .B({H3[31:2], n71, 
        H3[0]}), .SUM({N922, N921, N920, N919, N918, N917, N916, N915, N914, 
        N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, 
        N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891}) );
  hash_core_DW01_add_5 add_312 ( .A({SHA256_result[223:194], n79, n89}), .B({
        H2, n99}), .SUM({N890, N889, N888, N887, N886, N885, N884, N883, N882, 
        N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, 
        N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859}) );
  hash_core_DW01_add_6 add_311 ( .A({n25, n131, n132, SHA256_result[252], n133, 
        n134, n135, n136, n137, SHA256_result[246], n138, n139, n140, n141, 
        n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
        n154, n155, n156, n157, n65, SHA256_result[224]}), .B(H1), .SUM({N858, 
        N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, 
        N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, 
        N833, N832, N831, N830, N829, N828, N827}) );
  hash_core_DW01_inc_0 add_119 ( .A({round[6], n160, n159, round[3:2], n347, 
        n161}), .SUM({N127, N126, N125, N124, N123, N122, N121}) );
  hash_core_DW01_add_16 add_314 ( .A({next_E[31:19], n47, next_E[17:0]}), .B(
        H4), .SUM({N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, 
        N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, 
        N932, N931, N930, N929, N928, N927, N926, N925, N924, N923}) );
  hash_core_DW01_add_18 add_310 ( .A({next_A[31:21], n43, next_A[19:0]}), .B(
        H0), .SUM({N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, 
        N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, 
        N804, N803, N802, N801, N800, N799, N798, N797, N796, N795}) );
  hash_core_DW01_add_26 add_1_root_add_0_root_add_113 ( .A(f2_ABC_32), .B(
        f3_A_32), .SUM({T2_32_31_, T2_32_30_, T2_32_29_, T2_32_28_, T2_32_27_, 
        T2_32_26_, T2_32_25_, T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_, 
        T2_32_20_, T2_32_19_, T2_32_18_, T2_32_17_, T2_32_16_, T2_32_15_, 
        T2_32_14_, T2_32_13_, T2_32_12_, T2_32_11_, T2_32_10_, T2_32_9_, 
        T2_32_8_, T2_32_7_, T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_, T2_32_2_, 
        T2_32_1_, T2_32_0_}) );
  hash_core_DW01_add_24 add_0_root_add_0_root_add_108_4 ( .A({N119, N118, N117, 
        N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, 
        N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, 
        N91, N90, N89, N88}), .B({N87, N86, N85, N84, N83, N82, N81, N80, N79, 
        N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, 
        N64, N63, N62, N61, N60, N59, N58, N57, N56}), .SUM(T1_32) );
  hash_core_DW01_add_38 add_112 ( .A(SHA256_result[159:128]), .B({T1_32[31:14], 
        n45, T1_32[12:0]}), .SUM(next_E) );
  hash_core_DW01_add_40 add_0_root_add_0_root_add_113 ( .A({T2_32_31_, 
        T2_32_30_, T2_32_29_, T2_32_28_, T2_32_27_, T2_32_26_, T2_32_25_, 
        T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_, T2_32_20_, T2_32_19_, 
        T2_32_18_, T2_32_17_, T2_32_16_, T2_32_15_, T2_32_14_, T2_32_13_, 
        T2_32_12_, T2_32_11_, T2_32_10_, T2_32_9_, T2_32_8_, T2_32_7_, 
        T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_, T2_32_2_, T2_32_1_, T2_32_0_}), 
        .B({T1_32[31:14], n45, T1_32[12:0]}), .SUM(next_A) );
  hash_core_DW01_add_46 add_2_root_add_0_root_add_108_4 ( .A(
        SHA256_result[31:0]), .B({f1_EFG_32[31:5], n40, f1_EFG_32[3], n39, 
        f1_EFG_32[1:0]}), .SUM({N119, N118, N117, N116, N115, N114, N113, N112, 
        N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, 
        N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88}) );
  hash_core_DW01_add_50 add_3_root_add_0_root_add_108_4 ( .A(Kt), .B(Wt), 
        .SUM({N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24}) );
  hash_core_DW01_add_56 add_1_root_add_0_root_add_108_4 ( .A(f4_E_32), .B({N55, 
        N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, 
        N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24}), .SUM({N87, N86, N85, N84, N83, N82, N81, N80, N79, 
        N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, 
        N64, N63, N62, N61, N60, N59, N58, N57, N56}) );
  DFFHQX1 read_counter_reg_2_ ( .D(N3081), .CK(clk), .Q(read_counter[2]) );
  DFFHQX1 read_counter_reg_0_ ( .D(N3079), .CK(clk), .Q(read_counter[0]) );
  DFFHQX1 Kt_reg_31_ ( .D(N2977), .CK(clk), .Q(Kt[31]) );
  DFFHQX1 Kt_reg_30_ ( .D(N2976), .CK(clk), .Q(Kt[30]) );
  DFFHQX1 Kt_reg_29_ ( .D(N2975), .CK(clk), .Q(Kt[29]) );
  DFFHQX1 Kt_reg_28_ ( .D(N2974), .CK(clk), .Q(Kt[28]) );
  DFFHQX1 Kt_reg_27_ ( .D(N2973), .CK(clk), .Q(Kt[27]) );
  DFFHQX1 Kt_reg_26_ ( .D(N2972), .CK(clk), .Q(Kt[26]) );
  DFFHQX1 Kt_reg_25_ ( .D(N2971), .CK(clk), .Q(Kt[25]) );
  DFFHQX1 Kt_reg_24_ ( .D(N2970), .CK(clk), .Q(Kt[24]) );
  DFFHQX1 Kt_reg_23_ ( .D(N2969), .CK(clk), .Q(Kt[23]) );
  DFFHQX1 H_reg_16_ ( .D(n2463), .CK(clk), .Q(SHA256_result[16]) );
  DFFHQX1 C_reg_10_ ( .D(n2788), .CK(clk), .Q(SHA256_result[170]) );
  DFFHQX1 B_reg_12_ ( .D(n2819), .CK(clk), .Q(SHA256_result[204]) );
  DFFHQX1 B_reg_14_ ( .D(n2817), .CK(clk), .Q(SHA256_result[206]) );
  DFFHQX1 C_reg_11_ ( .D(n2787), .CK(clk), .Q(SHA256_result[171]) );
  DFFHQX1 A_reg_6_ ( .D(n2889), .CK(clk), .Q(SHA256_result[230]) );
  DFFHQX1 A_reg_7_ ( .D(n2888), .CK(clk), .Q(SHA256_result[231]) );
  DFFHQX1 A_reg_16_ ( .D(n2879), .CK(clk), .Q(SHA256_result[240]) );
  DFFHQX1 A_reg_25_ ( .D(n2870), .CK(clk), .Q(SHA256_result[249]) );
  DFFHQXL A_reg_26_ ( .D(n2869), .CK(clk), .Q(SHA256_result[250]) );
  DFFHQXL A_reg_27_ ( .D(n2868), .CK(clk), .Q(SHA256_result[251]) );
  DFFHQXL A_reg_29_ ( .D(n2866), .CK(clk), .Q(SHA256_result[253]) );
  DFFHQXL A_reg_30_ ( .D(n2865), .CK(clk), .Q(SHA256_result[254]) );
  DFFHQX1 Kt_reg_22_ ( .D(N2968), .CK(clk), .Q(Kt[22]) );
  DFFHQX1 Kt_reg_21_ ( .D(N2967), .CK(clk), .Q(Kt[21]) );
  DFFHQX1 Kt_reg_20_ ( .D(N2966), .CK(clk), .Q(Kt[20]) );
  DFFHQX1 H_reg_14_ ( .D(n2465), .CK(clk), .Q(SHA256_result[14]) );
  DFFHQX1 H_reg_15_ ( .D(n2464), .CK(clk), .Q(SHA256_result[15]) );
  DFFHQX1 H_reg_17_ ( .D(n2462), .CK(clk), .Q(SHA256_result[17]) );
  DFFHQX1 F_reg_19_ ( .D(n2683), .CK(clk), .Q(SHA256_result[83]) );
  DFFHQX1 G_reg_16_ ( .D(n2495), .CK(clk), .Q(SHA256_result[48]) );
  DFFHQX1 G_reg_17_ ( .D(n2494), .CK(clk), .Q(SHA256_result[49]) );
  DFFHQX1 C_reg_5_ ( .D(n2793), .CK(clk), .Q(SHA256_result[165]) );
  DFFHQX1 B_reg_5_ ( .D(n2826), .CK(clk), .Q(SHA256_result[197]) );
  DFFHQX1 B_reg_6_ ( .D(n2825), .CK(clk), .Q(SHA256_result[198]) );
  DFFHQX1 B_reg_8_ ( .D(n2823), .CK(clk), .Q(SHA256_result[200]) );
  DFFX1 F_reg_17_ ( .D(n2685), .CK(clk), .Q(SHA256_result[81]), .QN(n1151) );
  DFFHQX1 C_reg_6_ ( .D(n2792), .CK(clk), .Q(SHA256_result[166]) );
  DFFHQX1 C_reg_7_ ( .D(n2791), .CK(clk), .Q(SHA256_result[167]) );
  DFFHQX1 E_reg_24_ ( .D(n2710), .CK(clk), .Q(SHA256_result[120]) );
  DFFHQX1 A_reg_3_ ( .D(n2892), .CK(clk), .Q(SHA256_result[227]) );
  DFFHQX1 A_reg_4_ ( .D(n2891), .CK(clk), .Q(SHA256_result[228]) );
  DFFHQX1 A_reg_5_ ( .D(n2890), .CK(clk), .Q(SHA256_result[229]) );
  DFFHQX1 Kt_reg_19_ ( .D(N2965), .CK(clk), .Q(Kt[19]) );
  DFFHQX1 Kt_reg_18_ ( .D(N2964), .CK(clk), .Q(Kt[18]) );
  DFFHQX1 Kt_reg_17_ ( .D(N2963), .CK(clk), .Q(Kt[17]) );
  DFFHQX1 Kt_reg_16_ ( .D(N2962), .CK(clk), .Q(Kt[16]) );
  DFFHQX1 H3_reg_2_ ( .D(n2604), .CK(clk), .Q(H3[2]) );
  DFFHQX1 H7_reg_2_ ( .D(n2445), .CK(clk), .Q(H7[2]) );
  DFFHQX1 H2_reg_2_ ( .D(n2573), .CK(clk), .Q(H2[2]) );
  DFFHQX1 H6_reg_2_ ( .D(n2540), .CK(clk), .Q(H6[2]) );
  DFFHQX1 H6_reg_3_ ( .D(n2539), .CK(clk), .Q(H6[3]) );
  DFFHQX1 H_reg_3_ ( .D(n2476), .CK(clk), .Q(SHA256_result[3]) );
  DFFHQX1 H_reg_4_ ( .D(n2475), .CK(clk), .Q(SHA256_result[4]) );
  DFFHQX1 H_reg_6_ ( .D(n2473), .CK(clk), .Q(SHA256_result[6]) );
  DFFHQX1 H_reg_7_ ( .D(n2472), .CK(clk), .Q(SHA256_result[7]) );
  DFFHQX1 H_reg_8_ ( .D(n2471), .CK(clk), .Q(SHA256_result[8]) );
  DFFHQX1 H_reg_9_ ( .D(n2470), .CK(clk), .Q(SHA256_result[9]) );
  DFFHQX1 H_reg_10_ ( .D(n2469), .CK(clk), .Q(SHA256_result[10]) );
  DFFHQX1 C_reg_4_ ( .D(n2794), .CK(clk), .Q(SHA256_result[164]) );
  DFFHQX1 E_reg_18_ ( .D(n2716), .CK(clk), .Q(SHA256_result[114]) );
  DFFHQX1 E_reg_23_ ( .D(n2711), .CK(clk), .Q(SHA256_result[119]) );
  DFFHQX1 digest_reg_31_ ( .D(N3078), .CK(clk), .Q(digest[31]) );
  DFFHQX1 digest_reg_30_ ( .D(N3077), .CK(clk), .Q(digest[30]) );
  DFFHQX1 digest_reg_29_ ( .D(N3076), .CK(clk), .Q(digest[29]) );
  DFFHQX1 digest_reg_28_ ( .D(N3075), .CK(clk), .Q(digest[28]) );
  DFFHQX1 digest_reg_27_ ( .D(N3074), .CK(clk), .Q(digest[27]) );
  DFFHQX1 digest_reg_26_ ( .D(N3073), .CK(clk), .Q(digest[26]) );
  DFFHQX1 digest_reg_25_ ( .D(N3072), .CK(clk), .Q(digest[25]) );
  DFFHQX1 digest_reg_24_ ( .D(N3071), .CK(clk), .Q(digest[24]) );
  DFFHQX1 digest_reg_23_ ( .D(N3070), .CK(clk), .Q(digest[23]) );
  DFFHQX1 digest_reg_22_ ( .D(N3069), .CK(clk), .Q(digest[22]) );
  DFFHQX1 digest_reg_21_ ( .D(N3068), .CK(clk), .Q(digest[21]) );
  DFFHQX1 digest_reg_20_ ( .D(N3067), .CK(clk), .Q(digest[20]) );
  DFFHQX1 digest_reg_19_ ( .D(N3066), .CK(clk), .Q(digest[19]) );
  DFFHQX1 digest_reg_18_ ( .D(N3065), .CK(clk), .Q(digest[18]) );
  DFFHQX1 digest_reg_17_ ( .D(N3064), .CK(clk), .Q(digest[17]) );
  DFFHQX1 digest_reg_16_ ( .D(N3063), .CK(clk), .Q(digest[16]) );
  DFFHQX1 digest_reg_15_ ( .D(N3062), .CK(clk), .Q(digest[15]) );
  DFFHQX1 digest_reg_14_ ( .D(N3061), .CK(clk), .Q(digest[14]) );
  DFFHQX1 digest_reg_13_ ( .D(N3060), .CK(clk), .Q(digest[13]) );
  DFFHQX1 digest_reg_12_ ( .D(N3059), .CK(clk), .Q(digest[12]) );
  DFFHQX1 digest_reg_11_ ( .D(N3058), .CK(clk), .Q(digest[11]) );
  DFFHQX1 digest_reg_10_ ( .D(N3057), .CK(clk), .Q(digest[10]) );
  DFFHQX1 digest_reg_9_ ( .D(N3056), .CK(clk), .Q(digest[9]) );
  DFFHQX1 digest_reg_8_ ( .D(N3055), .CK(clk), .Q(digest[8]) );
  DFFHQX1 digest_reg_7_ ( .D(N3054), .CK(clk), .Q(digest[7]) );
  DFFHQX1 digest_reg_6_ ( .D(N3053), .CK(clk), .Q(digest[6]) );
  DFFHQX1 digest_reg_5_ ( .D(N3052), .CK(clk), .Q(digest[5]) );
  DFFHQX1 digest_reg_4_ ( .D(N3051), .CK(clk), .Q(digest[4]) );
  DFFHQX1 digest_reg_3_ ( .D(N3050), .CK(clk), .Q(digest[3]) );
  DFFHQX1 digest_reg_2_ ( .D(N3049), .CK(clk), .Q(digest[2]) );
  DFFHQX1 digest_reg_1_ ( .D(N3048), .CK(clk), .Q(digest[1]) );
  DFFHQX1 digest_reg_0_ ( .D(N3047), .CK(clk), .Q(digest[0]) );
  DFFHQX4 C_reg_1_ ( .D(n2797), .CK(clk), .Q(SHA256_result[161]) );
  DFFHQXL H3_reg_31_ ( .D(n2575), .CK(clk), .Q(H3[31]) );
  DFFHQXL C_reg_31_ ( .D(n2767), .CK(clk), .Q(SHA256_result[191]) );
  DFFHQXL D_reg_31_ ( .D(n2735), .CK(clk), .Q(SHA256_result[159]) );
  DFFHQX4 A_reg_0_ ( .D(n2895), .CK(clk), .Q(SHA256_result[224]) );
  DFFHQXL H1_reg_31_ ( .D(n2832), .CK(clk), .Q(H1[31]) );
  DFFHQXL B_reg_31_ ( .D(n2800), .CK(clk), .Q(SHA256_result[223]) );
  DFFHQXL G_reg_31_ ( .D(n2480), .CK(clk), .Q(SHA256_result[63]) );
  DFFHQXL H2_reg_11_ ( .D(n2564), .CK(clk), .Q(H2[11]) );
  DFFHQXL H3_reg_11_ ( .D(n2595), .CK(clk), .Q(H3[11]) );
  DFFHQXL H5_reg_9_ ( .D(n2661), .CK(clk), .Q(H5[9]) );
  DFFHQXL H2_reg_10_ ( .D(n2565), .CK(clk), .Q(H2[10]) );
  DFFHQXL H5_reg_10_ ( .D(n2660), .CK(clk), .Q(H5[10]) );
  DFFHQXL G_reg_23_ ( .D(n2488), .CK(clk), .Q(SHA256_result[55]) );
  DFFHQXL D_reg_0_ ( .D(n2766), .CK(clk), .Q(SHA256_result[128]) );
  DFFHQXL D_reg_2_ ( .D(n2764), .CK(clk), .Q(SHA256_result[130]) );
  DFFHQXL H_reg_21_ ( .D(n2458), .CK(clk), .Q(SHA256_result[21]) );
  DFFXL F_reg_23_ ( .D(n2679), .CK(clk), .Q(SHA256_result[87]), .QN(n1145) );
  DFFHQXL A_reg_21_ ( .D(n2874), .CK(clk), .Q(SHA256_result[245]) );
  DFFHQXL A_reg_10_ ( .D(n2885), .CK(clk), .Q(SHA256_result[234]) );
  DFFHQXL A_reg_12_ ( .D(n2883), .CK(clk), .Q(SHA256_result[236]) );
  DFFHQXL A_reg_11_ ( .D(n2884), .CK(clk), .Q(SHA256_result[235]) );
  DFFHQXL A_reg_9_ ( .D(n2886), .CK(clk), .Q(SHA256_result[233]) );
  DFFHQXL A_reg_20_ ( .D(n2875), .CK(clk), .Q(SHA256_result[244]) );
  DFFHQXL A_reg_8_ ( .D(n2887), .CK(clk), .Q(SHA256_result[232]) );
  DFFHQXL H3_reg_9_ ( .D(n2597), .CK(clk), .Q(H3[9]) );
  DFFHQXL H1_reg_8_ ( .D(n2855), .CK(clk), .Q(H1[8]) );
  DFFHQXL H7_reg_7_ ( .D(n2440), .CK(clk), .Q(H7[7]) );
  DFFHQXL H2_reg_7_ ( .D(n2568), .CK(clk), .Q(H2[7]) );
  DFFHQXL H2_reg_9_ ( .D(n2566), .CK(clk), .Q(H2[9]) );
  DFFHQXL H3_reg_8_ ( .D(n2598), .CK(clk), .Q(H3[8]) );
  DFFHQXL H5_reg_6_ ( .D(n2664), .CK(clk), .Q(H5[6]) );
  DFFXL F_reg_16_ ( .D(n2686), .CK(clk), .Q(SHA256_result[80]), .QN(n1152) );
  DFFHQXL A_reg_18_ ( .D(n2877), .CK(clk), .Q(SHA256_result[242]) );
  DFFHQXL A_reg_17_ ( .D(n2878), .CK(clk), .Q(SHA256_result[241]) );
  DFFHQXL A_reg_19_ ( .D(n2876), .CK(clk), .Q(SHA256_result[243]) );
  DFFHQXL A_reg_24_ ( .D(n2871), .CK(clk), .Q(SHA256_result[248]) );
  DFFHQXL A_reg_15_ ( .D(n2880), .CK(clk), .Q(SHA256_result[239]) );
  DFFHQXL A_reg_13_ ( .D(n2882), .CK(clk), .Q(SHA256_result[237]) );
  DFFHQXL H5_reg_5_ ( .D(n2665), .CK(clk), .Q(H5[5]) );
  DFFHQXL H3_reg_6_ ( .D(n2600), .CK(clk), .Q(H3[6]) );
  DFFHQXL H1_reg_6_ ( .D(n2857), .CK(clk), .Q(H1[6]) );
  DFFHQXL H2_reg_6_ ( .D(n2569), .CK(clk), .Q(H2[6]) );
  DFFHQXL H2_reg_5_ ( .D(n2570), .CK(clk), .Q(H2[5]) );
  DFFHQXL H3_reg_5_ ( .D(n2601), .CK(clk), .Q(H3[5]) );
  DFFHQXL H5_reg_3_ ( .D(n2667), .CK(clk), .Q(H5[3]) );
  DFFHQXL H_reg_11_ ( .D(n2468), .CK(clk), .Q(SHA256_result[11]) );
  DFFHQXL A_reg_14_ ( .D(n2881), .CK(clk), .Q(SHA256_result[238]) );
  DFFHQXL H1_reg_4_ ( .D(n2859), .CK(clk), .Q(H1[4]) );
  DFFHQXL H2_reg_4_ ( .D(n2571), .CK(clk), .Q(H2[4]) );
  DFFHQXL H3_reg_4_ ( .D(n2602), .CK(clk), .Q(H3[4]) );
  DFFHQXL H2_reg_3_ ( .D(n2572), .CK(clk), .Q(H2[3]) );
  DFFHQXL H4_reg_23_ ( .D(n2615), .CK(clk), .Q(H4[23]) );
  DFFHQX1 F_reg_20_ ( .D(n2682), .CK(clk), .Q(SHA256_result[84]) );
  DFFHQX1 H_reg_18_ ( .D(n2461), .CK(clk), .Q(SHA256_result[18]) );
  DFFHQX1 H_reg_19_ ( .D(n2460), .CK(clk), .Q(SHA256_result[19]) );
  DFFHQX1 H1_reg_5_ ( .D(n2858), .CK(clk), .Q(H1[5]) );
  DFFHQX1 H7_reg_4_ ( .D(n2443), .CK(clk), .Q(H7[4]) );
  DFFX1 F_reg_7_ ( .D(n2695), .CK(clk), .Q(SHA256_result[71]), .QN(n1161) );
  DFFHQX1 H1_reg_3_ ( .D(n2860), .CK(clk), .Q(H1[3]) );
  DFFHQX1 H3_reg_3_ ( .D(n2603), .CK(clk), .Q(H3[3]) );
  DFFHQX1 H5_reg_2_ ( .D(n2668), .CK(clk), .Q(H5[2]) );
  DFFHQX1 H7_reg_3_ ( .D(n2444), .CK(clk), .Q(H7[3]) );
  DFFHQX1 C_reg_8_ ( .D(n2790), .CK(clk), .Q(SHA256_result[168]) );
  DFFHQX1 C_reg_12_ ( .D(n2786), .CK(clk), .Q(SHA256_result[172]) );
  DFFHQX1 B_reg_9_ ( .D(n2822), .CK(clk), .Q(SHA256_result[201]) );
  DFFHQX1 B_reg_13_ ( .D(n2818), .CK(clk), .Q(SHA256_result[205]) );
  DFFHQX1 B_reg_10_ ( .D(n2821), .CK(clk), .Q(SHA256_result[202]) );
  DFFHQX1 B_reg_11_ ( .D(n2820), .CK(clk), .Q(SHA256_result[203]) );
  DFFHQXL C_reg_30_ ( .D(n2768), .CK(clk), .Q(SHA256_result[190]) );
  DFFHQXL D_reg_30_ ( .D(n2736), .CK(clk), .Q(SHA256_result[158]) );
  DFFHQXL B_reg_30_ ( .D(n2801), .CK(clk), .Q(SHA256_result[222]) );
  DFFHQX1 H2_reg_18_ ( .D(n2557), .CK(clk), .Q(H2[18]) );
  DFFHQX1 B_reg_18_ ( .D(n2813), .CK(clk), .Q(SHA256_result[210]) );
  DFFHQXL H0_reg_31_ ( .D(n2896), .CK(clk), .Q(H0[31]) );
  DFFHQXL H1_reg_30_ ( .D(n2833), .CK(clk), .Q(H1[30]) );
  DFFHQXL H6_reg_30_ ( .D(n2512), .CK(clk), .Q(H6[30]) );
  DFFHQXL H2_reg_30_ ( .D(n2545), .CK(clk), .Q(H2[30]) );
  DFFHQXL H3_reg_30_ ( .D(n2576), .CK(clk), .Q(H3[30]) );
  DFFHQXL H4_reg_31_ ( .D(n2607), .CK(clk), .Q(H4[31]) );
  DFFHQXL H5_reg_30_ ( .D(n2640), .CK(clk), .Q(H5[30]) );
  DFFHQXL H7_reg_30_ ( .D(n2417), .CK(clk), .Q(H7[30]) );
  DFFHQXL H6_reg_31_ ( .D(n2511), .CK(clk), .Q(H6[31]) );
  DFFHQXL H2_reg_31_ ( .D(n2544), .CK(clk), .Q(H2[31]) );
  DFFHQXL H7_reg_31_ ( .D(n2416), .CK(clk), .Q(H7[31]) );
  DFFHQXL H5_reg_31_ ( .D(n2639), .CK(clk), .Q(H5[31]) );
  DFFHQXL H4_reg_28_ ( .D(n2610), .CK(clk), .Q(H4[28]) );
  DFFHQXL H0_reg_28_ ( .D(n2899), .CK(clk), .Q(H0[28]) );
  DFFHQXL H0_reg_29_ ( .D(n2898), .CK(clk), .Q(H0[29]) );
  DFFHQXL H4_reg_29_ ( .D(n2609), .CK(clk), .Q(H4[29]) );
  DFFHQXL H0_reg_30_ ( .D(n2897), .CK(clk), .Q(H0[30]) );
  DFFHQXL H3_reg_27_ ( .D(n2579), .CK(clk), .Q(H3[27]) );
  DFFHQXL H6_reg_28_ ( .D(n2514), .CK(clk), .Q(H6[28]) );
  DFFHQXL H1_reg_27_ ( .D(n2836), .CK(clk), .Q(H1[27]) );
  DFFHQXL H1_reg_29_ ( .D(n2834), .CK(clk), .Q(H1[29]) );
  DFFHQXL H2_reg_28_ ( .D(n2547), .CK(clk), .Q(H2[28]) );
  DFFHQXL H3_reg_29_ ( .D(n2577), .CK(clk), .Q(H3[29]) );
  DFFHQXL H5_reg_28_ ( .D(n2642), .CK(clk), .Q(H5[28]) );
  DFFHQXL H7_reg_27_ ( .D(n2420), .CK(clk), .Q(H7[27]) );
  DFFHQXL H7_reg_28_ ( .D(n2419), .CK(clk), .Q(H7[28]) );
  DFFHQXL H3_reg_28_ ( .D(n2578), .CK(clk), .Q(H3[28]) );
  DFFHQXL H6_reg_29_ ( .D(n2513), .CK(clk), .Q(H6[29]) );
  DFFHQXL H7_reg_29_ ( .D(n2418), .CK(clk), .Q(H7[29]) );
  DFFHQXL H5_reg_29_ ( .D(n2641), .CK(clk), .Q(H5[29]) );
  DFFHQXL H2_reg_27_ ( .D(n2548), .CK(clk), .Q(H2[27]) );
  DFFHQXL H2_reg_29_ ( .D(n2546), .CK(clk), .Q(H2[29]) );
  DFFHQXL H0_reg_21_ ( .D(n2906), .CK(clk), .Q(H0[21]) );
  DFFHQXL H0_reg_23_ ( .D(n2904), .CK(clk), .Q(H0[23]) );
  DFFHQXL H0_reg_27_ ( .D(n2900), .CK(clk), .Q(H0[27]) );
  DFFHQXL H4_reg_22_ ( .D(n2616), .CK(clk), .Q(H4[22]) );
  DFFHQXL H0_reg_22_ ( .D(n2905), .CK(clk), .Q(H0[22]) );
  DFFHQXL H4_reg_27_ ( .D(n2611), .CK(clk), .Q(H4[27]) );
  DFFHQXL H4_reg_20_ ( .D(n2618), .CK(clk), .Q(H4[20]) );
  DFFHQXL H0_reg_20_ ( .D(n2907), .CK(clk), .Q(H0[20]) );
  DFFHQXL H0_reg_26_ ( .D(n2901), .CK(clk), .Q(H0[26]) );
  DFFHQXL H4_reg_26_ ( .D(n2612), .CK(clk), .Q(H4[26]) );
  DFFHQXL H0_reg_24_ ( .D(n2903), .CK(clk), .Q(H0[24]) );
  DFFHQXL H0_reg_25_ ( .D(n2902), .CK(clk), .Q(H0[25]) );
  DFFHQXL H4_reg_24_ ( .D(n2614), .CK(clk), .Q(H4[24]) );
  DFFHQXL H4_reg_25_ ( .D(n2613), .CK(clk), .Q(H4[25]) );
  DFFHQXL H4_reg_30_ ( .D(n2608), .CK(clk), .Q(H4[30]) );
  DFFHQXL H2_reg_24_ ( .D(n2551), .CK(clk), .Q(H2[24]) );
  DFFHQXL H5_reg_26_ ( .D(n2644), .CK(clk), .Q(H5[26]) );
  DFFHQXL H1_reg_24_ ( .D(n2839), .CK(clk), .Q(H1[24]) );
  DFFHQXL H1_reg_25_ ( .D(n2838), .CK(clk), .Q(H1[25]) );
  DFFHQXL H2_reg_26_ ( .D(n2549), .CK(clk), .Q(H2[26]) );
  DFFHQXL H3_reg_24_ ( .D(n2582), .CK(clk), .Q(H3[24]) );
  DFFHQXL H3_reg_26_ ( .D(n2580), .CK(clk), .Q(H3[26]) );
  DFFHQXL H5_reg_25_ ( .D(n2645), .CK(clk), .Q(H5[25]) );
  DFFHQXL H5_reg_27_ ( .D(n2643), .CK(clk), .Q(H5[27]) );
  DFFHQXL H6_reg_24_ ( .D(n2518), .CK(clk), .Q(H6[24]) );
  DFFHQXL H6_reg_26_ ( .D(n2516), .CK(clk), .Q(H6[26]) );
  DFFHQXL H7_reg_25_ ( .D(n2422), .CK(clk), .Q(H7[25]) );
  DFFHQXL H1_reg_26_ ( .D(n2837), .CK(clk), .Q(H1[26]) );
  DFFHQXL H2_reg_25_ ( .D(n2550), .CK(clk), .Q(H2[25]) );
  DFFHQXL H3_reg_25_ ( .D(n2581), .CK(clk), .Q(H3[25]) );
  DFFHQXL H7_reg_26_ ( .D(n2421), .CK(clk), .Q(H7[26]) );
  DFFHQXL H4_reg_15_ ( .D(n2623), .CK(clk), .Q(H4[15]) );
  DFFHQXL H0_reg_17_ ( .D(n2910), .CK(clk), .Q(H0[17]) );
  DFFHQXL H4_reg_21_ ( .D(n2617), .CK(clk), .Q(H4[21]) );
  DFFHQXL H0_reg_18_ ( .D(n2909), .CK(clk), .Q(H0[18]) );
  DFFHQXL H0_reg_15_ ( .D(n2912), .CK(clk), .Q(H0[15]) );
  DFFHQXL H0_reg_19_ ( .D(n2908), .CK(clk), .Q(H0[19]) );
  DFFHQXL H4_reg_17_ ( .D(n2621), .CK(clk), .Q(H4[17]) );
  DFFHQXL H4_reg_19_ ( .D(n2619), .CK(clk), .Q(H4[19]) );
  DFFHQXL H4_reg_12_ ( .D(n2626), .CK(clk), .Q(H4[12]) );
  DFFHQXL H0_reg_11_ ( .D(n2916), .CK(clk), .Q(H0[11]) );
  DFFHQXL H0_reg_10_ ( .D(n2917), .CK(clk), .Q(H0[10]) );
  DFFHQXL H4_reg_14_ ( .D(n2624), .CK(clk), .Q(H4[14]) );
  DFFHQXL H4_reg_18_ ( .D(n2620), .CK(clk), .Q(H4[18]) );
  DFFHQXL H0_reg_14_ ( .D(n2913), .CK(clk), .Q(H0[14]) );
  DFFHQXL H0_reg_13_ ( .D(n2914), .CK(clk), .Q(H0[13]) );
  DFFHQXL H_reg_31_ ( .D(n2448), .CK(clk), .Q(SHA256_result[31]) );
  DFFHQXL H4_reg_16_ ( .D(n2622), .CK(clk), .Q(H4[16]) );
  DFFHQXL H0_reg_12_ ( .D(n2915), .CK(clk), .Q(H0[12]) );
  DFFHQXL H0_reg_16_ ( .D(n2911), .CK(clk), .Q(H0[16]) );
  DFFHQXL H4_reg_13_ ( .D(n2625), .CK(clk), .Q(H4[13]) );
  DFFHQXL D_reg_29_ ( .D(n2737), .CK(clk), .Q(SHA256_result[157]) );
  DFFHQXL D_reg_25_ ( .D(n2741), .CK(clk), .Q(SHA256_result[153]) );
  DFFHQXL D_reg_28_ ( .D(n2738), .CK(clk), .Q(SHA256_result[156]) );
  DFFHQXL D_reg_26_ ( .D(n2740), .CK(clk), .Q(SHA256_result[154]) );
  DFFHQXL D_reg_27_ ( .D(n2739), .CK(clk), .Q(SHA256_result[155]) );
  DFFHQXL H6_reg_22_ ( .D(n2520), .CK(clk), .Q(H6[22]) );
  DFFHQXL H5_reg_23_ ( .D(n2647), .CK(clk), .Q(H5[23]) );
  DFFHQXL H2_reg_22_ ( .D(n2553), .CK(clk), .Q(H2[22]) );
  DFFHQXL H3_reg_22_ ( .D(n2584), .CK(clk), .Q(H3[22]) );
  DFFHQXL H5_reg_24_ ( .D(n2646), .CK(clk), .Q(H5[24]) );
  DFFHQXL H6_reg_23_ ( .D(n2519), .CK(clk), .Q(H6[23]) );
  DFFHQXL H7_reg_23_ ( .D(n2424), .CK(clk), .Q(H7[23]) );
  DFFHQXL H1_reg_22_ ( .D(n2841), .CK(clk), .Q(H1[22]) );
  DFFHQXL H7_reg_22_ ( .D(n2425), .CK(clk), .Q(H7[22]) );
  DFFHQXL H2_reg_23_ ( .D(n2552), .CK(clk), .Q(H2[23]) );
  DFFHQXL H3_reg_21_ ( .D(n2585), .CK(clk), .Q(H3[21]) );
  DFFHQXL H3_reg_23_ ( .D(n2583), .CK(clk), .Q(H3[23]) );
  DFFHQXL H5_reg_22_ ( .D(n2648), .CK(clk), .Q(H5[22]) );
  DFFHQXL H4_reg_7_ ( .D(n2631), .CK(clk), .Q(H4[7]) );
  DFFHQXL H4_reg_4_ ( .D(n2634), .CK(clk), .Q(H4[4]) );
  DFFHQXL H0_reg_4_ ( .D(n2923), .CK(clk), .Q(H0[4]) );
  DFFHQXL H4_reg_3_ ( .D(n2635), .CK(clk), .Q(H4[3]) );
  DFFHQXL H4_reg_5_ ( .D(n2633), .CK(clk), .Q(H4[5]) );
  DFFHQXL H0_reg_3_ ( .D(n2924), .CK(clk), .Q(H0[3]) );
  DFFHQXL H4_reg_8_ ( .D(n2630), .CK(clk), .Q(H4[8]) );
  DFFHQXL H4_reg_6_ ( .D(n2632), .CK(clk), .Q(H4[6]) );
  DFFHQXL H0_reg_6_ ( .D(n2921), .CK(clk), .Q(H0[6]) );
  DFFHQXL H0_reg_7_ ( .D(n2920), .CK(clk), .Q(H0[7]) );
  DFFHQXL H0_reg_8_ ( .D(n2919), .CK(clk), .Q(H0[8]) );
  DFFHQXL H4_reg_9_ ( .D(n2629), .CK(clk), .Q(H4[9]) );
  DFFHQXL H0_reg_2_ ( .D(n2925), .CK(clk), .Q(H0[2]) );
  DFFHQXL H4_reg_2_ ( .D(n2636), .CK(clk), .Q(H4[2]) );
  DFFHQXL H4_reg_10_ ( .D(n2628), .CK(clk), .Q(H4[10]) );
  DFFHQXL H4_reg_11_ ( .D(n2627), .CK(clk), .Q(H4[11]) );
  DFFHQXL H0_reg_9_ ( .D(n2918), .CK(clk), .Q(H0[9]) );
  DFFHQXL D_reg_18_ ( .D(n2748), .CK(clk), .Q(SHA256_result[146]) );
  DFFHQXL D_reg_19_ ( .D(n2747), .CK(clk), .Q(SHA256_result[147]) );
  DFFHQXL D_reg_23_ ( .D(n2743), .CK(clk), .Q(SHA256_result[151]) );
  DFFHQXL D_reg_22_ ( .D(n2744), .CK(clk), .Q(SHA256_result[150]) );
  DFFHQXL D_reg_21_ ( .D(n2745), .CK(clk), .Q(SHA256_result[149]) );
  DFFHQXL D_reg_20_ ( .D(n2746), .CK(clk), .Q(SHA256_result[148]) );
  DFFHQXL D_reg_24_ ( .D(n2742), .CK(clk), .Q(SHA256_result[152]) );
  DFFHQXL H1_reg_20_ ( .D(n2843), .CK(clk), .Q(H1[20]) );
  DFFHQXL H3_reg_20_ ( .D(n2586), .CK(clk), .Q(H3[20]) );
  DFFHQXL H6_reg_19_ ( .D(n2523), .CK(clk), .Q(H6[19]) );
  DFFHQXL H5_reg_21_ ( .D(n2649), .CK(clk), .Q(H5[21]) );
  DFFHQXL H6_reg_21_ ( .D(n2521), .CK(clk), .Q(H6[21]) );
  DFFHQXL H2_reg_21_ ( .D(n2554), .CK(clk), .Q(H2[21]) );
  DFFHQXL H2_reg_19_ ( .D(n2556), .CK(clk), .Q(H2[19]) );
  DFFHQXL H7_reg_21_ ( .D(n2426), .CK(clk), .Q(H7[21]) );
  DFFHQXL H1_reg_19_ ( .D(n2844), .CK(clk), .Q(H1[19]) );
  DFFHQXL H2_reg_20_ ( .D(n2555), .CK(clk), .Q(H2[20]) );
  DFFHQXL H5_reg_20_ ( .D(n2650), .CK(clk), .Q(H5[20]) );
  DFFHQXL H6_reg_20_ ( .D(n2522), .CK(clk), .Q(H6[20]) );
  DFFHQXL H1_reg_21_ ( .D(n2842), .CK(clk), .Q(H1[21]) );
  DFFHQXL H3_reg_19_ ( .D(n2587), .CK(clk), .Q(H3[19]) );
  DFFHQXL H0_reg_0_ ( .D(n2927), .CK(clk), .Q(H0[0]) );
  DFFHQXL H4_reg_0_ ( .D(n2638), .CK(clk), .Q(H4[0]) );
  DFFHQXL H4_reg_1_ ( .D(n2637), .CK(clk), .Q(H4[1]) );
  DFFHQXL H_reg_28_ ( .D(n2451), .CK(clk), .Q(SHA256_result[28]) );
  DFFHQXL H_reg_30_ ( .D(n2449), .CK(clk), .Q(SHA256_result[30]) );
  DFFHQXL H_reg_29_ ( .D(n2450), .CK(clk), .Q(SHA256_result[29]) );
  DFFHQXL D_reg_17_ ( .D(n2749), .CK(clk), .Q(SHA256_result[145]) );
  DFFHQXL C_reg_29_ ( .D(n2769), .CK(clk), .Q(SHA256_result[189]) );
  DFFHQXL F_reg_30_ ( .D(n2672), .CK(clk), .Q(SHA256_result[94]) );
  DFFHQXL G_reg_30_ ( .D(n2481), .CK(clk), .Q(SHA256_result[62]) );
  DFFHQXL D_reg_10_ ( .D(n2756), .CK(clk), .Q(SHA256_result[138]) );
  DFFHQXL D_reg_16_ ( .D(n2750), .CK(clk), .Q(SHA256_result[144]) );
  DFFHQXL D_reg_14_ ( .D(n2752), .CK(clk), .Q(SHA256_result[142]) );
  DFFHQXL D_reg_15_ ( .D(n2751), .CK(clk), .Q(SHA256_result[143]) );
  DFFHQXL B_reg_29_ ( .D(n2802), .CK(clk), .Q(SHA256_result[221]) );
  DFFHQXL D_reg_12_ ( .D(n2754), .CK(clk), .Q(SHA256_result[140]) );
  DFFHQXL D_reg_11_ ( .D(n2755), .CK(clk), .Q(SHA256_result[139]) );
  DFFHQXL B_reg_28_ ( .D(n2803), .CK(clk), .Q(SHA256_result[220]) );
  DFFHQXL C_reg_28_ ( .D(n2770), .CK(clk), .Q(SHA256_result[188]) );
  DFFHQXL D_reg_13_ ( .D(n2753), .CK(clk), .Q(SHA256_result[141]) );
  DFFHQXL H7_reg_17_ ( .D(n2430), .CK(clk), .Q(H7[17]) );
  DFFHQXL H7_reg_18_ ( .D(n2429), .CK(clk), .Q(H7[18]) );
  DFFHQXL H5_reg_19_ ( .D(n2651), .CK(clk), .Q(H5[19]) );
  DFFHQXL H1_reg_18_ ( .D(n2845), .CK(clk), .Q(H1[18]) );
  DFFHQXL H6_reg_17_ ( .D(n2525), .CK(clk), .Q(H6[17]) );
  DFFHQXL H3_reg_17_ ( .D(n2589), .CK(clk), .Q(H3[17]) );
  DFFHQXL H3_reg_18_ ( .D(n2588), .CK(clk), .Q(H3[18]) );
  DFFHQXL H5_reg_18_ ( .D(n2652), .CK(clk), .Q(H5[18]) );
  DFFHQXL H2_reg_17_ ( .D(n2558), .CK(clk), .Q(H2[17]) );
  DFFHQXL H7_reg_19_ ( .D(n2428), .CK(clk), .Q(H7[19]) );
  DFFHQXL G_reg_28_ ( .D(n2483), .CK(clk), .Q(SHA256_result[60]) );
  DFFHQXL D_reg_7_ ( .D(n2759), .CK(clk), .Q(SHA256_result[135]) );
  DFFHQXL D_reg_8_ ( .D(n2758), .CK(clk), .Q(SHA256_result[136]) );
  DFFHQXL D_reg_9_ ( .D(n2757), .CK(clk), .Q(SHA256_result[137]) );
  DFFHQXL F_reg_29_ ( .D(n2673), .CK(clk), .Q(SHA256_result[93]) );
  DFFHQXL C_reg_26_ ( .D(n2772), .CK(clk), .Q(SHA256_result[186]) );
  DFFHQXL C_reg_24_ ( .D(n2774), .CK(clk), .Q(SHA256_result[184]) );
  DFFXL F_reg_28_ ( .D(n2674), .CK(clk), .Q(SHA256_result[92]), .QN(n1140) );
  DFFHQXL B_reg_27_ ( .D(n2804), .CK(clk), .Q(SHA256_result[219]) );
  DFFHQXL B_reg_26_ ( .D(n2805), .CK(clk), .Q(SHA256_result[218]) );
  DFFHQXL C_reg_25_ ( .D(n2773), .CK(clk), .Q(SHA256_result[185]) );
  DFFHQXL G_reg_29_ ( .D(n2482), .CK(clk), .Q(SHA256_result[61]) );
  DFFHQXL C_reg_27_ ( .D(n2771), .CK(clk), .Q(SHA256_result[187]) );
  DFFHQXL B_reg_25_ ( .D(n2806), .CK(clk), .Q(SHA256_result[217]) );
  DFFHQXL B_reg_24_ ( .D(n2807), .CK(clk), .Q(SHA256_result[216]) );
  DFFHQXL H7_reg_16_ ( .D(n2431), .CK(clk), .Q(H7[16]) );
  DFFHQXL H5_reg_17_ ( .D(n2653), .CK(clk), .Q(H5[17]) );
  DFFHQXL H1_reg_15_ ( .D(n2848), .CK(clk), .Q(H1[15]) );
  DFFHQXL H1_reg_16_ ( .D(n2847), .CK(clk), .Q(H1[16]) );
  DFFHQXL H6_reg_14_ ( .D(n2528), .CK(clk), .Q(H6[14]) );
  DFFHQXL H6_reg_15_ ( .D(n2527), .CK(clk), .Q(H6[15]) );
  DFFHQXL H6_reg_16_ ( .D(n2526), .CK(clk), .Q(H6[16]) );
  DFFHQXL H7_reg_15_ ( .D(n2432), .CK(clk), .Q(H7[15]) );
  DFFHQXL H2_reg_15_ ( .D(n2560), .CK(clk), .Q(H2[15]) );
  DFFHQXL H3_reg_15_ ( .D(n2591), .CK(clk), .Q(H3[15]) );
  DFFHQXL H3_reg_16_ ( .D(n2590), .CK(clk), .Q(H3[16]) );
  DFFHQXL H1_reg_14_ ( .D(n2849), .CK(clk), .Q(H1[14]) );
  DFFHQXL H5_reg_16_ ( .D(n2654), .CK(clk), .Q(H5[16]) );
  DFFHQXL H_reg_24_ ( .D(n2455), .CK(clk), .Q(SHA256_result[24]) );
  DFFHQXL H_reg_25_ ( .D(n2454), .CK(clk), .Q(SHA256_result[25]) );
  DFFHQXL H_reg_26_ ( .D(n2453), .CK(clk), .Q(SHA256_result[26]) );
  DFFHQXL D_reg_5_ ( .D(n2761), .CK(clk), .Q(SHA256_result[133]) );
  DFFHQXL H_reg_27_ ( .D(n2452), .CK(clk), .Q(SHA256_result[27]) );
  DFFHQXL D_reg_3_ ( .D(n2763), .CK(clk), .Q(SHA256_result[131]) );
  DFFHQXL D_reg_6_ ( .D(n2760), .CK(clk), .Q(SHA256_result[134]) );
  DFFHQXL C_reg_22_ ( .D(n2776), .CK(clk), .Q(SHA256_result[182]) );
  DFFHQXL D_reg_4_ ( .D(n2762), .CK(clk), .Q(SHA256_result[132]) );
  DFFHQXL B_reg_21_ ( .D(n2810), .CK(clk), .Q(SHA256_result[213]) );
  DFFHQXL B_reg_22_ ( .D(n2809), .CK(clk), .Q(SHA256_result[214]) );
  DFFHQXL C_reg_21_ ( .D(n2777), .CK(clk), .Q(SHA256_result[181]) );
  DFFHQXL C_reg_20_ ( .D(n2778), .CK(clk), .Q(SHA256_result[180]) );
  DFFHQXL C_reg_23_ ( .D(n2775), .CK(clk), .Q(SHA256_result[183]) );
  DFFHQXL B_reg_20_ ( .D(n2811), .CK(clk), .Q(SHA256_result[212]) );
  DFFHQXL B_reg_23_ ( .D(n2808), .CK(clk), .Q(SHA256_result[215]) );
  DFFTRX1 round_reg_0_ ( .D(N121), .RN(n129), .CK(clk), .Q(n344), .QN(n1396)
         );
  DFFHQXL H6_reg_13_ ( .D(n2529), .CK(clk), .Q(H6[13]) );
  DFFHQXL H7_reg_12_ ( .D(n2435), .CK(clk), .Q(H7[12]) );
  DFFHQXL H7_reg_13_ ( .D(n2434), .CK(clk), .Q(H7[13]) );
  DFFHQXL H5_reg_15_ ( .D(n2655), .CK(clk), .Q(H5[15]) );
  DFFHQXL H1_reg_11_ ( .D(n2852), .CK(clk), .Q(H1[11]) );
  DFFHQXL H1_reg_13_ ( .D(n2850), .CK(clk), .Q(H1[13]) );
  DFFHQXL H5_reg_13_ ( .D(n2657), .CK(clk), .Q(H5[13]) );
  DFFHQXL H6_reg_12_ ( .D(n2530), .CK(clk), .Q(H6[12]) );
  DFFHQXL H7_reg_14_ ( .D(n2433), .CK(clk), .Q(H7[14]) );
  DFFHQXL H2_reg_13_ ( .D(n2562), .CK(clk), .Q(H2[13]) );
  DFFHQXL H2_reg_14_ ( .D(n2561), .CK(clk), .Q(H2[14]) );
  DFFHQXL H3_reg_13_ ( .D(n2593), .CK(clk), .Q(H3[13]) );
  DFFHQXL H3_reg_14_ ( .D(n2592), .CK(clk), .Q(H3[14]) );
  DFFHQXL H2_reg_12_ ( .D(n2563), .CK(clk), .Q(H2[12]) );
  DFFHQXL H3_reg_12_ ( .D(n2594), .CK(clk), .Q(H3[12]) );
  DFFHQXL H1_reg_12_ ( .D(n2851), .CK(clk), .Q(H1[12]) );
  DFFHQXL H5_reg_14_ ( .D(n2656), .CK(clk), .Q(H5[14]) );
  DFFHQXL G_reg_25_ ( .D(n2486), .CK(clk), .Q(SHA256_result[57]) );
  DFFHQXL G_reg_27_ ( .D(n2484), .CK(clk), .Q(SHA256_result[59]) );
  DFFHQXL C_reg_16_ ( .D(n2782), .CK(clk), .Q(SHA256_result[176]) );
  DFFHQXL C_reg_17_ ( .D(n2781), .CK(clk), .Q(SHA256_result[177]) );
  DFFHQXL C_reg_18_ ( .D(n2780), .CK(clk), .Q(SHA256_result[178]) );
  DFFHQXL H_reg_20_ ( .D(n2459), .CK(clk), .Q(SHA256_result[20]) );
  DFFHQXL H_reg_22_ ( .D(n2457), .CK(clk), .Q(SHA256_result[22]) );
  DFFHQXL H_reg_23_ ( .D(n2456), .CK(clk), .Q(SHA256_result[23]) );
  DFFHQXL D_reg_1_ ( .D(n2765), .CK(clk), .Q(SHA256_result[129]) );
  DFFHQXL C_reg_19_ ( .D(n2779), .CK(clk), .Q(SHA256_result[179]) );
  DFFXL F_reg_26_ ( .D(n2676), .CK(clk), .Q(SHA256_result[90]), .QN(n1142) );
  DFFHQXL G_reg_26_ ( .D(n2485), .CK(clk), .Q(SHA256_result[58]) );
  DFFXL F_reg_24_ ( .D(n2678), .CK(clk), .Q(SHA256_result[88]), .QN(n1144) );
  DFFHQXL B_reg_19_ ( .D(n2812), .CK(clk), .Q(SHA256_result[211]) );
  DFFHQXL H0_reg_5_ ( .D(n2922), .CK(clk), .Q(H0[5]) );
  DFFHQXL H0_reg_1_ ( .D(n2926), .CK(clk), .Q(H0[1]) );
  DFFHQX1 H_reg_12_ ( .D(n2467), .CK(clk), .Q(SHA256_result[12]) );
  DFFHQX1 H_reg_13_ ( .D(n2466), .CK(clk), .Q(SHA256_result[13]) );
  DFFHQX1 H_reg_5_ ( .D(n2474), .CK(clk), .Q(SHA256_result[5]) );
  DFFHQX1 G_reg_18_ ( .D(n2493), .CK(clk), .Q(SHA256_result[50]) );
  DFFHQX1 G_reg_19_ ( .D(n2492), .CK(clk), .Q(SHA256_result[51]) );
  DFFHQX1 G_reg_6_ ( .D(n2505), .CK(clk), .Q(SHA256_result[38]) );
  DFFHQX1 C_reg_13_ ( .D(n2785), .CK(clk), .Q(SHA256_result[173]) );
  DFFX1 F_reg_27_ ( .D(n2675), .CK(clk), .Q(SHA256_result[91]), .QN(n1141) );
  DFFHQX1 H6_reg_27_ ( .D(n2515), .CK(clk), .Q(H6[27]) );
  DFFHQXL H5_reg_12_ ( .D(n2658), .CK(clk), .Q(H5[12]) );
  DFFHQXL H6_reg_11_ ( .D(n2531), .CK(clk), .Q(H6[11]) );
  DFFHQXL H7_reg_11_ ( .D(n2436), .CK(clk), .Q(H7[11]) );
  DFFHQXL H5_reg_11_ ( .D(n2659), .CK(clk), .Q(H5[11]) );
  DFFHQXL C_reg_15_ ( .D(n2783), .CK(clk), .Q(SHA256_result[175]) );
  DFFHQXL F_reg_22_ ( .D(n2680), .CK(clk), .Q(SHA256_result[86]) );
  DFFHQXL G_reg_21_ ( .D(n2490), .CK(clk), .Q(SHA256_result[53]) );
  DFFHQXL F_reg_21_ ( .D(n2681), .CK(clk), .Q(SHA256_result[85]) );
  DFFHQXL G_reg_22_ ( .D(n2489), .CK(clk), .Q(SHA256_result[54]) );
  DFFHQXL B_reg_15_ ( .D(n2816), .CK(clk), .Q(SHA256_result[207]) );
  DFFHQX1 C_reg_14_ ( .D(n2784), .CK(clk), .Q(SHA256_result[174]) );
  DFFHQX1 H7_reg_24_ ( .D(n2423), .CK(clk), .Q(H7[24]) );
  DFFHQX1 G_reg_24_ ( .D(n2487), .CK(clk), .Q(SHA256_result[56]) );
  DFFHQX1 H2_reg_16_ ( .D(n2559), .CK(clk), .Q(H2[16]) );
  DFFHQXL H6_reg_10_ ( .D(n2532), .CK(clk), .Q(H6[10]) );
  DFFHQX4 H6_reg_0_ ( .D(n2542), .CK(clk), .Q(H6[0]) );
  DFFHQXL H3_reg_10_ ( .D(n2596), .CK(clk), .Q(H3[10]) );
  DFFHQX1 B_reg_17_ ( .D(n2814), .CK(clk), .Q(SHA256_result[209]) );
  DFFHQX1 B_reg_16_ ( .D(n2815), .CK(clk), .Q(SHA256_result[208]) );
  DFFX4 F_reg_0_ ( .D(n2702), .CK(clk), .Q(SHA256_result[64]), .QN(n1168) );
  DFFHQX4 H2_reg_1_ ( .D(n2574), .CK(clk), .Q(H2[1]) );
  DFFTRX1 round_reg_5_ ( .D(N126), .RN(n129), .CK(clk), .Q(round[5]), .QN(
        n1370) );
  DFFHQX1 H3_reg_7_ ( .D(n2599), .CK(clk), .Q(H3[7]) );
  DFFHQX1 H5_reg_8_ ( .D(n2662), .CK(clk), .Q(H5[8]) );
  DFFHQX1 H6_reg_9_ ( .D(n2533), .CK(clk), .Q(H6[9]) );
  DFFHQX1 H7_reg_9_ ( .D(n2438), .CK(clk), .Q(H7[9]) );
  DFFHQX1 H1_reg_9_ ( .D(n2854), .CK(clk), .Q(H1[9]) );
  DFFHQX1 H7_reg_10_ ( .D(n2437), .CK(clk), .Q(H7[10]) );
  DFFHQX1 E_reg_20_ ( .D(n2714), .CK(clk), .Q(SHA256_result[116]) );
  DFFHQX1 E_reg_21_ ( .D(n2713), .CK(clk), .Q(SHA256_result[117]) );
  DFFHQX1 H7_reg_6_ ( .D(n2441), .CK(clk), .Q(H7[6]) );
  DFFHQX1 H1_reg_7_ ( .D(n2856), .CK(clk), .Q(H1[7]) );
  DFFHQX1 H2_reg_8_ ( .D(n2567), .CK(clk), .Q(H2[8]) );
  DFFHQX1 H5_reg_7_ ( .D(n2663), .CK(clk), .Q(H5[7]) );
  DFFHQX1 H6_reg_7_ ( .D(n2535), .CK(clk), .Q(H6[7]) );
  DFFHQX1 H6_reg_8_ ( .D(n2534), .CK(clk), .Q(H6[8]) );
  DFFHQX1 H7_reg_8_ ( .D(n2439), .CK(clk), .Q(H7[8]) );
  DFFHQX1 G_reg_11_ ( .D(n2500), .CK(clk), .Q(SHA256_result[43]) );
  DFFHQX1 H_reg_2_ ( .D(n2477), .CK(clk), .Q(SHA256_result[2]) );
  DFFHQX1 H6_reg_6_ ( .D(n2536), .CK(clk), .Q(H6[6]) );
  DFFHQX1 H5_reg_4_ ( .D(n2666), .CK(clk), .Q(H5[4]) );
  DFFHQX1 H6_reg_5_ ( .D(n2537), .CK(clk), .Q(H6[5]) );
  DFFHQX1 H_reg_1_ ( .D(n2478), .CK(clk), .Q(SHA256_result[1]) );
  DFFHQX1 C_reg_3_ ( .D(n2795), .CK(clk), .Q(SHA256_result[163]) );
  DFFHQX1 E_reg_22_ ( .D(n2712), .CK(clk), .Q(SHA256_result[118]) );
  DFFHQX1 H_reg_0_ ( .D(n2479), .CK(clk), .Q(SHA256_result[0]) );
  DFFHQX4 H7_reg_0_ ( .D(n2447), .CK(clk), .Q(H7[0]) );
  DFFHQX4 H7_reg_1_ ( .D(n2446), .CK(clk), .Q(H7[1]) );
  DFFX4 A_reg_1_ ( .D(n2894), .CK(clk), .Q(n91), .QN(n92) );
  DFFHQX4 E_reg_30_ ( .D(n2704), .CK(clk), .Q(SHA256_result[126]) );
  DFFX4 B_reg_0_ ( .D(n2831), .CK(clk), .Q(n89), .QN(n88) );
  DFFHQX4 E_reg_5_ ( .D(n2729), .CK(clk), .Q(SHA256_result[101]) );
  DFFX4 G_reg_0_ ( .D(n2543), .CK(clk), .Q(n82), .QN(n81) );
  DFFX4 B_reg_1_ ( .D(n2830), .CK(clk), .Q(n79), .QN(n78) );
  DFFHQXL F_reg_31_ ( .D(n2671), .CK(clk), .Q(SHA256_result[95]) );
  DFFHQX4 H1_reg_0_ ( .D(n2863), .CK(clk), .Q(H1[0]) );
  DFFHQX4 F_reg_4_ ( .D(n2698), .CK(clk), .Q(SHA256_result[68]) );
  DFFHQX2 G_reg_13_ ( .D(n2498), .CK(clk), .Q(SHA256_result[45]) );
  DFFX2 F_reg_15_ ( .D(n2687), .CK(clk), .Q(SHA256_result[79]), .QN(n1153) );
  DFFHQXL E_reg_29_ ( .D(n2705), .CK(clk), .Q(SHA256_result[125]) );
  DFFX2 F_reg_14_ ( .D(n2688), .CK(clk), .Q(SHA256_result[78]), .QN(n1154) );
  DFFX2 F_reg_8_ ( .D(n2694), .CK(clk), .Q(SHA256_result[72]), .QN(n1160) );
  DFFHQX2 G_reg_9_ ( .D(n2502), .CK(clk), .Q(SHA256_result[41]) );
  DFFHQX4 G_reg_8_ ( .D(n2503), .CK(clk), .Q(SHA256_result[40]) );
  DFFHQX4 E_reg_31_ ( .D(n2703), .CK(clk), .Q(SHA256_result[127]) );
  DFFHQX2 F_reg_9_ ( .D(n2693), .CK(clk), .Q(SHA256_result[73]) );
  DFFHQXL A_reg_23_ ( .D(n2872), .CK(clk), .Q(SHA256_result[247]) );
  DFFTRXL round_reg_4_ ( .D(N125), .RN(n129), .CK(clk), .Q(round[4]), .QN(n32)
         );
  DFFHQX4 H2_reg_0_ ( .D(n2799), .CK(clk), .Q(n99) );
  DFFXL read_counter_reg_1_ ( .D(N3080), .CK(clk), .Q(read_counter[1]), .QN(
        n972) );
  DFFHQX2 B_reg_2_ ( .D(n2829), .CK(clk), .Q(SHA256_result[194]) );
  DFFHQX1 B_reg_3_ ( .D(n2828), .CK(clk), .Q(SHA256_result[195]) );
  DFFTRX1 round_reg_1_ ( .D(N122), .RN(n129), .CK(clk), .Q(round[1]), .QN(
        n1393) );
  DFFTRX2 round_reg_2_ ( .D(N123), .RN(n129), .CK(clk), .Q(round[2]), .QN(
        n1388) );
  DFFTRX2 round_reg_3_ ( .D(N124), .RN(n129), .CK(clk), .Q(round[3]), .QN(
        n1383) );
  DFFHQX2 E_reg_26_ ( .D(n2708), .CK(clk), .Q(SHA256_result[122]) );
  DFFHQX2 E_reg_27_ ( .D(n2707), .CK(clk), .Q(SHA256_result[123]) );
  DFFHQX2 E_reg_28_ ( .D(n2706), .CK(clk), .Q(SHA256_result[124]) );
  DFFHQX2 F_reg_2_ ( .D(n2700), .CK(clk), .Q(SHA256_result[66]) );
  DFFHQX2 G_reg_2_ ( .D(n2509), .CK(clk), .Q(SHA256_result[34]) );
  DFFHQX2 G_reg_3_ ( .D(n2508), .CK(clk), .Q(SHA256_result[35]) );
  DFFHQX2 G_reg_7_ ( .D(n2504), .CK(clk), .Q(SHA256_result[39]) );
  DFFHQX2 Kt_reg_15_ ( .D(N2961), .CK(clk), .Q(Kt[15]) );
  DFFHQX2 Kt_reg_14_ ( .D(N2960), .CK(clk), .Q(Kt[14]) );
  DFFHQX2 Kt_reg_12_ ( .D(N2958), .CK(clk), .Q(Kt[12]) );
  DFFHQX2 Kt_reg_11_ ( .D(N2957), .CK(clk), .Q(Kt[11]) );
  DFFHQX2 Kt_reg_10_ ( .D(N2956), .CK(clk), .Q(Kt[10]) );
  DFFHQX2 Kt_reg_9_ ( .D(N2955), .CK(clk), .Q(Kt[9]) );
  DFFHQX2 Kt_reg_5_ ( .D(N2951), .CK(clk), .Q(Kt[5]) );
  DFFHQXL A_reg_31_ ( .D(n2864), .CK(clk), .Q(SHA256_result[255]) );
  DFFHQX1 H6_reg_25_ ( .D(n2517), .CK(clk), .Q(H6[25]) );
  DFFX1 F_reg_25_ ( .D(n2677), .CK(clk), .Q(SHA256_result[89]), .QN(n1143) );
  DFFHQX1 H1_reg_17_ ( .D(n2846), .CK(clk), .Q(H1[17]) );
  DFFHQX1 H1_reg_28_ ( .D(n2835), .CK(clk), .Q(H1[28]) );
  DFFHQX2 A_reg_28_ ( .D(n2867), .CK(clk), .Q(SHA256_result[252]) );
  DFFHQX1 H6_reg_18_ ( .D(n2524), .CK(clk), .Q(H6[18]) );
  DFFHQX1 F_reg_18_ ( .D(n2684), .CK(clk), .Q(SHA256_result[82]) );
  DFFHQX1 H7_reg_5_ ( .D(n2442), .CK(clk), .Q(H7[5]) );
  DFFX2 F_reg_5_ ( .D(n2697), .CK(clk), .Q(SHA256_result[69]), .QN(n1163) );
  DFFHQX2 C_reg_2_ ( .D(n2796), .CK(clk), .Q(SHA256_result[162]) );
  DFFHQX1 H7_reg_20_ ( .D(n2427), .CK(clk), .Q(H7[20]) );
  DFFHQX1 G_reg_20_ ( .D(n2491), .CK(clk), .Q(SHA256_result[52]) );
  DFFHQX1 H1_reg_10_ ( .D(n2853), .CK(clk), .Q(H1[10]) );
  DFFHQX1 H6_reg_4_ ( .D(n2538), .CK(clk), .Q(H6[4]) );
  DFFHQX2 H1_reg_1_ ( .D(n2862), .CK(clk), .Q(H1[1]) );
  DFFHQX1 H1_reg_2_ ( .D(n2861), .CK(clk), .Q(H1[2]) );
  DFFHQX2 E_reg_16_ ( .D(n2718), .CK(clk), .Q(SHA256_result[112]) );
  DFFHQX2 E_reg_17_ ( .D(n2717), .CK(clk), .Q(SHA256_result[113]) );
  DFFHQX1 B_reg_4_ ( .D(n2827), .CK(clk), .Q(SHA256_result[196]) );
  DFFHQX2 G_reg_14_ ( .D(n2497), .CK(clk), .Q(SHA256_result[46]) );
  DFFHQX2 G_reg_12_ ( .D(n2499), .CK(clk), .Q(SHA256_result[44]) );
  DFFHQX2 G_reg_15_ ( .D(n2496), .CK(clk), .Q(SHA256_result[47]) );
  DFFHQX2 G_reg_4_ ( .D(n2507), .CK(clk), .Q(SHA256_result[36]) );
  DFFHQX1 H1_reg_23_ ( .D(n2840), .CK(clk), .Q(H1[23]) );
  DFFHQX2 B_reg_7_ ( .D(n2824), .CK(clk), .Q(SHA256_result[199]) );
  DFFHQX1 E_reg_19_ ( .D(n2715), .CK(clk), .Q(SHA256_result[115]) );
  DFFX2 F_reg_12_ ( .D(n2690), .CK(clk), .Q(SHA256_result[76]), .QN(n1156) );
  DFFHQX2 F_reg_13_ ( .D(n2689), .CK(clk), .Q(SHA256_result[77]) );
  EDFFTRX1 round_reg_6_ ( .RN(N127), .D(n129), .E(1'b1), .CK(clk), .Q(round[6]), .QN(n392) );
  DFFHQX2 H3_reg_1_ ( .D(n2605), .CK(clk), .Q(n71) );
  DFFHQX1 A_reg_2_ ( .D(n2893), .CK(clk), .Q(SHA256_result[226]) );
  DFFHQX4 H5_reg_1_ ( .D(n2669), .CK(clk), .Q(H5[1]) );
  DFFHQX4 H5_reg_0_ ( .D(n2670), .CK(clk), .Q(H5[0]) );
  DFFHQX4 H6_reg_1_ ( .D(n2541), .CK(clk), .Q(n96) );
  DFFHQX4 H3_reg_0_ ( .D(n2606), .CK(clk), .Q(H3[0]) );
  DFFHQX2 F_reg_10_ ( .D(n2692), .CK(clk), .Q(SHA256_result[74]) );
  DFFHQX4 E_reg_7_ ( .D(n2727), .CK(clk), .Q(SHA256_result[103]) );
  DFFHQX4 A_reg_22_ ( .D(n2873), .CK(clk), .Q(SHA256_result[246]) );
  DFFHQX2 G_reg_10_ ( .D(n2501), .CK(clk), .Q(SHA256_result[42]) );
  DFFHQX4 E_reg_25_ ( .D(n2709), .CK(clk), .Q(SHA256_result[121]) );
  DFFHQX1 C_reg_9_ ( .D(n2789), .CK(clk), .Q(SHA256_result[169]) );
  DFFX2 F_reg_11_ ( .D(n2691), .CK(clk), .Q(SHA256_result[75]), .QN(n1157) );
  DFFHQX4 E_reg_3_ ( .D(n2731), .CK(clk), .Q(SHA256_result[99]) );
  DFFHQX2 F_reg_6_ ( .D(n2696), .CK(clk), .Q(SHA256_result[70]) );
  DFFX2 F_reg_3_ ( .D(n2699), .CK(clk), .Q(SHA256_result[67]), .QN(n1165) );
  DFFHQX4 Kt_reg_7_ ( .D(N2953), .CK(clk), .Q(Kt[7]) );
  CLKINVX3 U3 ( .A(n211), .Y(n210) );
  NAND2X2 U4 ( .A(N814), .B(n202), .Y(n653) );
  OAI2BB1X4 U5 ( .A0N(n199), .A1N(N952), .B0(n454), .Y(n2705) );
  NOR2BX4 U15 ( .AN(first_block), .B(n1490), .Y(n128) );
  INVX8 U16 ( .A(n128), .Y(n677) );
  CLKINVX8 U17 ( .A(n91), .Y(n64) );
  CLKBUFX8 U18 ( .A(SHA256_result[242]), .Y(n141) );
  NAND2X2 U19 ( .A(N951), .B(n196), .Y(n456) );
  NAND2X4 U20 ( .A(N822), .B(n204), .Y(n626) );
  NAND2X4 U21 ( .A(n120), .B(n121), .Y(n10) );
  NAND2X4 U22 ( .A(n11), .B(n1755), .Y(n2800) );
  CLKINVX4 U23 ( .A(n10), .Y(n11) );
  NOR2XL U24 ( .A(round[6]), .B(n1849), .Y(n12) );
  NOR2XL U25 ( .A(n13), .B(n224), .Y(n126) );
  INVX1 U26 ( .A(n12), .Y(n13) );
  INVX12 U27 ( .A(n126), .Y(n23) );
  NAND2X1 U28 ( .A(n619), .B(n620), .Y(n14) );
  NAND2X4 U29 ( .A(n15), .B(n618), .Y(n2865) );
  CLKINVX3 U30 ( .A(n14), .Y(n15) );
  OAI2BB1X2 U31 ( .A0N(N950), .A1N(n717), .B0(n462), .Y(n2707) );
  XOR3X4 U32 ( .A(n140), .B(n151), .C(SHA256_result[252]), .Y(f3_A_32[6]) );
  OAI2BB1X2 U33 ( .A0N(SHA256_result[200]), .A1N(n151), .B0(n607), .Y(
        f2_ABC_32[8]) );
  BUFX8 U34 ( .A(SHA256_result[232]), .Y(n151) );
  NAND2X4 U35 ( .A(n117), .B(n1493), .Y(n2480) );
  NAND2X4 U36 ( .A(N825), .B(n197), .Y(n618) );
  OAI2BB1X4 U37 ( .A0N(N823), .A1N(n205), .B0(n625), .Y(n2867) );
  OAI211X4 U38 ( .A0(n283), .A1(n445), .B0(n413), .C0(n412), .Y(n2509) );
  NAND2X1 U39 ( .A(n445), .B(SHA256_result[98]), .Y(n74) );
  INVX2 U40 ( .A(SHA256_result[66]), .Y(n445) );
  OAI2BB1X4 U41 ( .A0N(n205), .A1N(N826), .B0(n617), .Y(n2864) );
  MXI2X4 U42 ( .A(n444), .B(n1165), .S0(SHA256_result[99]), .Y(f1_EFG_32[3])
         );
  MXI2X4 U43 ( .A(n918), .B(n1157), .S0(SHA256_result[107]), .Y(f1_EFG_32[11])
         );
  OAI221X4 U44 ( .A0(n315), .A1(n1157), .B0(n194), .B1(n918), .C0(n1513), .Y(
        n2500) );
  OAI21X1 U45 ( .A0(SHA256_result[201]), .A1(n150), .B0(SHA256_result[169]), 
        .Y(n606) );
  CLKBUFX8 U46 ( .A(SHA256_result[243]), .Y(n140) );
  OAI2BB1X4 U47 ( .A0N(N948), .A1N(n202), .B0(n470), .Y(n2709) );
  MXI2X4 U48 ( .A(n921), .B(n1154), .S0(SHA256_result[110]), .Y(f1_EFG_32[14])
         );
  INVX8 U49 ( .A(SHA256_result[46]), .Y(n921) );
  MX2X4 U50 ( .A(SHA256_result[41]), .B(SHA256_result[73]), .S0(
        SHA256_result[105]), .Y(f1_EFG_32[9]) );
  XOR3X2 U51 ( .A(SHA256_result[110]), .B(SHA256_result[105]), .C(
        SHA256_result[124]), .Y(f4_E_32[3]) );
  NOR3XL U52 ( .A(n1849), .B(round[6]), .C(n224), .Y(n16) );
  BUFX3 U53 ( .A(n340), .Y(n17) );
  BUFX4 U54 ( .A(n27), .Y(n18) );
  BUFX12 U55 ( .A(n26), .Y(n19) );
  BUFX3 U56 ( .A(n28), .Y(n20) );
  BUFX3 U57 ( .A(n30), .Y(n21) );
  BUFX3 U58 ( .A(n29), .Y(n22) );
  INVX4 U59 ( .A(n16), .Y(n24) );
  CLKINVX3 U60 ( .A(n340), .Y(n341) );
  INVXL U61 ( .A(n126), .Y(n340) );
  INVX1 U62 ( .A(n341), .Y(n27) );
  INVXL U63 ( .A(n126), .Y(n28) );
  BUFX3 U64 ( .A(n27), .Y(n30) );
  MXI2X4 U65 ( .A(n919), .B(n1156), .S0(SHA256_result[108]), .Y(f1_EFG_32[12])
         );
  INVX8 U66 ( .A(SHA256_result[44]), .Y(n919) );
  MXI2X2 U67 ( .A(n81), .B(n1168), .S0(SHA256_result[96]), .Y(f1_EFG_32[0]) );
  OAI2BB1X4 U68 ( .A0N(N817), .A1N(n200), .B0(n648), .Y(n2873) );
  XOR3X4 U69 ( .A(SHA256_result[108]), .B(SHA256_result[103]), .C(
        SHA256_result[122]), .Y(f4_E_32[1]) );
  MXI2X4 U70 ( .A(n914), .B(n1161), .S0(SHA256_result[103]), .Y(f1_EFG_32[7])
         );
  NAND2X4 U71 ( .A(n105), .B(n1724), .Y(n2768) );
  NOR2X4 U72 ( .A(n106), .B(n107), .Y(n1724) );
  MX2X4 U73 ( .A(SHA256_result[42]), .B(SHA256_result[74]), .S0(
        SHA256_result[106]), .Y(f1_EFG_32[10]) );
  NAND3X4 U74 ( .A(n123), .B(n124), .C(n1691), .Y(n2735) );
  AND2X4 U75 ( .A(n125), .B(n677), .Y(n1691) );
  NAND2X4 U76 ( .A(N922), .B(n197), .Y(n125) );
  OAI211XL U77 ( .A0(n23), .A1(n447), .B0(n62), .C0(n1540), .Y(n2541) );
  BUFX8 U78 ( .A(SHA256_result[255]), .Y(n25) );
  OAI2BB2X1 U79 ( .B0(n342), .B1(n1168), .A0N(H5[0]), .A1N(n226), .Y(n2670) );
  OAI2BB1X4 U80 ( .A0N(n1489), .A1N(SHA256_result[31]), .B0(n1454), .Y(n2448)
         );
  NAND3X4 U81 ( .A(n97), .B(n98), .C(n1458), .Y(n2449) );
  NAND2X4 U82 ( .A(n104), .B(n1723), .Y(n2767) );
  OAI2BB2XL U83 ( .B0(n342), .B1(n1167), .A0N(H5[1]), .A1N(n226), .Y(n2669) );
  OAI21X1 U84 ( .A0(n157), .A1(SHA256_result[194]), .B0(SHA256_result[162]), 
        .Y(n613) );
  OAI2BB1X2 U85 ( .A0N(SHA256_result[194]), .A1N(n157), .B0(n613), .Y(
        f2_ABC_32[2]) );
  BUFX12 U86 ( .A(SHA256_result[226]), .Y(n157) );
  NAND2X2 U87 ( .A(n85), .B(n86), .Y(n87) );
  MXI2X2 U88 ( .A(n915), .B(n1160), .S0(SHA256_result[104]), .Y(f1_EFG_32[8])
         );
  NAND2X2 U89 ( .A(n1859), .B(n392), .Y(n390) );
  CLKINVX3 U90 ( .A(n266), .Y(n338) );
  INVX1 U91 ( .A(n188), .Y(n186) );
  INVX1 U92 ( .A(n339), .Y(n277) );
  NAND2X2 U93 ( .A(N1016), .B(n206), .Y(n94) );
  BUFX3 U94 ( .A(SHA256_result[125]), .Y(n51) );
  CLKBUFX8 U95 ( .A(SHA256_result[247]), .Y(n137) );
  INVX1 U96 ( .A(n278), .Y(n274) );
  MX2X2 U97 ( .A(SHA256_result[45]), .B(SHA256_result[77]), .S0(
        SHA256_result[109]), .Y(f1_EFG_32[13]) );
  MX2X1 U98 ( .A(SHA256_result[51]), .B(SHA256_result[83]), .S0(
        SHA256_result[115]), .Y(f1_EFG_32[19]) );
  MXI2X1 U99 ( .A(n923), .B(n1152), .S0(SHA256_result[112]), .Y(f1_EFG_32[16])
         );
  XOR3X2 U100 ( .A(SHA256_result[112]), .B(SHA256_result[107]), .C(
        SHA256_result[126]), .Y(f4_E_32[5]) );
  OAI2BB1X1 U101 ( .A0N(SHA256_result[196]), .A1N(n155), .B0(n611), .Y(
        f2_ABC_32[4]) );
  OAI2BB1X1 U102 ( .A0N(SHA256_result[195]), .A1N(n156), .B0(n612), .Y(
        f2_ABC_32[3]) );
  XOR3X2 U103 ( .A(SHA256_result[107]), .B(SHA256_result[102]), .C(
        SHA256_result[121]), .Y(f4_E_32[0]) );
  CLKINVX3 U104 ( .A(n46), .Y(n47) );
  CLKINVX3 U105 ( .A(n1491), .Y(n389) );
  BUFX3 U106 ( .A(next_A[20]), .Y(n43) );
  INVX1 U107 ( .A(n1437), .Y(n52) );
  INVX1 U108 ( .A(n189), .Y(n185) );
  BUFX3 U109 ( .A(next_E[30]), .Y(n44) );
  INVX1 U110 ( .A(SHA256_result[37]), .Y(n441) );
  INVX1 U111 ( .A(n53), .Y(n61) );
  INVX8 U112 ( .A(n228), .Y(n224) );
  BUFX3 U113 ( .A(SHA256_result[224]), .Y(n158) );
  BUFX3 U114 ( .A(SHA256_result[233]), .Y(n150) );
  BUFX3 U115 ( .A(SHA256_result[234]), .Y(n149) );
  BUFX3 U116 ( .A(SHA256_result[235]), .Y(n148) );
  CLKBUFX8 U117 ( .A(SHA256_result[241]), .Y(n142) );
  BUFX3 U118 ( .A(SHA256_result[244]), .Y(n139) );
  BUFX3 U119 ( .A(SHA256_result[245]), .Y(n138) );
  BUFX3 U120 ( .A(SHA256_result[248]), .Y(n136) );
  BUFX3 U121 ( .A(SHA256_result[250]), .Y(n134) );
  BUFX3 U122 ( .A(SHA256_result[38]), .Y(n50) );
  INVX2 U123 ( .A(SHA256_result[36]), .Y(n443) );
  INVX1 U124 ( .A(SHA256_result[35]), .Y(n444) );
  INVX1 U125 ( .A(SHA256_result[34]), .Y(n446) );
  INVX8 U126 ( .A(n37), .Y(n342) );
  BUFX3 U127 ( .A(SHA256_result[227]), .Y(n156) );
  BUFX4 U128 ( .A(SHA256_result[229]), .Y(n154) );
  INVX1 U129 ( .A(SHA256_result[49]), .Y(n924) );
  INVX1 U130 ( .A(SHA256_result[48]), .Y(n923) );
  INVX2 U131 ( .A(SHA256_result[47]), .Y(n922) );
  BUFX3 U132 ( .A(SHA256_result[253]), .Y(n132) );
  BUFX3 U133 ( .A(SHA256_result[240]), .Y(n143) );
  BUFX3 U134 ( .A(SHA256_result[231]), .Y(n152) );
  BUFX3 U135 ( .A(SHA256_result[230]), .Y(n153) );
  BUFX3 U136 ( .A(SHA256_result[238]), .Y(n145) );
  BUFX3 U137 ( .A(SHA256_result[236]), .Y(n147) );
  NOR2X1 U138 ( .A(n792), .B(n161), .Y(n1878) );
  NOR2X1 U139 ( .A(n797), .B(n160), .Y(n2148) );
  BUFX3 U140 ( .A(round[5]), .Y(n160) );
  INVX1 U141 ( .A(SHA256_result[39]), .Y(n914) );
  OAI2BB1X2 U142 ( .A0N(N818), .A1N(n203), .B0(n644), .Y(n2872) );
  OAI221XL U143 ( .A0(n303), .A1(n1160), .B0(n191), .B1(n915), .C0(n1516), .Y(
        n2503) );
  OAI211X1 U144 ( .A0(n484), .A1(n320), .B0(n483), .C0(n482), .Y(n2715) );
  NAND2X1 U145 ( .A(N942), .B(n195), .Y(n482) );
  OAI211X1 U146 ( .A0(n282), .A1(n442), .B0(n408), .C0(n407), .Y(n2507) );
  OAI21XL U147 ( .A0(n163), .A1(n1160), .B0(n1633), .Y(n2694) );
  OAI21XL U148 ( .A0(n164), .A1(n1153), .B0(n1626), .Y(n2687) );
  OAI21XL U149 ( .A0(n88), .A1(n176), .B0(n677), .Y(n583) );
  OAI21XL U150 ( .A0(n342), .A1(n442), .B0(n431), .Y(n2666) );
  NAND2X1 U151 ( .A(n93), .B(n1495), .Y(n2482) );
  AND2X2 U152 ( .A(n94), .B(n95), .Y(n1495) );
  NAND2X1 U153 ( .A(SHA256_result[93]), .B(n274), .Y(n95) );
  OR2X2 U154 ( .A(n311), .B(n937), .Y(n97) );
  OR2X2 U155 ( .A(n1457), .B(n970), .Y(n98) );
  NAND2X1 U156 ( .A(N810), .B(n203), .Y(n663) );
  AOI221X1 U157 ( .A0(n254), .A1(SHA256_result[13]), .B0(n248), .B1(
        SHA256_result[45]), .C0(n2061), .Y(n2060) );
  AOI221X1 U158 ( .A0(n254), .A1(SHA256_result[15]), .B0(n248), .B1(
        SHA256_result[47]), .C0(n2053), .Y(n2052) );
  OAI2BB1X1 U159 ( .A0N(N946), .A1N(n199), .B0(n475), .Y(n2711) );
  NAND2X1 U160 ( .A(N941), .B(n204), .Y(n485) );
  NAND2X2 U161 ( .A(n38), .B(n626), .Y(n2868) );
  AOI21X1 U162 ( .A0(n182), .A1(n133), .B0(n256), .Y(n628) );
  NAND3X1 U163 ( .A(n636), .B(n635), .C(n634), .Y(n2870) );
  NAND2X1 U164 ( .A(N820), .B(n199), .Y(n634) );
  NAND3X1 U165 ( .A(n458), .B(n457), .C(n456), .Y(n2706) );
  OAI2BB1X1 U166 ( .A0N(N949), .A1N(n200), .B0(n466), .Y(n2708) );
  OAI2BB1X1 U167 ( .A0N(N938), .A1N(n197), .B0(n493), .Y(n2719) );
  NAND2X2 U168 ( .A(n441), .B(n84), .Y(n85) );
  CLKINVX3 U169 ( .A(SHA256_result[101]), .Y(n84) );
  NAND2X2 U170 ( .A(n446), .B(n72), .Y(n73) );
  INVX2 U171 ( .A(SHA256_result[98]), .Y(n72) );
  NAND2X2 U172 ( .A(n443), .B(n531), .Y(n76) );
  INVX4 U173 ( .A(SHA256_result[100]), .Y(n531) );
  INVXL U174 ( .A(n341), .Y(n26) );
  BUFX3 U175 ( .A(n26), .Y(n29) );
  CLKINVX3 U176 ( .A(n209), .Y(n203) );
  CLKINVX3 U177 ( .A(n171), .Y(n162) );
  CLKINVX3 U178 ( .A(n207), .Y(n197) );
  CLKINVX3 U179 ( .A(n208), .Y(n202) );
  CLKINVX3 U180 ( .A(n53), .Y(n58) );
  CLKINVX3 U181 ( .A(n209), .Y(n199) );
  CLKINVX2 U182 ( .A(n53), .Y(n62) );
  CLKINVX3 U183 ( .A(n53), .Y(n60) );
  CLKINVX3 U184 ( .A(n207), .Y(n204) );
  OAI21XL U185 ( .A0(first_block), .A1(n393), .B0(n1491), .Y(n703) );
  INVX1 U186 ( .A(SHA256_result[96]), .Y(n70) );
  CLKINVX3 U187 ( .A(n209), .Y(n195) );
  INVX1 U188 ( .A(n208), .Y(n198) );
  INVX1 U189 ( .A(n677), .Y(n257) );
  CLKINVX3 U190 ( .A(n52), .Y(n54) );
  INVX1 U191 ( .A(n53), .Y(n59) );
  INVX1 U192 ( .A(n113), .Y(n769) );
  INVX1 U193 ( .A(n224), .Y(n211) );
  INVX1 U194 ( .A(n209), .Y(n196) );
  INVXL U195 ( .A(n1985), .Y(n245) );
  CLKINVX3 U196 ( .A(SHA256_result[97]), .Y(n68) );
  BUFX4 U197 ( .A(n69), .Y(n67) );
  NOR2X1 U198 ( .A(n1370), .B(n346), .Y(n31) );
  INVX1 U199 ( .A(n1456), .Y(n267) );
  CLKINVX3 U200 ( .A(n208), .Y(n200) );
  INVX1 U201 ( .A(n188), .Y(n187) );
  INVX1 U202 ( .A(round[4]), .Y(n346) );
  OR3XL U203 ( .A(n971), .B(read_counter[1]), .C(n973), .Y(n33) );
  OR3XL U204 ( .A(read_counter[1]), .B(read_counter[2]), .C(read_counter[0]), 
        .Y(n34) );
  OR3XL U205 ( .A(n972), .B(read_counter[0]), .C(n973), .Y(n35) );
  OR3XL U206 ( .A(n972), .B(n971), .C(n973), .Y(n36) );
  NOR2X1 U207 ( .A(first_block), .B(n23), .Y(n37) );
  CLKINVX3 U208 ( .A(n52), .Y(n57) );
  CLKINVX3 U209 ( .A(n52), .Y(n55) );
  CLKINVX3 U210 ( .A(n52), .Y(n56) );
  AND2X2 U211 ( .A(n627), .B(n628), .Y(n38) );
  AND2X2 U212 ( .A(n73), .B(n74), .Y(n39) );
  AND2X2 U213 ( .A(n76), .B(n77), .Y(n40) );
  INVX1 U214 ( .A(n81), .Y(n83) );
  INVX1 U215 ( .A(n208), .Y(n201) );
  NOR2X1 U216 ( .A(n1370), .B(n159), .Y(n41) );
  INVX1 U217 ( .A(n78), .Y(n80) );
  INVX1 U218 ( .A(n88), .Y(n90) );
  AOI21XL U220 ( .A0(N886), .A1(n199), .B0(n261), .Y(n1727) );
  XOR3X2 U221 ( .A(n157), .B(n146), .C(SHA256_result[246]), .Y(f3_A_32[0]) );
  AOI21XL U222 ( .A0(N1027), .A1(n205), .B0(n258), .Y(n1481) );
  AOI21XL U223 ( .A0(N979), .A1(n200), .B0(n259), .Y(n1617) );
  AOI21XL U224 ( .A0(N917), .A1(n199), .B0(n259), .Y(n1696) );
  AOI21XL U225 ( .A0(N920), .A1(n200), .B0(n259), .Y(n1693) );
  OAI21X1 U226 ( .A0(n164), .A1(n827), .B0(n1756), .Y(n2801) );
  OAI221XL U227 ( .A0(n304), .A1(n1153), .B0(n191), .B1(n922), .C0(n1509), .Y(
        n2496) );
  AOI21XL U228 ( .A0(N1014), .A1(n202), .B0(n258), .Y(n1497) );
  AOI21XL U229 ( .A0(N1013), .A1(n717), .B0(n258), .Y(n1498) );
  AOI21XL U230 ( .A0(N1015), .A1(n200), .B0(n258), .Y(n1496) );
  AOI21X1 U231 ( .A0(N995), .A1(n204), .B0(n259), .Y(n1516) );
  AOI21XL U232 ( .A0(N968), .A1(n197), .B0(n259), .Y(n1628) );
  AOI21XL U233 ( .A0(N994), .A1(n204), .B0(n259), .Y(n1517) );
  AOI21XL U234 ( .A0(N969), .A1(n204), .B0(n259), .Y(n1627) );
  AOI21XL U235 ( .A0(SHA256_result[124]), .A1(n179), .B0(n262), .Y(n458) );
  AOI21XL U236 ( .A0(n83), .A1(n179), .B0(n262), .Y(n416) );
  AOI21XL U237 ( .A0(n184), .A1(SHA256_result[120]), .B0(n258), .Y(n473) );
  AOI21XL U238 ( .A0(SHA256_result[37]), .A1(n184), .B0(n262), .Y(n404) );
  AOI21XL U239 ( .A0(n184), .A1(SHA256_result[113]), .B0(n261), .Y(n488) );
  AOI21XL U240 ( .A0(n135), .A1(n181), .B0(n256), .Y(n636) );
  AOI21XL U241 ( .A0(n157), .A1(n179), .B0(n256), .Y(n708) );
  AOI21XL U242 ( .A0(n183), .A1(n143), .B0(n256), .Y(n661) );
  NAND2BX1 U243 ( .AN(n24), .B(first_block), .Y(n1437) );
  OAI211X1 U244 ( .A0(n22), .A1(n455), .B0(n58), .C0(n1582), .Y(n2610) );
  OAI211X1 U245 ( .A0(n23), .A1(n944), .B0(n54), .C0(n1451), .Y(n2443) );
  BUFX16 U246 ( .A(T1_32[13]), .Y(n45) );
  NAND2X4 U247 ( .A(N1049), .B(n202), .Y(n100) );
  CLKINVX3 U248 ( .A(SHA256_result[40]), .Y(n915) );
  AOI2BB2X4 U249 ( .B0(N890), .B1(n202), .A0N(n798), .A1N(n280), .Y(n1723) );
  OAI2BB2XL U250 ( .B0(n342), .B1(n1156), .A0N(H5[12]), .A1N(n227), .Y(n2658)
         );
  OAI221XL U251 ( .A0(n304), .A1(n1156), .B0(n192), .B1(n919), .C0(n1512), .Y(
        n2499) );
  AOI2BB2X4 U252 ( .B0(N1050), .B1(n197), .A0N(n938), .A1N(n279), .Y(n1454) );
  INVX4 U253 ( .A(next_E[18]), .Y(n46) );
  NAND2BX2 U254 ( .AN(n1849), .B(output_enable), .Y(n1491) );
  CLKINVX3 U255 ( .A(n173), .Y(n166) );
  INVX1 U256 ( .A(n174), .Y(n173) );
  OAI2BB1X4 U257 ( .A0N(n198), .A1N(N954), .B0(n552), .Y(n2703) );
  INVXL U258 ( .A(next_E[9]), .Y(n513) );
  INVX1 U259 ( .A(n717), .Y(n48) );
  INVX1 U260 ( .A(n204), .Y(n49) );
  INVX4 U261 ( .A(n716), .Y(n721) );
  INVX1 U262 ( .A(n207), .Y(n205) );
  OR2XL U263 ( .A(n389), .B(n111), .Y(n716) );
  INVX1 U264 ( .A(n721), .Y(n207) );
  OAI221XL U265 ( .A0(n304), .A1(n1154), .B0(n190), .B1(n921), .C0(n1510), .Y(
        n2497) );
  OAI22XL U266 ( .A0(n1985), .A1(n445), .B0(n246), .B1(n72), .Y(n354) );
  OAI2BB2X1 U267 ( .B0(n342), .B1(n1160), .A0N(H5[8]), .A1N(n226), .Y(n2662)
         );
  MXI2X4 U268 ( .A(n922), .B(n1153), .S0(SHA256_result[111]), .Y(f1_EFG_32[15]) );
  OAI2BB2XL U269 ( .B0(n342), .B1(n1153), .A0N(H5[15]), .A1N(n227), .Y(n2655)
         );
  NAND3X4 U270 ( .A(n448), .B(n449), .C(n450), .Y(n2704) );
  NAND2X4 U271 ( .A(N953), .B(n203), .Y(n448) );
  NAND2XL U272 ( .A(n442), .B(SHA256_result[100]), .Y(n77) );
  INVX4 U273 ( .A(SHA256_result[68]), .Y(n442) );
  NAND2XL U274 ( .A(H7[0]), .B(n223), .Y(n1453) );
  INVX12 U275 ( .A(n1437), .Y(n53) );
  MXI2X4 U276 ( .A(n924), .B(n1151), .S0(SHA256_result[113]), .Y(f1_EFG_32[17]) );
  INVXL U277 ( .A(next_A[7]), .Y(n688) );
  XOR3X4 U278 ( .A(n155), .B(n144), .C(n136), .Y(f3_A_32[2]) );
  CLKINVX2 U279 ( .A(n70), .Y(n63) );
  INVX4 U280 ( .A(n64), .Y(n65) );
  CLKINVX2 U281 ( .A(n64), .Y(n66) );
  INVX4 U282 ( .A(n68), .Y(n69) );
  AOI22X2 U283 ( .A0(N985), .A1(n717), .B0(SHA256_result[126]), .B1(n273), .Y(
        n1611) );
  NOR2X1 U284 ( .A(n345), .B(n161), .Y(n113) );
  AND2X2 U285 ( .A(N889), .B(n203), .Y(n106) );
  OAI21X1 U286 ( .A0(n156), .A1(SHA256_result[195]), .B0(SHA256_result[163]), 
        .Y(n612) );
  INVXL U287 ( .A(n447), .Y(n75) );
  OAI211X2 U288 ( .A0(n283), .A1(n550), .B0(n439), .C0(n438), .Y(n2671) );
  NAND2X4 U289 ( .A(N986), .B(n196), .Y(n438) );
  NAND2XL U290 ( .A(n1163), .B(SHA256_result[101]), .Y(n86) );
  CLKINVX8 U291 ( .A(n87), .Y(f1_EFG_32[5]) );
  OAI2BB2X1 U292 ( .B0(n342), .B1(n857), .A0N(H3[0]), .A1N(n226), .Y(n2606) );
  AND2X4 U293 ( .A(n122), .B(n677), .Y(n1755) );
  NAND2X4 U294 ( .A(N858), .B(n198), .Y(n122) );
  OAI2BB2XL U295 ( .B0(n342), .B1(n941), .A0N(H7[1]), .A1N(n227), .Y(n2446) );
  OR2XL U296 ( .A(n162), .B(n936), .Y(n93) );
  AND2X4 U297 ( .A(n118), .B(n119), .Y(n1493) );
  OAI211XL U298 ( .A0(n19), .A1(n565), .B0(n59), .C0(n1561), .Y(n2574) );
  INVX1 U299 ( .A(n328), .Y(n311) );
  INVX1 U300 ( .A(n400), .Y(n1457) );
  INVX1 U301 ( .A(SHA256_result[62]), .Y(n937) );
  NAND2X4 U302 ( .A(N1018), .B(n199), .Y(n118) );
  AND2X4 U303 ( .A(n100), .B(n677), .Y(n1458) );
  NAND2XL U304 ( .A(n99), .B(n221), .Y(n570) );
  INVXL U305 ( .A(n174), .Y(n172) );
  NAND2X1 U306 ( .A(n101), .B(n1494), .Y(n2481) );
  NAND2X1 U307 ( .A(N1017), .B(n200), .Y(n102) );
  NAND2X1 U308 ( .A(SHA256_result[94]), .B(n274), .Y(n103) );
  AND2X2 U309 ( .A(n102), .B(n103), .Y(n1494) );
  OR2XL U310 ( .A(n162), .B(n937), .Y(n101) );
  INVX1 U311 ( .A(n280), .Y(n270) );
  INVX1 U312 ( .A(n280), .Y(n271) );
  INVX2 U313 ( .A(n173), .Y(n165) );
  NAND2X1 U314 ( .A(n393), .B(n1491), .Y(n715) );
  INVX1 U315 ( .A(SHA256_result[55]), .Y(n930) );
  OAI2BB1X1 U316 ( .A0N(n80), .A1N(n66), .B0(n614), .Y(f2_ABC_32[1]) );
  OAI21XL U317 ( .A0(n80), .A1(n66), .B0(SHA256_result[161]), .Y(n614) );
  OR2X2 U318 ( .A(n165), .B(n855), .Y(n104) );
  INVX1 U319 ( .A(n279), .Y(n272) );
  NOR2XL U320 ( .A(n113), .B(n2138), .Y(n2396) );
  NAND2X1 U321 ( .A(N809), .B(n201), .Y(n666) );
  NAND2X1 U322 ( .A(N808), .B(n202), .Y(n669) );
  NOR2X1 U323 ( .A(n166), .B(n468), .Y(n469) );
  NAND2X1 U324 ( .A(N807), .B(n200), .Y(n672) );
  NAND2XL U325 ( .A(n169), .B(n147), .Y(n673) );
  NAND2X1 U326 ( .A(N804), .B(n205), .Y(n681) );
  AOI21XL U327 ( .A0(n184), .A1(n153), .B0(n256), .Y(n689) );
  AOI21XL U328 ( .A0(n154), .A1(n179), .B0(n256), .Y(n693) );
  INVXL U329 ( .A(n116), .Y(n793) );
  AOI211XL U330 ( .A0(n761), .A1(round[2]), .B0(n2214), .C0(n2215), .Y(n2213)
         );
  AOI221XL U331 ( .A0(n2144), .A1(round[1]), .B0(n113), .B1(n31), .C0(n2215), 
        .Y(n2260) );
  AOI211XL U332 ( .A0(n761), .A1(n116), .B0(n2163), .C0(n2164), .Y(n2153) );
  AOI21XL U333 ( .A0(n116), .A1(n2350), .B0(n2151), .Y(n2156) );
  INVXL U334 ( .A(SHA256_result[33]), .Y(n447) );
  AOI21XL U335 ( .A0(n184), .A1(SHA256_result[114]), .B0(n262), .Y(n486) );
  AOI21XL U336 ( .A0(n184), .A1(SHA256_result[115]), .B0(n262), .Y(n483) );
  AOI22X1 U337 ( .A0(N882), .A1(n717), .B0(SHA256_result[215]), .B1(n270), .Y(
        n1731) );
  OAI2BB2X1 U338 ( .B0(n342), .B1(n802), .A0N(H1[5]), .A1N(n212), .Y(n2858) );
  OAI2BB2X1 U339 ( .B0(n342), .B1(n800), .A0N(H1[3]), .A1N(n219), .Y(n2860) );
  NAND2X1 U340 ( .A(N937), .B(n197), .Y(n494) );
  AOI21XL U341 ( .A0(n183), .A1(SHA256_result[110]), .B0(n258), .Y(n495) );
  BUFX4 U342 ( .A(SHA256_result[228]), .Y(n155) );
  AOI22X1 U343 ( .A0(N912), .A1(n198), .B0(SHA256_result[181]), .B1(n271), .Y(
        n1701) );
  AOI22X1 U344 ( .A0(N879), .A1(n204), .B0(SHA256_result[212]), .B1(n270), .Y(
        n1734) );
  AOI22X1 U345 ( .A0(N911), .A1(n206), .B0(SHA256_result[180]), .B1(n271), .Y(
        n1702) );
  OAI2BB2X1 U346 ( .B0(n342), .B1(n801), .A0N(H1[4]), .A1N(n216), .Y(n2859) );
  AOI22XL U347 ( .A0(next_E[12]), .A1(n269), .B0(N935), .B1(n201), .Y(n500) );
  OAI21XL U348 ( .A0(SHA256_result[202]), .A1(n149), .B0(SHA256_result[170]), 
        .Y(n605) );
  BUFX8 U349 ( .A(SHA256_result[254]), .Y(n131) );
  BUFX3 U350 ( .A(n344), .Y(n161) );
  AOI222XL U351 ( .A0(n113), .A1(n2122), .B0(n2195), .B1(n1393), .C0(n2304), 
        .C1(n1396), .Y(n2357) );
  AOI211XL U352 ( .A0(n2397), .A1(n116), .B0(n2323), .C0(n2325), .Y(n2392) );
  NAND2X1 U353 ( .A(n108), .B(n1692), .Y(n2736) );
  NAND2X1 U354 ( .A(N921), .B(n203), .Y(n109) );
  AND2X2 U355 ( .A(n109), .B(n110), .Y(n1692) );
  OR2XL U356 ( .A(n165), .B(n854), .Y(n105) );
  AND2X1 U357 ( .A(SHA256_result[222]), .B(n270), .Y(n107) );
  OR2X2 U358 ( .A(n165), .B(n887), .Y(n108) );
  NAND2XL U359 ( .A(SHA256_result[190]), .B(n271), .Y(n110) );
  INVX1 U360 ( .A(n187), .Y(n178) );
  INVX1 U361 ( .A(n186), .Y(n176) );
  INVX1 U362 ( .A(n677), .Y(n259) );
  NOR2XL U363 ( .A(n166), .B(n638), .Y(n639) );
  NAND2XL U364 ( .A(n1490), .B(n1491), .Y(n400) );
  INVXL U365 ( .A(n1456), .Y(n268) );
  AOI222XL U366 ( .A0(n2304), .A1(n2135), .B0(n2286), .B1(n2305), .C0(n2306), 
        .C1(n32), .Y(n2298) );
  NAND2XL U367 ( .A(n113), .B(n2378), .Y(n2184) );
  AOI21XL U368 ( .A0(n182), .A1(n144), .B0(n256), .Y(n664) );
  AOI21XL U369 ( .A0(n182), .A1(n145), .B0(n256), .Y(n667) );
  AOI21XL U370 ( .A0(n182), .A1(n140), .B0(n256), .Y(n654) );
  AOI21XL U371 ( .A0(n181), .A1(n146), .B0(n256), .Y(n670) );
  NAND2BX4 U372 ( .AN(n1859), .B(round[6]), .Y(n388) );
  AOI21XL U373 ( .A0(next_E[31]), .A1(n276), .B0(n551), .Y(n552) );
  AOI21XL U374 ( .A0(n183), .A1(n131), .B0(n256), .Y(n620) );
  NAND2X2 U375 ( .A(N824), .B(n198), .Y(n621) );
  NAND3X2 U376 ( .A(n623), .B(n622), .C(n621), .Y(n2866) );
  AOI21XL U377 ( .A0(n182), .A1(n132), .B0(n128), .Y(n623) );
  AOI21XL U378 ( .A0(next_A[31]), .A1(n276), .B0(n616), .Y(n617) );
  AOI21XL U379 ( .A0(N877), .A1(n195), .B0(n261), .Y(n1736) );
  AOI21XL U380 ( .A0(N876), .A1(n717), .B0(n261), .Y(n1737) );
  AOI21XL U381 ( .A0(N874), .A1(n717), .B0(n261), .Y(n1739) );
  AOI21XL U382 ( .A0(N873), .A1(n200), .B0(n257), .Y(n1740) );
  AOI21XL U383 ( .A0(N871), .A1(n198), .B0(n256), .Y(n1742) );
  AOI21XL U384 ( .A0(N868), .A1(n204), .B0(n259), .Y(n1745) );
  AOI21XL U385 ( .A0(N837), .A1(n202), .B0(n262), .Y(n1776) );
  AOI21XL U386 ( .A0(N836), .A1(n198), .B0(n262), .Y(n1777) );
  AOI21XL U387 ( .A0(N973), .A1(n206), .B0(n259), .Y(n1623) );
  AOI21XL U388 ( .A0(N867), .A1(n717), .B0(n257), .Y(n1746) );
  AOI21XL U389 ( .A0(N845), .A1(n721), .B0(n262), .Y(n1768) );
  AOI21XL U390 ( .A0(N844), .A1(n200), .B0(n262), .Y(n1769) );
  AOI21XL U391 ( .A0(N843), .A1(n206), .B0(n262), .Y(n1770) );
  AOI21XL U392 ( .A0(N842), .A1(n197), .B0(n262), .Y(n1771) );
  AOI21XL U393 ( .A0(N840), .A1(n196), .B0(n262), .Y(n1773) );
  AOI21XL U394 ( .A0(N838), .A1(n198), .B0(n262), .Y(n1775) );
  AOI21XL U395 ( .A0(N1040), .A1(n195), .B0(n257), .Y(n1468) );
  AOI21XL U396 ( .A0(N1030), .A1(n721), .B0(n257), .Y(n1478) );
  AOI21XL U397 ( .A0(n182), .A1(n150), .B0(n256), .Y(n680) );
  INVXL U398 ( .A(next_A[6]), .Y(n691) );
  INVXL U399 ( .A(next_A[5]), .Y(n695) );
  INVXL U400 ( .A(next_A[1]), .Y(n714) );
  NAND2XL U401 ( .A(N796), .B(n197), .Y(n713) );
  AOI21XL U402 ( .A0(n66), .A1(n184), .B0(n256), .Y(n712) );
  AOI22XL U403 ( .A0(next_A[0]), .A1(n269), .B0(n158), .B1(n179), .Y(n719) );
  AOI21XL U404 ( .A0(N795), .A1(n195), .B0(n257), .Y(n718) );
  OR2XL U405 ( .A(n1849), .B(n388), .Y(n111) );
  AOI22XL U406 ( .A0(N839), .A1(n205), .B0(n147), .B1(n269), .Y(n1774) );
  AOI22XL U407 ( .A0(N835), .A1(n721), .B0(n151), .B1(n269), .Y(n1778) );
  AOI22XL U408 ( .A0(N833), .A1(n203), .B0(n153), .B1(n269), .Y(n1780) );
  AOI22XL U409 ( .A0(N832), .A1(n206), .B0(n154), .B1(n271), .Y(n1781) );
  AOI22XL U410 ( .A0(N830), .A1(n202), .B0(n156), .B1(n269), .Y(n1783) );
  AOI2BB2XL U411 ( .B0(N894), .B1(n203), .A0N(n323), .A1N(n558), .Y(n553) );
  AOI2BB2XL U412 ( .B0(N892), .B1(n203), .A0N(n324), .A1N(n565), .Y(n555) );
  AOI2BB2XL U413 ( .B0(N849), .B1(n203), .A0N(n323), .A1N(n646), .Y(n578) );
  AOI2BB2XL U414 ( .B0(N829), .B1(n202), .A0N(n281), .A1N(n707), .Y(n580) );
  INVX1 U415 ( .A(round[1]), .Y(n345) );
  INVXL U416 ( .A(next_A[4]), .Y(n700) );
  INVXL U417 ( .A(next_A[3]), .Y(n706) );
  NAND2BXL U418 ( .AN(n49), .B(N1023), .Y(n395) );
  NAND2BXL U419 ( .AN(n48), .B(N1019), .Y(n402) );
  INVX1 U420 ( .A(n130), .Y(n233) );
  AOI222XL U421 ( .A0(n2276), .A1(n1396), .B0(n2185), .B1(n114), .C0(n2277), 
        .C1(n32), .Y(n2270) );
  AOI31XL U422 ( .A0(n781), .A1(n1393), .A2(n2226), .B0(n1878), .Y(n2211) );
  AOI22XL U423 ( .A0(n2202), .A1(n112), .B0(n2138), .B1(n2148), .Y(n2204) );
  AOI211XL U424 ( .A0(n2342), .A1(n32), .B0(n2373), .C0(n2414), .Y(n2411) );
  AOI22XL U425 ( .A0(n116), .A1(n2252), .B0(n2363), .B1(n161), .Y(n2405) );
  AOI222XL U426 ( .A0(n2356), .A1(n32), .B0(n2187), .B1(n41), .C0(n2176), .C1(
        n112), .Y(n2388) );
  AOI222XL U427 ( .A0(n2190), .A1(round[2]), .B0(n2185), .B1(n32), .C0(n2189), 
        .C1(n747), .Y(n2382) );
  AOI211XL U428 ( .A0(n2268), .A1(n116), .B0(n2283), .C0(n2348), .Y(n2344) );
  AOI222XL U429 ( .A0(n2221), .A1(n114), .B0(n2324), .B1(n113), .C0(n2315), 
        .C1(n41), .Y(n2317) );
  AOI222XL U430 ( .A0(n782), .A1(n161), .B0(n2315), .B1(n32), .C0(n2247), .C1(
        n160), .Y(n2307) );
  AOI222XL U431 ( .A0(n2304), .A1(n345), .B0(n2287), .B1(n112), .C0(n2314), 
        .C1(n2268), .Y(n2308) );
  NOR2X1 U432 ( .A(n161), .B(n347), .Y(n112) );
  NOR2XL U433 ( .A(n345), .B(n343), .Y(n2135) );
  OAI32XL U434 ( .A0(n781), .A1(round[1]), .A2(n797), .B0(round[2]), .B1(n2244), .Y(n2243) );
  AOI31XL U435 ( .A0(n795), .A1(n753), .A2(n762), .B0(n32), .Y(n2340) );
  AOI21XL U436 ( .A0(round[2]), .A1(n113), .B0(n2124), .Y(n2118) );
  AOI31XL U437 ( .A0(n160), .A1(round[2]), .A2(n113), .B0(n2404), .Y(n2403) );
  NOR2X1 U438 ( .A(n346), .B(n160), .Y(n114) );
  NOR2XL U439 ( .A(n343), .B(n797), .Y(n2187) );
  AOI21XL U440 ( .A0(n792), .A1(n2173), .B0(n345), .Y(n2303) );
  INVX1 U441 ( .A(n247), .Y(n246) );
  NAND2XL U442 ( .A(n116), .B(n160), .Y(n2146) );
  NOR2XL U443 ( .A(n345), .B(n160), .Y(n2268) );
  OAI2BB1X4 U444 ( .A0N(n387), .A1N(n348), .B0(n1434), .Y(n1849) );
  OAI211XL U445 ( .A0(n17), .A1(n951), .B0(n59), .C0(n1448), .Y(n2436) );
  NAND2XL U446 ( .A(H7[11]), .B(n223), .Y(n1448) );
  OAI211XL U447 ( .A0(n23), .A1(n950), .B0(n55), .C0(n1449), .Y(n2437) );
  NAND2XL U448 ( .A(H7[10]), .B(n223), .Y(n1449) );
  OAI211XL U449 ( .A0(n17), .A1(n948), .B0(n58), .C0(n1450), .Y(n2439) );
  NAND2XL U450 ( .A(H7[8]), .B(n223), .Y(n1450) );
  NAND2XL U451 ( .A(H7[4]), .B(n223), .Y(n1451) );
  OAI211XL U452 ( .A0(n24), .A1(n441), .B0(n55), .C0(n1538), .Y(n2537) );
  NAND2XL U453 ( .A(H6[5]), .B(n221), .Y(n1538) );
  OAI211XL U454 ( .A0(n24), .A1(n856), .B0(n58), .C0(n1562), .Y(n2575) );
  OAI211XL U455 ( .A0(n18), .A1(n798), .B0(n55), .C0(n1787), .Y(n2832) );
  OAI211XL U456 ( .A0(n17), .A1(n943), .B0(n58), .C0(n1452), .Y(n2444) );
  NAND2XL U457 ( .A(H7[3]), .B(n223), .Y(n1452) );
  NAND2XL U458 ( .A(H6[28]), .B(n224), .Y(n1524) );
  OAI211XL U459 ( .A0(n17), .A1(n918), .B0(n55), .C0(n1535), .Y(n2531) );
  NAND2XL U460 ( .A(H6[11]), .B(n221), .Y(n1535) );
  OAI211XL U461 ( .A0(n22), .A1(n915), .B0(n59), .C0(n1536), .Y(n2534) );
  NAND2XL U462 ( .A(H6[8]), .B(n221), .Y(n1536) );
  OAI211XL U463 ( .A0(n18), .A1(n914), .B0(n54), .C0(n1537), .Y(n2535) );
  NAND2XL U464 ( .A(H6[7]), .B(n221), .Y(n1537) );
  OAI211XL U465 ( .A0(n18), .A1(n1161), .B0(n60), .C0(n1607), .Y(n2663) );
  NAND2XL U466 ( .A(H5[7]), .B(n214), .Y(n1607) );
  OAI211XL U467 ( .A0(n17), .A1(n1165), .B0(n54), .C0(n1608), .Y(n2667) );
  OAI211XL U468 ( .A0(n24), .A1(n867), .B0(n56), .C0(n1575), .Y(n2596) );
  NAND2XL U469 ( .A(H3[10]), .B(n217), .Y(n1575) );
  OAI211XL U470 ( .A0(n21), .A1(n865), .B0(n55), .C0(n1576), .Y(n2598) );
  OAI211XL U471 ( .A0(n17), .A1(n862), .B0(n56), .C0(n1577), .Y(n2601) );
  OAI211XL U472 ( .A0(n17), .A1(n861), .B0(n57), .C0(n1578), .Y(n2602) );
  OAI211XL U473 ( .A0(n17), .A1(n860), .B0(n57), .C0(n1579), .Y(n2603) );
  NAND2XL U474 ( .A(H3[3]), .B(n216), .Y(n1579) );
  OAI211XL U475 ( .A0(n21), .A1(n858), .B0(n60), .C0(n1580), .Y(n2605) );
  OAI211XL U476 ( .A0(n21), .A1(n833), .B0(n60), .C0(n1556), .Y(n2566) );
  OAI211XL U477 ( .A0(n20), .A1(n832), .B0(n60), .C0(n1557), .Y(n2567) );
  NAND2XL U478 ( .A(H2[8]), .B(n218), .Y(n1557) );
  OAI211XL U479 ( .A0(n20), .A1(n830), .B0(n54), .C0(n1558), .Y(n2569) );
  OAI211XL U480 ( .A0(n24), .A1(n829), .B0(n61), .C0(n1559), .Y(n2570) );
  OAI211XL U481 ( .A0(n23), .A1(n828), .B0(n54), .C0(n1560), .Y(n2571) );
  NAND2XL U482 ( .A(H2[1]), .B(n218), .Y(n1561) );
  OAI211XL U483 ( .A0(n17), .A1(n808), .B0(n54), .C0(n1800), .Y(n2852) );
  NAND2XL U484 ( .A(H1[11]), .B(n213), .Y(n1800) );
  OAI211XL U485 ( .A0(n18), .A1(n807), .B0(n57), .C0(n1801), .Y(n2853) );
  OAI211XL U486 ( .A0(n22), .A1(n806), .B0(n61), .C0(n1802), .Y(n2854) );
  NAND2XL U487 ( .A(H1[9]), .B(n213), .Y(n1802) );
  OAI211XL U488 ( .A0(n19), .A1(n804), .B0(n62), .C0(n1803), .Y(n2856) );
  NAND2XL U489 ( .A(H1[7]), .B(n213), .Y(n1803) );
  OAI211XL U490 ( .A0(n17), .A1(n799), .B0(n58), .C0(n1804), .Y(n2861) );
  NAND2XL U491 ( .A(H1[0]), .B(n213), .Y(n1805) );
  NAND3XL U492 ( .A(n115), .B(n60), .C(n1873), .Y(n2922) );
  OR2XL U493 ( .A(n22), .B(n692), .Y(n115) );
  NAND3BXL U494 ( .AN(n711), .B(n59), .C(n1875), .Y(n2926) );
  NAND2XL U495 ( .A(H5[2]), .B(n214), .Y(n1609) );
  INVXL U496 ( .A(n155), .Y(n697) );
  INVXL U497 ( .A(n156), .Y(n702) );
  NAND2XL U498 ( .A(H2[3]), .B(n221), .Y(n557) );
  INVXL U499 ( .A(SHA256_result[162]), .Y(n562) );
  NAND2XL U500 ( .A(H2[2]), .B(n221), .Y(n561) );
  INVXL U501 ( .A(SHA256_result[160]), .Y(n571) );
  AOI22XL U502 ( .A0(N984), .A1(n721), .B0(n51), .B1(n273), .Y(n1612) );
  OAI211XL U503 ( .A0(n19), .A1(n444), .B0(n58), .C0(n1539), .Y(n2539) );
  NAND2XL U504 ( .A(H6[3]), .B(n220), .Y(n1539) );
  NAND2XL U505 ( .A(n96), .B(n220), .Y(n1540) );
  OAI211XL U506 ( .A0(n21), .A1(n81), .B0(n57), .C0(n1541), .Y(n2542) );
  NAND2XL U507 ( .A(H6[0]), .B(n220), .Y(n1541) );
  OAI211XL U508 ( .A0(n22), .A1(n440), .B0(n55), .C0(n1581), .Y(n2608) );
  OAI211XL U509 ( .A0(n23), .A1(n510), .B0(n56), .C0(n1589), .Y(n2629) );
  OAI211XL U510 ( .A0(n20), .A1(n524), .B0(n56), .C0(n1590), .Y(n2632) );
  OAI2BB2XL U511 ( .B0(n342), .B1(n949), .A0N(H7[9]), .A1N(n227), .Y(n2438) );
  OAI2BB2XL U512 ( .B0(n342), .B1(n947), .A0N(H7[7]), .A1N(n227), .Y(n2440) );
  OAI2BB2XL U513 ( .B0(n342), .B1(n946), .A0N(H7[6]), .A1N(n227), .Y(n2441) );
  OAI2BB2XL U514 ( .B0(n342), .B1(n945), .A0N(H7[5]), .A1N(n225), .Y(n2442) );
  OAI2BB2XL U515 ( .B0(n342), .B1(n917), .A0N(H6[10]), .A1N(n225), .Y(n2532)
         );
  OAI2BB2XL U516 ( .B0(n342), .B1(n916), .A0N(H6[9]), .A1N(n215), .Y(n2533) );
  OAI2BB2XL U517 ( .B0(n342), .B1(n913), .A0N(H6[6]), .A1N(n217), .Y(n2536) );
  OAI2BB2XL U518 ( .B0(n342), .B1(n904), .A0N(H5[10]), .A1N(n226), .Y(n2660)
         );
  OAI2BB2XL U519 ( .B0(n342), .B1(n903), .A0N(H5[9]), .A1N(n226), .Y(n2661) );
  OAI2BB2XL U520 ( .B0(n342), .B1(n902), .A0N(H5[6]), .A1N(n226), .Y(n2664) );
  OAI2BB2XL U521 ( .B0(n342), .B1(n1163), .A0N(H5[5]), .A1N(n226), .Y(n2665)
         );
  OAI2BB2XL U522 ( .B0(n342), .B1(n868), .A0N(H3[11]), .A1N(n225), .Y(n2595)
         );
  OAI2BB2XL U523 ( .B0(n342), .B1(n866), .A0N(H3[9]), .A1N(n225), .Y(n2597) );
  OAI2BB2XL U524 ( .B0(n342), .B1(n864), .A0N(H3[7]), .A1N(n225), .Y(n2599) );
  OAI2BB2XL U525 ( .B0(n342), .B1(n863), .A0N(H3[6]), .A1N(n225), .Y(n2600) );
  OAI2BB2XL U526 ( .B0(n342), .B1(n805), .A0N(H1[8]), .A1N(n225), .Y(n2855) );
  OAI2BB2XL U527 ( .B0(n342), .B1(n803), .A0N(H1[6]), .A1N(n222), .Y(n2857) );
  OAI2BB2XL U528 ( .B0(n342), .B1(n738), .A0N(H0[21]), .A1N(n221), .Y(n2906)
         );
  OAI2BB2XL U529 ( .B0(n342), .B1(n737), .A0N(H0[20]), .A1N(n213), .Y(n2907)
         );
  OAI2BB2XL U530 ( .B0(n342), .B1(n735), .A0N(H0[18]), .A1N(n215), .Y(n2909)
         );
  AOI21XL U531 ( .A0(n185), .A1(SHA256_result[95]), .B0(n260), .Y(n439) );
  AOI2BB2XL U532 ( .B0(n169), .B1(SHA256_result[117]), .A0N(n324), .A1N(n478), 
        .Y(n479) );
  AOI2BB2XL U533 ( .B0(SHA256_result[107]), .B1(n169), .A0N(n324), .A1N(n503), 
        .Y(n504) );
  AOI21XL U534 ( .A0(N1012), .A1(n195), .B0(n258), .Y(n1499) );
  AOI21XL U535 ( .A0(N1011), .A1(n199), .B0(n258), .Y(n1500) );
  AOI21XL U536 ( .A0(N1010), .A1(n204), .B0(n258), .Y(n1501) );
  AOI21XL U537 ( .A0(N1002), .A1(n197), .B0(n258), .Y(n1509) );
  AOI21XL U538 ( .A0(N1001), .A1(n195), .B0(n258), .Y(n1510) );
  AOI21XL U539 ( .A0(N999), .A1(n195), .B0(n259), .Y(n1512) );
  AOI21XL U540 ( .A0(N998), .A1(n195), .B0(n259), .Y(n1513) );
  AOI21XL U541 ( .A0(N971), .A1(n717), .B0(n259), .Y(n1625) );
  INVX4 U542 ( .A(SHA256_result[43]), .Y(n918) );
  CLKBUFX8 U543 ( .A(SHA256_result[237]), .Y(n146) );
  CLKBUFX8 U544 ( .A(SHA256_result[249]), .Y(n135) );
  CLKBUFX8 U545 ( .A(SHA256_result[239]), .Y(n144) );
  CLKBUFX8 U546 ( .A(SHA256_result[251]), .Y(n133) );
  NAND2XL U547 ( .A(H6[4]), .B(n219), .Y(n406) );
  NAND2XL U548 ( .A(H5[4]), .B(n219), .Y(n431) );
  NAND2XL U549 ( .A(H6[2]), .B(n219), .Y(n411) );
  OAI211XL U550 ( .A0(n1168), .A1(n321), .B0(n417), .C0(n416), .Y(n2543) );
  NAND2XL U551 ( .A(N987), .B(n202), .Y(n417) );
  NAND2XL U552 ( .A(N988), .B(n717), .Y(n415) );
  AOI21XL U553 ( .A0(n75), .A1(n179), .B0(n259), .Y(n414) );
  INVXL U554 ( .A(next_E[6]), .Y(n527) );
  INVXL U555 ( .A(next_E[2]), .Y(n541) );
  INVXL U556 ( .A(next_E[1]), .Y(n545) );
  INVXL U557 ( .A(next_E[4]), .Y(n534) );
  AOI21XL U558 ( .A0(SHA256_result[100]), .A1(n180), .B0(n256), .Y(n532) );
  NAND2XL U559 ( .A(N990), .B(n197), .Y(n410) );
  NAND2XL U560 ( .A(N860), .B(n201), .Y(n567) );
  AOI21XL U561 ( .A0(SHA256_result[161]), .A1(n183), .B0(n261), .Y(n566) );
  INVXL U562 ( .A(next_E[5]), .Y(n530) );
  NAND2XL U563 ( .A(N928), .B(n197), .Y(n529) );
  AOI21XL U564 ( .A0(SHA256_result[101]), .A1(n181), .B0(n257), .Y(n528) );
  AOI2BB2XL U565 ( .B0(n168), .B1(SHA256_result[112]), .A0N(n324), .A1N(n490), 
        .Y(n491) );
  AOI2BB2XL U566 ( .B0(n169), .B1(SHA256_result[116]), .A0N(n323), .A1N(n480), 
        .Y(n481) );
  NAND2BXL U567 ( .AN(n310), .B(SHA256_result[124]), .Y(n419) );
  NAND2BXL U568 ( .AN(n314), .B(SHA256_result[123]), .Y(n422) );
  MXI2XL U569 ( .A(n930), .B(n1145), .S0(SHA256_result[119]), .Y(f1_EFG_32[23]) );
  AOI22XL U570 ( .A0(N875), .A1(n200), .B0(SHA256_result[208]), .B1(n270), .Y(
        n1738) );
  AOI22XL U571 ( .A0(N869), .A1(n200), .B0(SHA256_result[202]), .B1(n270), .Y(
        n1744) );
  AOI22XL U572 ( .A0(N866), .A1(n199), .B0(SHA256_result[199]), .B1(n270), .Y(
        n1747) );
  AOI22XL U573 ( .A0(N1008), .A1(n721), .B0(SHA256_result[85]), .B1(n273), .Y(
        n1503) );
  AOI22XL U574 ( .A0(N1007), .A1(n204), .B0(SHA256_result[84]), .B1(n273), .Y(
        n1504) );
  AOI22XL U575 ( .A0(N1006), .A1(n202), .B0(SHA256_result[83]), .B1(n273), .Y(
        n1505) );
  AOI22XL U576 ( .A0(N1005), .A1(n201), .B0(SHA256_result[82]), .B1(n273), .Y(
        n1506) );
  AOI22XL U577 ( .A0(N891), .A1(n196), .B0(SHA256_result[160]), .B1(n270), .Y(
        n1722) );
  AOI22XL U578 ( .A0(N1009), .A1(n203), .B0(SHA256_result[86]), .B1(n274), .Y(
        n1502) );
  AOI22XL U579 ( .A0(N902), .A1(n204), .B0(SHA256_result[171]), .B1(n271), .Y(
        n1711) );
  AOI22XL U580 ( .A0(N900), .A1(n202), .B0(SHA256_result[169]), .B1(n271), .Y(
        n1713) );
  AOI22XL U581 ( .A0(N897), .A1(n205), .B0(SHA256_result[166]), .B1(n271), .Y(
        n1716) );
  AOI22XL U582 ( .A0(N898), .A1(n199), .B0(SHA256_result[167]), .B1(n272), .Y(
        n1715) );
  AOI22XL U583 ( .A0(N961), .A1(n203), .B0(SHA256_result[102]), .B1(n272), .Y(
        n1635) );
  AOI22XL U584 ( .A0(N1000), .A1(n202), .B0(SHA256_result[77]), .B1(n273), .Y(
        n1511) );
  AOI22XL U585 ( .A0(N997), .A1(n199), .B0(SHA256_result[74]), .B1(n273), .Y(
        n1514) );
  AOI22XL U586 ( .A0(N996), .A1(n195), .B0(SHA256_result[73]), .B1(n273), .Y(
        n1515) );
  AOI22XL U587 ( .A0(N993), .A1(n197), .B0(SHA256_result[70]), .B1(n273), .Y(
        n1518) );
  AOI22XL U588 ( .A0(N977), .A1(n717), .B0(SHA256_result[118]), .B1(n273), .Y(
        n1619) );
  AOI22XL U589 ( .A0(N976), .A1(n199), .B0(SHA256_result[117]), .B1(n272), .Y(
        n1620) );
  AOI22XL U590 ( .A0(N975), .A1(n204), .B0(SHA256_result[116]), .B1(n272), .Y(
        n1621) );
  AOI22XL U591 ( .A0(N974), .A1(n197), .B0(SHA256_result[115]), .B1(n272), .Y(
        n1622) );
  AOI22XL U592 ( .A0(N955), .A1(n200), .B0(n63), .B1(n271), .Y(n1641) );
  AOI22XL U593 ( .A0(N970), .A1(n197), .B0(SHA256_result[111]), .B1(n272), .Y(
        n1626) );
  AOI22XL U594 ( .A0(N960), .A1(n204), .B0(SHA256_result[101]), .B1(n272), .Y(
        n1636) );
  AOI22XL U595 ( .A0(N963), .A1(n202), .B0(SHA256_result[104]), .B1(n272), .Y(
        n1633) );
  AOI22XL U596 ( .A0(N978), .A1(n204), .B0(SHA256_result[119]), .B1(n273), .Y(
        n1618) );
  AOI22XL U597 ( .A0(N972), .A1(n721), .B0(SHA256_result[113]), .B1(n272), .Y(
        n1624) );
  AOI22XL U598 ( .A0(N1020), .A1(n199), .B0(n75), .B1(n274), .Y(n1488) );
  AOI22XL U599 ( .A0(N1039), .A1(n196), .B0(SHA256_result[52]), .B1(n275), .Y(
        n1469) );
  AOI22XL U600 ( .A0(N1036), .A1(n204), .B0(SHA256_result[49]), .B1(n275), .Y(
        n1472) );
  AOI22XL U601 ( .A0(N1035), .A1(n204), .B0(SHA256_result[48]), .B1(n274), .Y(
        n1473) );
  AOI22XL U602 ( .A0(N1032), .A1(n198), .B0(SHA256_result[45]), .B1(n274), .Y(
        n1476) );
  AOI22XL U603 ( .A0(N1031), .A1(n202), .B0(SHA256_result[44]), .B1(n274), .Y(
        n1477) );
  AOI22XL U604 ( .A0(N1025), .A1(n201), .B0(n50), .B1(n274), .Y(n1483) );
  AOI22XL U605 ( .A0(N1038), .A1(n195), .B0(SHA256_result[51]), .B1(n275), .Y(
        n1470) );
  AOI22XL U606 ( .A0(N1037), .A1(n721), .B0(SHA256_result[50]), .B1(n275), .Y(
        n1471) );
  AOI22XL U607 ( .A0(N1028), .A1(n202), .B0(SHA256_result[41]), .B1(n274), .Y(
        n1480) );
  AOI22XL U608 ( .A0(N1024), .A1(n203), .B0(SHA256_result[37]), .B1(n274), .Y(
        n1484) );
  INVXL U609 ( .A(next_E[8]), .Y(n518) );
  INVXL U610 ( .A(next_E[7]), .Y(n523) );
  NAND2XL U611 ( .A(SHA256_result[160]), .B(n170), .Y(n569) );
  NAND2XL U612 ( .A(SHA256_result[68]), .B(n170), .Y(n433) );
  NAND2XL U613 ( .A(N959), .B(n721), .Y(n432) );
  NAND2XL U614 ( .A(SHA256_result[163]), .B(n170), .Y(n560) );
  NAND2XL U615 ( .A(N862), .B(n203), .Y(n559) );
  NAND2XL U616 ( .A(SHA256_result[162]), .B(n171), .Y(n564) );
  NAND2XL U617 ( .A(N861), .B(n196), .Y(n563) );
  NAND2XL U618 ( .A(SHA256_result[36]), .B(n170), .Y(n408) );
  NAND2XL U619 ( .A(N991), .B(n200), .Y(n407) );
  NAND2BXL U620 ( .AN(n265), .B(SHA256_result[121]), .Y(n425) );
  NAND2XL U621 ( .A(N980), .B(n201), .Y(n424) );
  AOI2BB2XL U622 ( .B0(N958), .B1(n203), .A0N(n321), .A1N(n535), .Y(n434) );
  AOI2BB2XL U623 ( .B0(N827), .B1(n202), .A0N(n322), .A1N(n720), .Y(n582) );
  AOI2BB2XL U624 ( .B0(N966), .B1(n195), .A0N(n322), .A1N(n502), .Y(n427) );
  AOI2BB2XL U625 ( .B0(N962), .B1(n206), .A0N(n325), .A1N(n520), .Y(n429) );
  MXI2XL U626 ( .A(n931), .B(n1144), .S0(SHA256_result[120]), .Y(f1_EFG_32[24]) );
  MXI2XL U627 ( .A(n934), .B(n1141), .S0(SHA256_result[123]), .Y(f1_EFG_32[27]) );
  MXI2XL U628 ( .A(n933), .B(n1142), .S0(SHA256_result[122]), .Y(f1_EFG_32[26]) );
  MXI2XL U629 ( .A(n935), .B(n1140), .S0(SHA256_result[124]), .Y(f1_EFG_32[28]) );
  MX2X1 U630 ( .A(SHA256_result[61]), .B(SHA256_result[93]), .S0(n51), .Y(
        f1_EFG_32[29]) );
  NOR3XL U631 ( .A(output_enable), .B(round[6]), .C(n1849), .Y(n129) );
  NAND2XL U632 ( .A(output_enable), .B(n1434), .Y(n1978) );
  AOI222XL U633 ( .A0(n2285), .A1(n345), .B0(n2286), .B1(n32), .C0(n2287), 
        .C1(n1396), .Y(n2278) );
  AOI31XL U634 ( .A0(n161), .A1(n1388), .A2(n2234), .B0(n2284), .Y(n2279) );
  AOI22XL U635 ( .A0(n2137), .A1(n345), .B0(n2259), .B1(n1370), .Y(n2253) );
  AOI221XL U636 ( .A0(n761), .A1(n1383), .B0(n2185), .B1(n160), .C0(n2186), 
        .Y(n2179) );
  AOI2BB2XL U637 ( .B0(n2177), .B1(round[2]), .A0N(n2166), .A1N(n1396), .Y(
        n2167) );
  AOI22XL U638 ( .A0(n237), .A1(n90), .B0(n235), .B1(n158), .Y(n2110) );
  AOI22XL U639 ( .A0(n242), .A1(SHA256_result[128]), .B0(n239), .B1(
        SHA256_result[160]), .Y(n2111) );
  AOI211XL U640 ( .A0(n249), .A1(n83), .B0(n350), .C0(n349), .Y(n2112) );
  AOI22XL U641 ( .A0(n237), .A1(n80), .B0(n235), .B1(n66), .Y(n2106) );
  AOI22XL U642 ( .A0(n237), .A1(SHA256_result[194]), .B0(n235), .B1(n157), .Y(
        n2102) );
  AOI22XL U643 ( .A0(n242), .A1(SHA256_result[130]), .B0(n239), .B1(
        SHA256_result[162]), .Y(n2103) );
  AOI22XL U644 ( .A0(n237), .A1(SHA256_result[195]), .B0(n235), .B1(n156), .Y(
        n2098) );
  AOI22XL U645 ( .A0(n242), .A1(SHA256_result[131]), .B0(n239), .B1(
        SHA256_result[163]), .Y(n2099) );
  AOI22XL U646 ( .A0(n237), .A1(SHA256_result[196]), .B0(n235), .B1(n155), .Y(
        n2094) );
  AOI22XL U647 ( .A0(n242), .A1(SHA256_result[132]), .B0(n239), .B1(
        SHA256_result[164]), .Y(n2095) );
  AOI211XL U648 ( .A0(n249), .A1(SHA256_result[36]), .B0(n358), .C0(n357), .Y(
        n2096) );
  AOI22XL U649 ( .A0(n237), .A1(SHA256_result[197]), .B0(n235), .B1(n154), .Y(
        n2090) );
  AOI22XL U650 ( .A0(n241), .A1(SHA256_result[133]), .B0(n239), .B1(
        SHA256_result[165]), .Y(n2091) );
  AOI211XL U651 ( .A0(n249), .A1(SHA256_result[37]), .B0(n360), .C0(n359), .Y(
        n2092) );
  AOI22XL U652 ( .A0(n237), .A1(SHA256_result[198]), .B0(n235), .B1(n153), .Y(
        n2086) );
  AOI22XL U653 ( .A0(n242), .A1(SHA256_result[134]), .B0(n239), .B1(
        SHA256_result[166]), .Y(n2087) );
  AOI211XL U654 ( .A0(n249), .A1(n50), .B0(n362), .C0(n361), .Y(n2088) );
  AOI22XL U655 ( .A0(n237), .A1(SHA256_result[199]), .B0(n235), .B1(n152), .Y(
        n2082) );
  AOI22XL U656 ( .A0(n241), .A1(SHA256_result[135]), .B0(n239), .B1(
        SHA256_result[167]), .Y(n2083) );
  AOI211XL U657 ( .A0(n249), .A1(SHA256_result[39]), .B0(n364), .C0(n363), .Y(
        n2084) );
  AOI22XL U658 ( .A0(n237), .A1(SHA256_result[200]), .B0(n235), .B1(n151), .Y(
        n2078) );
  AOI22XL U659 ( .A0(n1986), .A1(SHA256_result[136]), .B0(n239), .B1(
        SHA256_result[168]), .Y(n2079) );
  AOI211XL U660 ( .A0(n249), .A1(SHA256_result[40]), .B0(n366), .C0(n365), .Y(
        n2080) );
  AOI22XL U661 ( .A0(n237), .A1(SHA256_result[201]), .B0(n235), .B1(n150), .Y(
        n2074) );
  AOI22XL U662 ( .A0(n1986), .A1(SHA256_result[137]), .B0(n239), .B1(
        SHA256_result[169]), .Y(n2075) );
  AOI211XL U663 ( .A0(n249), .A1(SHA256_result[41]), .B0(n368), .C0(n367), .Y(
        n2076) );
  AOI22XL U664 ( .A0(n237), .A1(SHA256_result[202]), .B0(n235), .B1(n149), .Y(
        n2070) );
  AOI22XL U665 ( .A0(n1986), .A1(SHA256_result[138]), .B0(n239), .B1(
        SHA256_result[170]), .Y(n2071) );
  AOI211XL U666 ( .A0(n249), .A1(SHA256_result[42]), .B0(n370), .C0(n369), .Y(
        n2072) );
  AOI22XL U667 ( .A0(n237), .A1(SHA256_result[203]), .B0(n235), .B1(n148), .Y(
        n2066) );
  AOI22XL U668 ( .A0(n1986), .A1(SHA256_result[139]), .B0(n239), .B1(
        SHA256_result[171]), .Y(n2067) );
  AOI211XL U669 ( .A0(n248), .A1(SHA256_result[43]), .B0(n372), .C0(n371), .Y(
        n2068) );
  AOI22XL U670 ( .A0(n238), .A1(SHA256_result[204]), .B0(n236), .B1(n147), .Y(
        n2062) );
  AOI22XL U671 ( .A0(n241), .A1(SHA256_result[140]), .B0(n240), .B1(
        SHA256_result[172]), .Y(n2063) );
  AOI221XL U672 ( .A0(n254), .A1(SHA256_result[12]), .B0(n248), .B1(
        SHA256_result[44]), .C0(n2065), .Y(n2064) );
  AOI22XL U673 ( .A0(n238), .A1(SHA256_result[205]), .B0(n236), .B1(n146), .Y(
        n2058) );
  AOI22XL U674 ( .A0(n241), .A1(SHA256_result[141]), .B0(n240), .B1(
        SHA256_result[173]), .Y(n2059) );
  AOI22XL U675 ( .A0(n238), .A1(SHA256_result[206]), .B0(n236), .B1(n145), .Y(
        n2054) );
  AOI22XL U676 ( .A0(n241), .A1(SHA256_result[142]), .B0(n240), .B1(
        SHA256_result[174]), .Y(n2055) );
  AOI221XL U677 ( .A0(n254), .A1(SHA256_result[14]), .B0(n248), .B1(
        SHA256_result[46]), .C0(n2057), .Y(n2056) );
  AOI22XL U678 ( .A0(n238), .A1(SHA256_result[207]), .B0(n236), .B1(n144), .Y(
        n2050) );
  AOI22XL U679 ( .A0(n241), .A1(SHA256_result[143]), .B0(n240), .B1(
        SHA256_result[175]), .Y(n2051) );
  AOI22XL U680 ( .A0(n237), .A1(SHA256_result[208]), .B0(n236), .B1(n143), .Y(
        n2046) );
  AOI22XL U681 ( .A0(n241), .A1(SHA256_result[144]), .B0(n240), .B1(
        SHA256_result[176]), .Y(n2047) );
  AOI221XL U682 ( .A0(n254), .A1(SHA256_result[16]), .B0(n248), .B1(
        SHA256_result[48]), .C0(n2049), .Y(n2048) );
  AOI22XL U683 ( .A0(n238), .A1(SHA256_result[209]), .B0(n236), .B1(n142), .Y(
        n2042) );
  AOI22XL U684 ( .A0(n241), .A1(SHA256_result[145]), .B0(n240), .B1(
        SHA256_result[177]), .Y(n2043) );
  AOI221XL U685 ( .A0(n254), .A1(SHA256_result[17]), .B0(n248), .B1(
        SHA256_result[49]), .C0(n2045), .Y(n2044) );
  AOI22XL U686 ( .A0(n237), .A1(SHA256_result[210]), .B0(n236), .B1(n141), .Y(
        n2038) );
  AOI22XL U687 ( .A0(n241), .A1(SHA256_result[146]), .B0(n240), .B1(
        SHA256_result[178]), .Y(n2039) );
  AOI221XL U688 ( .A0(n254), .A1(SHA256_result[18]), .B0(n249), .B1(
        SHA256_result[50]), .C0(n2041), .Y(n2040) );
  AOI22XL U689 ( .A0(n238), .A1(SHA256_result[211]), .B0(n236), .B1(n140), .Y(
        n2034) );
  AOI221XL U690 ( .A0(n254), .A1(SHA256_result[19]), .B0(n249), .B1(
        SHA256_result[51]), .C0(n2037), .Y(n2036) );
  AOI22XL U691 ( .A0(n237), .A1(SHA256_result[212]), .B0(n236), .B1(n139), .Y(
        n2030) );
  AOI221XL U692 ( .A0(n254), .A1(SHA256_result[20]), .B0(n249), .B1(
        SHA256_result[52]), .C0(n2033), .Y(n2032) );
  AOI22XL U693 ( .A0(n238), .A1(SHA256_result[213]), .B0(n236), .B1(n138), .Y(
        n2026) );
  AOI221XL U694 ( .A0(n254), .A1(SHA256_result[21]), .B0(n249), .B1(
        SHA256_result[53]), .C0(n2029), .Y(n2028) );
  AOI22XL U695 ( .A0(n237), .A1(SHA256_result[214]), .B0(n236), .B1(
        SHA256_result[246]), .Y(n2022) );
  AOI221XL U696 ( .A0(n254), .A1(SHA256_result[22]), .B0(n249), .B1(
        SHA256_result[54]), .C0(n2025), .Y(n2024) );
  AOI22XL U697 ( .A0(n238), .A1(SHA256_result[215]), .B0(n236), .B1(n137), .Y(
        n2018) );
  AOI221XL U698 ( .A0(n254), .A1(SHA256_result[23]), .B0(n249), .B1(
        SHA256_result[55]), .C0(n2021), .Y(n2020) );
  AOI31XL U699 ( .A0(n2226), .A1(n346), .A2(n2138), .B0(n2190), .Y(n2399) );
  NOR3XL U700 ( .A(n2373), .B(n2148), .C(n2190), .Y(n2365) );
  AOI211XL U701 ( .A0(n2302), .A1(n32), .B0(n2339), .C0(n2340), .Y(n2338) );
  AOI22XL U702 ( .A0(n238), .A1(SHA256_result[216]), .B0(n236), .B1(n136), .Y(
        n2014) );
  AOI221XL U703 ( .A0(n254), .A1(SHA256_result[24]), .B0(n249), .B1(
        SHA256_result[56]), .C0(n2017), .Y(n2016) );
  AOI22XL U704 ( .A0(n238), .A1(SHA256_result[217]), .B0(n235), .B1(n135), .Y(
        n2010) );
  AOI211XL U705 ( .A0(n248), .A1(SHA256_result[57]), .B0(n374), .C0(n373), .Y(
        n2012) );
  AOI22XL U706 ( .A0(n238), .A1(SHA256_result[218]), .B0(n236), .B1(n134), .Y(
        n2006) );
  AOI22XL U707 ( .A0(n238), .A1(SHA256_result[219]), .B0(n235), .B1(n133), .Y(
        n2002) );
  AOI22XL U708 ( .A0(n238), .A1(SHA256_result[220]), .B0(n236), .B1(
        SHA256_result[252]), .Y(n1998) );
  AOI22XL U709 ( .A0(n238), .A1(SHA256_result[221]), .B0(n235), .B1(n132), .Y(
        n1994) );
  AOI22XL U710 ( .A0(n238), .A1(SHA256_result[222]), .B0(n236), .B1(n131), .Y(
        n1990) );
  AOI22XL U711 ( .A0(n238), .A1(SHA256_result[223]), .B0(n235), .B1(n25), .Y(
        n1979) );
  AND3X1 U712 ( .A(n1434), .B(n392), .C(inner_busy), .Y(n130) );
  NOR3XL U713 ( .A(n1370), .B(round[2]), .C(n127), .Y(n2323) );
  NOR3XL U714 ( .A(n781), .B(n1383), .C(n345), .Y(n2234) );
  NOR3XL U715 ( .A(n1383), .B(n160), .C(n756), .Y(n2140) );
  INVX1 U716 ( .A(n344), .Y(n343) );
  OAI22XL U717 ( .A0(round[3]), .A1(n2181), .B0(n2395), .B1(n1370), .Y(n2394)
         );
  NOR2XL U718 ( .A(n1383), .B(round[2]), .Y(n116) );
  NOR2XL U719 ( .A(n1388), .B(round[3]), .Y(n2139) );
  NOR2XL U720 ( .A(n1370), .B(round[3]), .Y(n2206) );
  AOI222XL U721 ( .A0(n2350), .A1(n1383), .B0(n2302), .B1(n1370), .C0(n2306), 
        .C1(n160), .Y(n2390) );
  OAI22XL U722 ( .A0(n888), .A1(n1984), .B0(n1156), .B1(n244), .Y(n2065) );
  OAI22XL U723 ( .A0(n890), .A1(n1984), .B0(n1154), .B1(n244), .Y(n2057) );
  OAI22XL U724 ( .A0(n891), .A1(n1984), .B0(n1153), .B1(n244), .Y(n2053) );
  OAI22XL U725 ( .A0(n893), .A1(n1984), .B0(n1151), .B1(n244), .Y(n2045) );
  OAI22XL U726 ( .A0(n1163), .A1(n244), .B0(n246), .B1(n84), .Y(n360) );
  OAI22XL U727 ( .A0(n1161), .A1(n244), .B0(n246), .B1(n520), .Y(n364) );
  OAI22XL U728 ( .A0(n1160), .A1(n244), .B0(n246), .B1(n515), .Y(n366) );
  OAI22XL U729 ( .A0(n1157), .A1(n244), .B0(n246), .B1(n502), .Y(n372) );
  OAI22XL U730 ( .A0(n892), .A1(n1984), .B0(n1152), .B1(n244), .Y(n2049) );
  OAI22XL U731 ( .A0(n1165), .A1(n244), .B0(n246), .B1(n535), .Y(n356) );
  OAI22XL U732 ( .A0(n1985), .A1(n1168), .B0(n246), .B1(n70), .Y(n350) );
  OAI22XL U733 ( .A0(n1167), .A1(n1985), .B0(n246), .B1(n542), .Y(n352) );
  OAI22XL U734 ( .A0(n899), .A1(n246), .B0(n1145), .B1(n1985), .Y(n2021) );
  AND2X1 U735 ( .A(n255), .B(SHA256_result[0]), .Y(n349) );
  AND2X1 U736 ( .A(n255), .B(SHA256_result[5]), .Y(n359) );
  AND2X1 U737 ( .A(n255), .B(SHA256_result[6]), .Y(n361) );
  AND2X1 U738 ( .A(n255), .B(SHA256_result[7]), .Y(n363) );
  AND2X1 U739 ( .A(n255), .B(SHA256_result[8]), .Y(n365) );
  AND2X1 U740 ( .A(n255), .B(SHA256_result[9]), .Y(n367) );
  AND2X1 U741 ( .A(n255), .B(SHA256_result[10]), .Y(n369) );
  AND2X1 U742 ( .A(n255), .B(SHA256_result[11]), .Y(n371) );
  INVXL U743 ( .A(SHA256_result[127]), .Y(n550) );
  INVXL U744 ( .A(SHA256_result[252]), .Y(n740) );
  INVXL U745 ( .A(SHA256_result[119]), .Y(n899) );
  INVXL U746 ( .A(SHA256_result[118]), .Y(n898) );
  INVXL U747 ( .A(SHA256_result[120]), .Y(n900) );
  INVXL U748 ( .A(SHA256_result[114]), .Y(n894) );
  INVXL U749 ( .A(SHA256_result[121]), .Y(n468) );
  INVXL U750 ( .A(SHA256_result[112]), .Y(n892) );
  INVXL U751 ( .A(n51), .Y(n452) );
  INVXL U752 ( .A(SHA256_result[115]), .Y(n895) );
  INVXL U753 ( .A(SHA256_result[126]), .Y(n440) );
  INVXL U754 ( .A(SHA256_result[116]), .Y(n896) );
  INVXL U755 ( .A(SHA256_result[117]), .Y(n897) );
  INVXL U756 ( .A(SHA256_result[113]), .Y(n893) );
  AND2X1 U757 ( .A(n254), .B(SHA256_result[4]), .Y(n357) );
  AND2X1 U758 ( .A(n254), .B(SHA256_result[2]), .Y(n353) );
  AND2X1 U759 ( .A(n254), .B(SHA256_result[1]), .Y(n351) );
  AND2X1 U760 ( .A(n254), .B(SHA256_result[3]), .Y(n355) );
  INVXL U761 ( .A(SHA256_result[246]), .Y(n646) );
  INVXL U762 ( .A(SHA256_result[82]), .Y(n906) );
  INVXL U763 ( .A(SHA256_result[77]), .Y(n905) );
  INVXL U764 ( .A(SHA256_result[70]), .Y(n902) );
  INVXL U765 ( .A(SHA256_result[73]), .Y(n903) );
  INVXL U766 ( .A(SHA256_result[74]), .Y(n904) );
  INVXL U767 ( .A(SHA256_result[86]), .Y(n910) );
  INVXL U768 ( .A(SHA256_result[85]), .Y(n909) );
  INVXL U769 ( .A(SHA256_result[84]), .Y(n908) );
  INVXL U770 ( .A(SHA256_result[83]), .Y(n907) );
  INVXL U771 ( .A(SHA256_result[210]), .Y(n815) );
  INVXL U772 ( .A(SHA256_result[209]), .Y(n814) );
  INVXL U773 ( .A(SHA256_result[207]), .Y(n812) );
  INVXL U774 ( .A(SHA256_result[205]), .Y(n810) );
  INVXL U775 ( .A(SHA256_result[201]), .Y(n806) );
  INVXL U776 ( .A(SHA256_result[206]), .Y(n811) );
  INVXL U777 ( .A(SHA256_result[204]), .Y(n809) );
  INVXL U778 ( .A(SHA256_result[200]), .Y(n805) );
  INVXL U779 ( .A(SHA256_result[198]), .Y(n803) );
  INVXL U780 ( .A(SHA256_result[197]), .Y(n802) );
  INVXL U781 ( .A(SHA256_result[196]), .Y(n801) );
  INVXL U782 ( .A(SHA256_result[178]), .Y(n842) );
  INVXL U783 ( .A(SHA256_result[177]), .Y(n841) );
  INVXL U784 ( .A(SHA256_result[175]), .Y(n839) );
  INVXL U785 ( .A(SHA256_result[174]), .Y(n838) );
  INVXL U786 ( .A(SHA256_result[173]), .Y(n837) );
  INVXL U787 ( .A(SHA256_result[172]), .Y(n836) );
  INVXL U788 ( .A(SHA256_result[168]), .Y(n832) );
  INVXL U789 ( .A(SHA256_result[165]), .Y(n829) );
  INVXL U790 ( .A(SHA256_result[164]), .Y(n828) );
  INVXL U791 ( .A(SHA256_result[42]), .Y(n917) );
  INVXL U792 ( .A(SHA256_result[54]), .Y(n929) );
  INVXL U793 ( .A(SHA256_result[53]), .Y(n928) );
  INVXL U794 ( .A(SHA256_result[176]), .Y(n840) );
  INVXL U795 ( .A(SHA256_result[170]), .Y(n834) );
  INVXL U796 ( .A(SHA256_result[123]), .Y(n460) );
  INVXL U797 ( .A(SHA256_result[122]), .Y(n464) );
  INVXL U798 ( .A(SHA256_result[107]), .Y(n502) );
  INVXL U799 ( .A(SHA256_result[208]), .Y(n813) );
  INVXL U800 ( .A(SHA256_result[203]), .Y(n808) );
  INVXL U801 ( .A(SHA256_result[202]), .Y(n807) );
  INVXL U802 ( .A(SHA256_result[199]), .Y(n804) );
  INVXL U803 ( .A(SHA256_result[194]), .Y(n799) );
  INVXL U804 ( .A(SHA256_result[195]), .Y(n800) );
  INVXL U805 ( .A(SHA256_result[41]), .Y(n916) );
  INVXL U806 ( .A(n50), .Y(n913) );
  INVXL U807 ( .A(SHA256_result[169]), .Y(n833) );
  INVXL U808 ( .A(SHA256_result[166]), .Y(n830) );
  INVXL U809 ( .A(SHA256_result[52]), .Y(n927) );
  INVXL U810 ( .A(SHA256_result[51]), .Y(n926) );
  INVXL U811 ( .A(SHA256_result[50]), .Y(n925) );
  INVXL U812 ( .A(SHA256_result[45]), .Y(n920) );
  INVXL U813 ( .A(SHA256_result[171]), .Y(n835) );
  INVXL U814 ( .A(SHA256_result[167]), .Y(n831) );
  INVXL U815 ( .A(SHA256_result[2]), .Y(n942) );
  NOR2XL U816 ( .A(n161), .B(n1383), .Y(n2334) );
  INVXL U817 ( .A(SHA256_result[129]), .Y(n858) );
  INVXL U818 ( .A(SHA256_result[161]), .Y(n565) );
  INVXL U819 ( .A(SHA256_result[1]), .Y(n941) );
  INVXL U820 ( .A(SHA256_result[10]), .Y(n950) );
  INVXL U821 ( .A(SHA256_result[21]), .Y(n961) );
  INVXL U822 ( .A(SHA256_result[15]), .Y(n955) );
  INVXL U823 ( .A(SHA256_result[14]), .Y(n954) );
  INVXL U824 ( .A(SHA256_result[11]), .Y(n951) );
  INVXL U825 ( .A(SHA256_result[8]), .Y(n948) );
  INVXL U826 ( .A(SHA256_result[6]), .Y(n946) );
  INVXL U827 ( .A(SHA256_result[20]), .Y(n960) );
  INVXL U828 ( .A(SHA256_result[17]), .Y(n957) );
  INVXL U829 ( .A(SHA256_result[16]), .Y(n956) );
  INVXL U830 ( .A(SHA256_result[13]), .Y(n953) );
  INVXL U831 ( .A(SHA256_result[12]), .Y(n952) );
  INVXL U832 ( .A(SHA256_result[19]), .Y(n959) );
  INVXL U833 ( .A(SHA256_result[18]), .Y(n958) );
  INVXL U834 ( .A(SHA256_result[9]), .Y(n949) );
  INVXL U835 ( .A(SHA256_result[128]), .Y(n857) );
  INVXL U836 ( .A(SHA256_result[7]), .Y(n947) );
  INVXL U837 ( .A(SHA256_result[5]), .Y(n945) );
  INVXL U838 ( .A(SHA256_result[124]), .Y(n455) );
  INVXL U839 ( .A(SHA256_result[0]), .Y(n940) );
  INVXL U840 ( .A(SHA256_result[111]), .Y(n891) );
  INVXL U841 ( .A(SHA256_result[3]), .Y(n943) );
  INVXL U842 ( .A(SHA256_result[4]), .Y(n944) );
  INVXL U843 ( .A(SHA256_result[163]), .Y(n558) );
  INVXL U844 ( .A(SHA256_result[106]), .Y(n506) );
  MXI2XL U845 ( .A(n932), .B(n1143), .S0(SHA256_result[121]), .Y(f1_EFG_32[25]) );
  NAND2X1 U846 ( .A(SHA256_result[95]), .B(n274), .Y(n119) );
  OR2X2 U847 ( .A(n162), .B(n938), .Y(n117) );
  OR2X2 U848 ( .A(n314), .B(n743), .Y(n120) );
  OR2XL U849 ( .A(n176), .B(n798), .Y(n121) );
  INVXL U850 ( .A(n25), .Y(n743) );
  OR2X2 U851 ( .A(n301), .B(n855), .Y(n123) );
  OR2XL U852 ( .A(n178), .B(n856), .Y(n124) );
  AOI22XL U853 ( .A0(n1986), .A1(SHA256_result[129]), .B0(n239), .B1(
        SHA256_result[161]), .Y(n2107) );
  INVX1 U854 ( .A(n281), .Y(n269) );
  INVX1 U855 ( .A(n281), .Y(n273) );
  INVX1 U856 ( .A(n279), .Y(n275) );
  INVX1 U857 ( .A(n277), .Y(n276) );
  INVX1 U858 ( .A(n337), .Y(n283) );
  INVX1 U859 ( .A(n337), .Y(n284) );
  INVX1 U860 ( .A(n336), .Y(n285) );
  INVX1 U861 ( .A(n335), .Y(n290) );
  INVX1 U862 ( .A(n335), .Y(n289) );
  INVX1 U863 ( .A(n337), .Y(n282) );
  INVX1 U864 ( .A(n335), .Y(n288) );
  INVX1 U865 ( .A(n336), .Y(n287) );
  INVX1 U866 ( .A(n334), .Y(n292) );
  INVX1 U867 ( .A(n336), .Y(n286) );
  INVX1 U868 ( .A(n334), .Y(n291) );
  INVX1 U869 ( .A(n334), .Y(n293) );
  INVX1 U870 ( .A(n329), .Y(n310) );
  INVX1 U871 ( .A(n329), .Y(n309) );
  INVX1 U872 ( .A(n329), .Y(n308) );
  INVX1 U873 ( .A(n326), .Y(n307) );
  INVX1 U874 ( .A(n332), .Y(n306) );
  INVX1 U875 ( .A(n333), .Y(n305) );
  INVX1 U876 ( .A(n330), .Y(n304) );
  INVX1 U877 ( .A(n330), .Y(n303) );
  INVX1 U878 ( .A(n331), .Y(n302) );
  INVX1 U879 ( .A(n333), .Y(n295) );
  INVX1 U880 ( .A(n332), .Y(n297) );
  INVX1 U881 ( .A(n331), .Y(n300) );
  INVX1 U882 ( .A(n333), .Y(n294) );
  INVX1 U883 ( .A(n333), .Y(n296) );
  INVX1 U884 ( .A(n332), .Y(n299) );
  INVX1 U885 ( .A(n332), .Y(n298) );
  INVX1 U886 ( .A(n331), .Y(n301) );
  INVX1 U887 ( .A(n328), .Y(n312) );
  INVX1 U888 ( .A(n328), .Y(n313) );
  INVX1 U889 ( .A(n327), .Y(n315) );
  INVX1 U890 ( .A(n327), .Y(n316) );
  INVX1 U891 ( .A(n326), .Y(n317) );
  INVX1 U892 ( .A(n326), .Y(n318) );
  INVX1 U893 ( .A(n327), .Y(n314) );
  INVX1 U894 ( .A(n326), .Y(n319) );
  INVX1 U895 ( .A(n338), .Y(n281) );
  INVX1 U896 ( .A(n338), .Y(n280) );
  INVX1 U897 ( .A(n339), .Y(n278) );
  INVX1 U898 ( .A(n338), .Y(n279) );
  INVX1 U899 ( .A(n327), .Y(n321) );
  INVX1 U900 ( .A(n328), .Y(n320) );
  INVX1 U901 ( .A(n327), .Y(n322) );
  INVX1 U902 ( .A(n328), .Y(n324) );
  INVX1 U903 ( .A(n327), .Y(n323) );
  INVX1 U904 ( .A(n328), .Y(n325) );
  INVX1 U905 ( .A(n186), .Y(n177) );
  INVX1 U906 ( .A(n230), .Y(n223) );
  INVX1 U907 ( .A(n232), .Y(n215) );
  INVX1 U908 ( .A(n231), .Y(n216) );
  INVX1 U909 ( .A(n229), .Y(n220) );
  INVX1 U910 ( .A(n230), .Y(n219) );
  INVX1 U911 ( .A(n230), .Y(n218) );
  INVX1 U912 ( .A(n232), .Y(n214) );
  INVX1 U913 ( .A(n232), .Y(n213) );
  INVX1 U914 ( .A(n229), .Y(n221) );
  INVX1 U915 ( .A(n229), .Y(n222) );
  INVX1 U916 ( .A(n231), .Y(n212) );
  INVX1 U917 ( .A(n231), .Y(n217) );
  INVX1 U918 ( .A(n185), .Y(n175) );
  INVX1 U919 ( .A(n266), .Y(n339) );
  INVX1 U920 ( .A(n264), .Y(n329) );
  INVX1 U921 ( .A(n264), .Y(n330) );
  INVX1 U922 ( .A(n264), .Y(n333) );
  INVX1 U923 ( .A(n264), .Y(n332) );
  INVX1 U924 ( .A(n264), .Y(n331) );
  INVX1 U925 ( .A(n263), .Y(n328) );
  INVX1 U926 ( .A(n263), .Y(n327) );
  INVX1 U927 ( .A(n265), .Y(n337) );
  INVX1 U928 ( .A(n264), .Y(n326) );
  INVX1 U929 ( .A(n265), .Y(n335) );
  INVX1 U930 ( .A(n265), .Y(n336) );
  INVX1 U931 ( .A(n265), .Y(n334) );
  INVX1 U932 ( .A(n211), .Y(n227) );
  INVX1 U933 ( .A(n211), .Y(n226) );
  INVX1 U934 ( .A(n211), .Y(n225) );
  INVX1 U935 ( .A(n193), .Y(n179) );
  INVX1 U936 ( .A(n193), .Y(n180) );
  INVX1 U937 ( .A(n192), .Y(n181) );
  INVX1 U938 ( .A(n189), .Y(n184) );
  INVX1 U939 ( .A(n191), .Y(n182) );
  INVX1 U940 ( .A(n190), .Y(n183) );
  INVX1 U941 ( .A(n210), .Y(n230) );
  INVX1 U942 ( .A(n210), .Y(n232) );
  INVX1 U943 ( .A(n210), .Y(n229) );
  INVX1 U944 ( .A(n210), .Y(n231) );
  INVX1 U945 ( .A(n207), .Y(n206) );
  INVX1 U946 ( .A(n722), .Y(n228) );
  INVX1 U947 ( .A(n172), .Y(n164) );
  INVX1 U948 ( .A(n172), .Y(n163) );
  INVX1 U949 ( .A(n677), .Y(n258) );
  INVX1 U950 ( .A(n677), .Y(n260) );
  INVX1 U951 ( .A(n677), .Y(n261) );
  INVX1 U952 ( .A(n677), .Y(n256) );
  INVX1 U953 ( .A(n677), .Y(n262) );
  INVX1 U954 ( .A(n173), .Y(n167) );
  INVX1 U955 ( .A(n721), .Y(n209) );
  INVX1 U956 ( .A(n721), .Y(n208) );
  INVX1 U957 ( .A(n267), .Y(n266) );
  INVX1 U958 ( .A(n268), .Y(n264) );
  INVX1 U959 ( .A(n268), .Y(n263) );
  INVX1 U960 ( .A(n267), .Y(n265) );
  INVX1 U961 ( .A(n715), .Y(n189) );
  INVX1 U962 ( .A(n715), .Y(n193) );
  INVX1 U963 ( .A(n715), .Y(n188) );
  INVX1 U964 ( .A(n715), .Y(n190) );
  INVX1 U965 ( .A(n715), .Y(n192) );
  INVX1 U966 ( .A(n715), .Y(n191) );
  INVX1 U967 ( .A(n715), .Y(n194) );
  INVX1 U968 ( .A(n2259), .Y(n749) );
  INVX1 U969 ( .A(n2325), .Y(n790) );
  INVX1 U970 ( .A(n2209), .Y(n785) );
  INVX1 U971 ( .A(n2277), .Y(n768) );
  NOR2X1 U972 ( .A(n769), .B(n788), .Y(n2190) );
  INVX1 U973 ( .A(n2249), .Y(n778) );
  NOR2X1 U974 ( .A(n795), .B(n791), .Y(n2162) );
  INVX1 U975 ( .A(n2134), .Y(n795) );
  INVX1 U976 ( .A(n2283), .Y(n755) );
  NAND4X1 U977 ( .A(n790), .B(n755), .C(n2199), .D(n766), .Y(n2242) );
  NAND2X1 U978 ( .A(n2266), .B(n127), .Y(n2200) );
  INVX1 U979 ( .A(n2276), .Y(n774) );
  AOI21X1 U980 ( .A0(n791), .A1(n758), .B0(n797), .Y(n2362) );
  INVX1 U981 ( .A(n2396), .Y(n747) );
  INVX1 U982 ( .A(n2224), .Y(n771) );
  NAND2X1 U983 ( .A(n764), .B(n756), .Y(n2251) );
  INVX1 U984 ( .A(n2306), .Y(n752) );
  INVX1 U985 ( .A(n2175), .Y(n746) );
  NAND2X1 U986 ( .A(n772), .B(n768), .Y(n2238) );
  NAND2X1 U987 ( .A(n765), .B(n795), .Y(n2275) );
  INVX1 U988 ( .A(n36), .Y(n236) );
  NOR2X1 U989 ( .A(n166), .B(n642), .Y(n643) );
  OAI2BB1X1 U990 ( .A0N(N821), .A1N(n195), .B0(n632), .Y(n2869) );
  NOR2X1 U991 ( .A(n166), .B(n630), .Y(n631) );
  OAI2BB1X1 U992 ( .A0N(N819), .A1N(n197), .B0(n640), .Y(n2871) );
  AOI21XL U993 ( .A0(next_A[24]), .A1(n275), .B0(n639), .Y(n640) );
  NAND2BX1 U994 ( .AN(n393), .B(n1491), .Y(n1490) );
  INVX1 U995 ( .A(n174), .Y(n169) );
  INVX1 U996 ( .A(n174), .Y(n170) );
  INVX1 U997 ( .A(n174), .Y(n171) );
  INVX1 U998 ( .A(n716), .Y(n717) );
  INVX1 U999 ( .A(n174), .Y(n168) );
  INVX1 U1000 ( .A(n2378), .Y(n797) );
  INVX1 U1001 ( .A(n2148), .Y(n792) );
  NAND3X1 U1002 ( .A(n345), .B(n32), .C(n1878), .Y(n1859) );
  AOI31X1 U1003 ( .A0(n2298), .A1(n2299), .A2(n2300), .B0(n233), .Y(N2961) );
  NOR3X1 U1004 ( .A(n2303), .B(n2219), .C(n2293), .Y(n2299) );
  AOI211X1 U1005 ( .A0(n2249), .A1(n1396), .B0(n2301), .C0(n2282), .Y(n2300)
         );
  AOI31X1 U1006 ( .A0(n763), .A1(n787), .A2(n2114), .B0(n233), .Y(N2977) );
  INVX1 U1007 ( .A(n2116), .Y(n787) );
  INVX1 U1008 ( .A(n2117), .Y(n763) );
  AND4X2 U1009 ( .A(n789), .B(n759), .C(n778), .D(n779), .Y(n2114) );
  INVX1 U1010 ( .A(n253), .Y(n251) );
  INVX1 U1011 ( .A(n253), .Y(n252) );
  NOR2X1 U1012 ( .A(n788), .B(n794), .Y(n2209) );
  NOR2X1 U1013 ( .A(n796), .B(n791), .Y(n2325) );
  NOR2X1 U1014 ( .A(n750), .B(n346), .Y(n2259) );
  NOR2X1 U1015 ( .A(n769), .B(n794), .Y(n2277) );
  OAI21XL U1016 ( .A0(n347), .A1(n749), .B0(n2372), .Y(n2386) );
  NAND4X1 U1017 ( .A(n2263), .B(n745), .C(n778), .D(n759), .Y(n2320) );
  INVX1 U1018 ( .A(n2322), .Y(n759) );
  NAND3BX1 U1019 ( .AN(n2174), .B(n749), .C(n745), .Y(n2170) );
  INVX1 U1020 ( .A(n2342), .Y(n750) );
  AOI21X1 U1021 ( .A0(n749), .A1(n2146), .B0(n345), .Y(n2236) );
  INVX1 U1022 ( .A(n2135), .Y(n756) );
  NOR2X1 U1023 ( .A(n783), .B(n756), .Y(n2283) );
  NOR2X1 U1024 ( .A(n786), .B(n769), .Y(n2177) );
  INVX1 U1025 ( .A(n2305), .Y(n788) );
  NOR2X1 U1026 ( .A(n796), .B(n781), .Y(n2174) );
  NOR2X1 U1027 ( .A(n781), .B(n794), .Y(n2249) );
  OAI222XL U1028 ( .A0(n781), .A1(n764), .B0(n796), .B1(n746), .C0(round[1]), 
        .C1(n2165), .Y(n2301) );
  NOR3X1 U1029 ( .A(n345), .B(n791), .C(n793), .Y(n2151) );
  NAND2X1 U1030 ( .A(n2398), .B(n347), .Y(n2166) );
  INVX1 U1031 ( .A(n2220), .Y(n764) );
  NOR2X1 U1032 ( .A(n127), .B(n346), .Y(n2175) );
  NOR2X1 U1033 ( .A(n788), .B(n347), .Y(n2350) );
  NOR2X1 U1034 ( .A(n793), .B(n756), .Y(n2183) );
  OAI22X1 U1035 ( .A0(n347), .A1(n796), .B0(n769), .B1(n793), .Y(n2356) );
  NOR2X1 U1036 ( .A(n765), .B(n794), .Y(n2247) );
  NOR2X1 U1037 ( .A(n2333), .B(n347), .Y(n2224) );
  NOR2X1 U1038 ( .A(n769), .B(n796), .Y(n2219) );
  NOR2X1 U1039 ( .A(n793), .B(n777), .Y(n2266) );
  NAND2X1 U1040 ( .A(n2249), .B(n347), .Y(n2199) );
  INVX1 U1041 ( .A(n2312), .Y(n789) );
  NOR2X1 U1042 ( .A(n777), .B(n794), .Y(n2161) );
  INVX1 U1043 ( .A(n114), .Y(n791) );
  INVX1 U1044 ( .A(n2372), .Y(n782) );
  NOR2X1 U1045 ( .A(n756), .B(n794), .Y(n2306) );
  NOR4BBX1 U1046 ( .AN(n2159), .BN(n2263), .C(n2225), .D(n2283), .Y(n2413) );
  AOI31X1 U1047 ( .A0(n773), .A1(n792), .A2(n2132), .B0(round[1]), .Y(n2131)
         );
  INVX1 U1048 ( .A(n2314), .Y(n772) );
  OAI22X1 U1049 ( .A0(n346), .A1(n2149), .B0(n796), .B1(n751), .Y(n2346) );
  INVX1 U1050 ( .A(n1878), .Y(n770) );
  INVX1 U1051 ( .A(n2252), .Y(n758) );
  NOR2X1 U1052 ( .A(n777), .B(n797), .Y(n2276) );
  NAND3X1 U1053 ( .A(n770), .B(n771), .C(n753), .Y(n2360) );
  INVX1 U1054 ( .A(n2248), .Y(n757) );
  NOR2X1 U1055 ( .A(n796), .B(n345), .Y(n2134) );
  AOI21X1 U1056 ( .A0(n2159), .A1(n774), .B0(n347), .Y(n2292) );
  INVX1 U1057 ( .A(n2294), .Y(n766) );
  INVX1 U1058 ( .A(n2258), .Y(n751) );
  NAND2X1 U1059 ( .A(n2195), .B(n2138), .Y(n2210) );
  NAND3X1 U1060 ( .A(n2199), .B(n766), .C(n2263), .Y(n2291) );
  NAND3X1 U1061 ( .A(n2184), .B(n753), .C(n752), .Y(n2376) );
  NAND3X1 U1062 ( .A(n2184), .B(n779), .C(n2132), .Y(n2182) );
  AOI21X1 U1063 ( .A0(n778), .A1(n790), .B0(n347), .Y(n2348) );
  AOI21X1 U1064 ( .A0(n2156), .A1(n790), .B0(n1396), .Y(n2197) );
  NAND2X1 U1065 ( .A(n347), .B(n1878), .Y(n2233) );
  NAND3X1 U1066 ( .A(n771), .B(n779), .C(n2233), .Y(n2230) );
  AOI21X1 U1067 ( .A0(n745), .A1(n770), .B0(n346), .Y(n2296) );
  OAI21XL U1068 ( .A0(n112), .A1(n777), .B0(n757), .Y(n2235) );
  OAI2BB1X1 U1069 ( .A0N(n113), .A1N(n2137), .B0(n2333), .Y(n2380) );
  NAND3X1 U1070 ( .A(n2184), .B(n2159), .C(n2149), .Y(n2207) );
  INVX1 U1071 ( .A(n2189), .Y(n776) );
  NAND2X1 U1072 ( .A(n2342), .B(n2305), .Y(n2160) );
  OAI2BB1X1 U1073 ( .A0N(n1393), .A1N(n2266), .B0(n753), .Y(n2321) );
  INVX1 U1074 ( .A(n245), .Y(n244) );
  INVX1 U1075 ( .A(n112), .Y(n765) );
  OAI222XL U1076 ( .A0(n788), .A1(n754), .B0(n756), .B1(n2146), .C0(n792), 
        .C1(n1396), .Y(n2273) );
  INVX1 U1077 ( .A(n2221), .Y(n754) );
  NOR2X1 U1078 ( .A(n346), .B(n797), .Y(n2304) );
  NOR3X1 U1079 ( .A(n781), .B(n797), .C(n345), .Y(n2152) );
  NAND2X1 U1080 ( .A(n2135), .B(n114), .Y(n2181) );
  INVX1 U1081 ( .A(n2223), .Y(n761) );
  NAND2X1 U1082 ( .A(n777), .B(n791), .Y(n2122) );
  INVX1 U1083 ( .A(n2187), .Y(n760) );
  INVX1 U1084 ( .A(n243), .Y(n241) );
  INVX1 U1085 ( .A(n36), .Y(n235) );
  INVX1 U1086 ( .A(n33), .Y(n240) );
  INVX1 U1087 ( .A(n250), .Y(n248) );
  INVX1 U1088 ( .A(n34), .Y(n255) );
  INVX1 U1089 ( .A(n35), .Y(n238) );
  INVX1 U1090 ( .A(n243), .Y(n242) );
  INVX1 U1091 ( .A(n250), .Y(n249) );
  AOI31X1 U1092 ( .A0(n387), .A1(n390), .A2(n388), .B0(n1849), .Y(n722) );
  OAI221XL U1093 ( .A0(n295), .A1(n935), .B0(n1457), .B1(n968), .C0(n1461), 
        .Y(n2451) );
  AOI21X1 U1094 ( .A0(N1047), .A1(n195), .B0(n257), .Y(n1461) );
  OAI221XL U1095 ( .A0(n315), .A1(n741), .B0(n176), .B1(n826), .C0(n1757), .Y(
        n2802) );
  AOI21X1 U1096 ( .A0(N856), .A1(n203), .B0(n258), .Y(n1757) );
  OAI221XL U1097 ( .A0(n315), .A1(n740), .B0(n176), .B1(n825), .C0(n1758), .Y(
        n2803) );
  AOI21X1 U1098 ( .A0(N855), .A1(n198), .B0(n259), .Y(n1758) );
  OAI221XL U1099 ( .A0(n294), .A1(n826), .B0(n177), .B1(n853), .C0(n1725), .Y(
        n2769) );
  AOI21X1 U1100 ( .A0(N888), .A1(n203), .B0(n261), .Y(n1725) );
  OAI221XL U1101 ( .A0(n296), .A1(n825), .B0(n177), .B1(n852), .C0(n1726), .Y(
        n2770) );
  AOI21X1 U1102 ( .A0(N887), .A1(n196), .B0(n261), .Y(n1726) );
  OAI221XL U1103 ( .A0(n299), .A1(n853), .B0(n178), .B1(n886), .C0(n1693), .Y(
        n2737) );
  OAI211X1 U1104 ( .A0(n655), .A1(n320), .B0(n654), .C0(n653), .Y(n2876) );
  OAI211X1 U1105 ( .A0(n287), .A1(n662), .B0(n661), .C0(n660), .Y(n2879) );
  INVXL U1106 ( .A(next_A[16]), .Y(n662) );
  NAND2X1 U1107 ( .A(N811), .B(n200), .Y(n660) );
  OAI211X1 U1108 ( .A0(n292), .A1(n665), .B0(n664), .C0(n663), .Y(n2880) );
  INVXL U1109 ( .A(next_A[15]), .Y(n665) );
  OAI211X1 U1110 ( .A0(n289), .A1(n668), .B0(n667), .C0(n666), .Y(n2881) );
  INVXL U1111 ( .A(next_A[14]), .Y(n668) );
  XOR3X2 U1112 ( .A(n154), .B(n143), .C(n135), .Y(f3_A_32[3]) );
  AOI22X1 U1113 ( .A0(N857), .A1(n202), .B0(n131), .B1(n270), .Y(n1756) );
  NAND2XL U1114 ( .A(next_A[30]), .B(n276), .Y(n619) );
  NOR2X1 U1115 ( .A(n899), .B(n167), .Y(n474) );
  OAI2BB1X1 U1116 ( .A0N(N945), .A1N(n199), .B0(n477), .Y(n2712) );
  NOR2X1 U1117 ( .A(n898), .B(n167), .Y(n476) );
  AOI21XL U1118 ( .A0(next_A[22]), .A1(n275), .B0(n647), .Y(n648) );
  NOR2X1 U1119 ( .A(n166), .B(n646), .Y(n647) );
  NOR2X1 U1120 ( .A(n167), .B(n464), .Y(n465) );
  OAI2BB1X1 U1121 ( .A0N(N816), .A1N(n204), .B0(n650), .Y(n2874) );
  AOI2BB2X1 U1122 ( .B0(n168), .B1(n138), .A0N(n320), .A1N(n649), .Y(n650) );
  INVXL U1123 ( .A(next_A[21]), .Y(n649) );
  AOI21XL U1124 ( .A0(next_A[28]), .A1(n275), .B0(n624), .Y(n625) );
  NOR2X1 U1125 ( .A(n740), .B(n167), .Y(n624) );
  AOI21XL U1126 ( .A0(next_E[27]), .A1(n276), .B0(n461), .Y(n462) );
  NOR2X1 U1127 ( .A(n167), .B(n460), .Y(n461) );
  NOR2X1 U1128 ( .A(n166), .B(n550), .Y(n551) );
  NOR2X1 U1129 ( .A(n743), .B(n167), .Y(n616) );
  OAI2BB1X1 U1130 ( .A0N(N815), .A1N(n203), .B0(n652), .Y(n2875) );
  AOI2BB2X1 U1131 ( .B0(n168), .B1(n139), .A0N(n322), .A1N(n651), .Y(n652) );
  OAI2BB1X1 U1132 ( .A0N(N812), .A1N(n200), .B0(n659), .Y(n2878) );
  AOI2BB2X1 U1133 ( .B0(n168), .B1(n142), .A0N(n278), .A1N(n658), .Y(n659) );
  INVXL U1134 ( .A(next_A[17]), .Y(n658) );
  OAI2BB1X1 U1135 ( .A0N(N813), .A1N(n721), .B0(n657), .Y(n2877) );
  AOI2BB2X1 U1136 ( .B0(n169), .B1(n141), .A0N(n280), .A1N(n656), .Y(n657) );
  OAI221XL U1137 ( .A0(n319), .A1(n685), .B0(n48), .B1(n684), .C0(n683), .Y(
        n2887) );
  INVX1 U1138 ( .A(next_A[8]), .Y(n685) );
  INVX1 U1139 ( .A(N803), .Y(n684) );
  NAND2X1 U1140 ( .A(n169), .B(n151), .Y(n683) );
  OAI221XL U1141 ( .A0(n319), .A1(n688), .B0(n48), .B1(n687), .C0(n686), .Y(
        n2888) );
  INVX1 U1142 ( .A(N802), .Y(n687) );
  NAND2X1 U1143 ( .A(n169), .B(n152), .Y(n686) );
  OAI221XL U1144 ( .A0(n310), .A1(n934), .B0(n1457), .B1(n967), .C0(n1462), 
        .Y(n2452) );
  AOI21X1 U1145 ( .A0(N1046), .A1(n202), .B0(n257), .Y(n1462) );
  OAI221XL U1146 ( .A0(n310), .A1(n932), .B0(n1457), .B1(n965), .C0(n1464), 
        .Y(n2454) );
  AOI21X1 U1147 ( .A0(N1044), .A1(n195), .B0(n257), .Y(n1464) );
  OAI221XL U1148 ( .A0(n310), .A1(n931), .B0(n1457), .B1(n964), .C0(n1465), 
        .Y(n2455) );
  AOI21X1 U1149 ( .A0(N1043), .A1(n201), .B0(n257), .Y(n1465) );
  OAI221XL U1150 ( .A0(n309), .A1(n930), .B0(n1457), .B1(n963), .C0(n1466), 
        .Y(n2456) );
  AOI21X1 U1151 ( .A0(N1042), .A1(n199), .B0(n257), .Y(n1466) );
  OAI221XL U1152 ( .A0(n309), .A1(n929), .B0(n1457), .B1(n962), .C0(n1467), 
        .Y(n2457) );
  AOI21X1 U1153 ( .A0(N1041), .A1(n206), .B0(n257), .Y(n1467) );
  OAI221XL U1154 ( .A0(n309), .A1(n928), .B0(n1457), .B1(n961), .C0(n1468), 
        .Y(n2458) );
  OAI221XL U1155 ( .A0(n308), .A1(n922), .B0(n1457), .B1(n955), .C0(n1474), 
        .Y(n2464) );
  AOI21X1 U1156 ( .A0(N1034), .A1(n195), .B0(n257), .Y(n1474) );
  OAI221XL U1157 ( .A0(n308), .A1(n921), .B0(n1457), .B1(n954), .C0(n1475), 
        .Y(n2465) );
  AOI21X1 U1158 ( .A0(N1033), .A1(n201), .B0(n257), .Y(n1475) );
  OAI221XL U1159 ( .A0(n308), .A1(n918), .B0(n1457), .B1(n951), .C0(n1478), 
        .Y(n2468) );
  OAI221XL U1160 ( .A0(n307), .A1(n917), .B0(n1457), .B1(n950), .C0(n1479), 
        .Y(n2469) );
  AOI21X1 U1161 ( .A0(N1029), .A1(n204), .B0(n258), .Y(n1479) );
  OAI221XL U1162 ( .A0(n307), .A1(n915), .B0(n1457), .B1(n948), .C0(n1481), 
        .Y(n2471) );
  OAI221XL U1163 ( .A0(n303), .A1(n894), .B0(n176), .B1(n906), .C0(n1623), .Y(
        n2684) );
  OAI221XL U1164 ( .A0(n302), .A1(n889), .B0(n178), .B1(n905), .C0(n1628), .Y(
        n2689) );
  OAI221XL U1165 ( .A0(n315), .A1(n739), .B0(n176), .B1(n824), .C0(n1759), .Y(
        n2804) );
  AOI21X1 U1166 ( .A0(N854), .A1(n717), .B0(n256), .Y(n1759) );
  OAI221XL U1167 ( .A0(n316), .A1(n738), .B0(n176), .B1(n818), .C0(n1765), .Y(
        n2810) );
  AOI21X1 U1168 ( .A0(N848), .A1(n204), .B0(n262), .Y(n1765) );
  OAI221XL U1169 ( .A0(n316), .A1(n735), .B0(n176), .B1(n815), .C0(n1768), .Y(
        n2813) );
  OAI221XL U1170 ( .A0(n316), .A1(n734), .B0(n176), .B1(n814), .C0(n1769), .Y(
        n2814) );
  OAI221XL U1171 ( .A0(n317), .A1(n732), .B0(n176), .B1(n812), .C0(n1771), .Y(
        n2816) );
  OAI221XL U1172 ( .A0(n317), .A1(n730), .B0(n176), .B1(n810), .C0(n1773), .Y(
        n2818) );
  OAI221XL U1173 ( .A0(n318), .A1(n726), .B0(n177), .B1(n806), .C0(n1777), .Y(
        n2822) );
  OAI221XL U1174 ( .A0(n296), .A1(n823), .B0(n177), .B1(n850), .C0(n1728), .Y(
        n2772) );
  AOI21X1 U1175 ( .A0(N885), .A1(n196), .B0(n261), .Y(n1728) );
  OAI221XL U1176 ( .A0(n293), .A1(n819), .B0(n177), .B1(n846), .C0(n1732), .Y(
        n2776) );
  AOI21X1 U1177 ( .A0(N881), .A1(n197), .B0(n261), .Y(n1732) );
  OAI221XL U1178 ( .A0(n298), .A1(n816), .B0(n177), .B1(n843), .C0(n1735), .Y(
        n2779) );
  AOI21X1 U1179 ( .A0(N878), .A1(n202), .B0(n261), .Y(n1735) );
  OAI221XL U1180 ( .A0(n301), .A1(n815), .B0(n177), .B1(n842), .C0(n1736), .Y(
        n2780) );
  OAI221XL U1181 ( .A0(n311), .A1(n814), .B0(n177), .B1(n841), .C0(n1737), .Y(
        n2781) );
  OAI221XL U1182 ( .A0(n311), .A1(n812), .B0(n177), .B1(n839), .C0(n1739), .Y(
        n2783) );
  OAI221XL U1183 ( .A0(n312), .A1(n811), .B0(n177), .B1(n838), .C0(n1740), .Y(
        n2784) );
  OAI221XL U1184 ( .A0(n312), .A1(n810), .B0(n177), .B1(n837), .C0(n1741), .Y(
        n2785) );
  AOI21X1 U1185 ( .A0(N872), .A1(n195), .B0(n259), .Y(n1741) );
  OAI221XL U1186 ( .A0(n312), .A1(n809), .B0(n178), .B1(n836), .C0(n1742), .Y(
        n2786) );
  OAI221XL U1187 ( .A0(n313), .A1(n805), .B0(n176), .B1(n832), .C0(n1746), .Y(
        n2790) );
  OAI221XL U1188 ( .A0(n314), .A1(n802), .B0(n176), .B1(n829), .C0(n1749), .Y(
        n2793) );
  AOI21X1 U1189 ( .A0(N864), .A1(n205), .B0(n257), .Y(n1749) );
  OAI221XL U1190 ( .A0(n314), .A1(n801), .B0(n176), .B1(n828), .C0(n1750), .Y(
        n2794) );
  AOI21X1 U1191 ( .A0(N863), .A1(n197), .B0(n262), .Y(n1750) );
  OAI221XL U1192 ( .A0(n317), .A1(n733), .B0(n176), .B1(n813), .C0(n1770), .Y(
        n2815) );
  OAI221XL U1193 ( .A0(n318), .A1(n728), .B0(n176), .B1(n808), .C0(n1775), .Y(
        n2820) );
  OAI221XL U1194 ( .A0(n318), .A1(n727), .B0(n177), .B1(n807), .C0(n1776), .Y(
        n2821) );
  OAI221XL U1195 ( .A0(n319), .A1(n724), .B0(n178), .B1(n804), .C0(n1779), .Y(
        n2824) );
  AOI21X1 U1196 ( .A0(N834), .A1(n197), .B0(n262), .Y(n1779) );
  OAI221XL U1197 ( .A0(n293), .A1(n824), .B0(n177), .B1(n851), .C0(n1727), .Y(
        n2771) );
  OAI221XL U1198 ( .A0(n299), .A1(n818), .B0(n177), .B1(n845), .C0(n1733), .Y(
        n2777) );
  AOI21X1 U1199 ( .A0(N880), .A1(n195), .B0(n261), .Y(n1733) );
  OAI221XL U1200 ( .A0(n313), .A1(n806), .B0(n178), .B1(n833), .C0(n1745), .Y(
        n2789) );
  OAI221XL U1201 ( .A0(n313), .A1(n803), .B0(n176), .B1(n830), .C0(n1748), .Y(
        n2792) );
  AOI21X1 U1202 ( .A0(N865), .A1(n195), .B0(n260), .Y(n1748) );
  OAI221XL U1203 ( .A0(n295), .A1(n839), .B0(n178), .B1(n872), .C0(n1707), .Y(
        n2751) );
  AOI21X1 U1204 ( .A0(N906), .A1(n203), .B0(n260), .Y(n1707) );
  OAI221XL U1205 ( .A0(n301), .A1(n850), .B0(n178), .B1(n883), .C0(n1696), .Y(
        n2740) );
  OAI221XL U1206 ( .A0(n298), .A1(n848), .B0(n178), .B1(n881), .C0(n1698), .Y(
        n2742) );
  AOI21X1 U1207 ( .A0(N915), .A1(n201), .B0(n260), .Y(n1698) );
  OAI221XL U1208 ( .A0(n299), .A1(n846), .B0(n178), .B1(n879), .C0(n1700), .Y(
        n2744) );
  AOI21X1 U1209 ( .A0(N913), .A1(n721), .B0(n260), .Y(n1700) );
  OAI221XL U1210 ( .A0(n300), .A1(n843), .B0(n178), .B1(n876), .C0(n1703), .Y(
        n2747) );
  AOI21X1 U1211 ( .A0(N910), .A1(n202), .B0(n260), .Y(n1703) );
  OAI221XL U1212 ( .A0(n298), .A1(n841), .B0(n178), .B1(n874), .C0(n1705), .Y(
        n2749) );
  AOI21X1 U1213 ( .A0(N908), .A1(n200), .B0(n260), .Y(n1705) );
  OAI221XL U1214 ( .A0(n297), .A1(n837), .B0(n193), .B1(n870), .C0(n1709), .Y(
        n2753) );
  AOI21X1 U1215 ( .A0(N904), .A1(n195), .B0(n260), .Y(n1709) );
  OAI221XL U1216 ( .A0(n294), .A1(n836), .B0(n192), .B1(n869), .C0(n1710), .Y(
        n2754) );
  AOI21X1 U1217 ( .A0(N903), .A1(n195), .B0(n260), .Y(n1710) );
  OAI221XL U1218 ( .A0(n300), .A1(n834), .B0(n194), .B1(n867), .C0(n1712), .Y(
        n2756) );
  AOI21X1 U1219 ( .A0(N901), .A1(n202), .B0(n260), .Y(n1712) );
  OAI221XL U1220 ( .A0(n294), .A1(n832), .B0(n177), .B1(n865), .C0(n1714), .Y(
        n2758) );
  AOI21X1 U1221 ( .A0(N899), .A1(n202), .B0(n260), .Y(n1714) );
  OAI221XL U1222 ( .A0(n297), .A1(n829), .B0(n177), .B1(n862), .C0(n1717), .Y(
        n2761) );
  AOI21X1 U1223 ( .A0(N896), .A1(n206), .B0(n261), .Y(n1717) );
  OAI221XL U1224 ( .A0(n300), .A1(n828), .B0(n177), .B1(n861), .C0(n1718), .Y(
        n2762) );
  AOI21X1 U1225 ( .A0(N895), .A1(n199), .B0(n261), .Y(n1718) );
  OAI221XL U1226 ( .A0(n297), .A1(n840), .B0(n178), .B1(n873), .C0(n1706), .Y(
        n2750) );
  AOI21X1 U1227 ( .A0(N907), .A1(n721), .B0(n260), .Y(n1706) );
  OAI221XL U1228 ( .A0(n295), .A1(n838), .B0(n178), .B1(n871), .C0(n1708), .Y(
        n2752) );
  AOI21X1 U1229 ( .A0(N905), .A1(n205), .B0(n260), .Y(n1708) );
  OAI221XL U1230 ( .A0(n296), .A1(n842), .B0(n178), .B1(n875), .C0(n1704), .Y(
        n2748) );
  AOI21X1 U1231 ( .A0(N909), .A1(n200), .B0(n260), .Y(n1704) );
  NAND3BX1 U1232 ( .AN(n1849), .B(n392), .C(n391), .Y(n393) );
  INVX1 U1233 ( .A(n1859), .Y(n391) );
  OAI211X1 U1234 ( .A0(n289), .A1(n674), .B0(n673), .C0(n672), .Y(n2883) );
  INVXL U1235 ( .A(next_A[12]), .Y(n674) );
  OAI211X1 U1236 ( .A0(n293), .A1(n671), .B0(n670), .C0(n669), .Y(n2882) );
  INVX1 U1237 ( .A(next_A[13]), .Y(n671) );
  OAI211X1 U1238 ( .A0(n282), .A1(n682), .B0(n681), .C0(n680), .Y(n2886) );
  INVX1 U1239 ( .A(next_A[9]), .Y(n682) );
  OAI211X1 U1240 ( .A0(n288), .A1(n691), .B0(n690), .C0(n689), .Y(n2889) );
  NAND2X1 U1241 ( .A(N801), .B(n200), .Y(n690) );
  OAI211X1 U1242 ( .A0(n292), .A1(n695), .B0(n694), .C0(n693), .Y(n2890) );
  NAND2X1 U1243 ( .A(N800), .B(n203), .Y(n694) );
  OAI211X1 U1244 ( .A0(n287), .A1(n700), .B0(n699), .C0(n698), .Y(n2891) );
  NAND2X1 U1245 ( .A(n155), .B(n171), .Y(n699) );
  NAND2X1 U1246 ( .A(N799), .B(n203), .Y(n698) );
  OAI211X1 U1247 ( .A0(n292), .A1(n706), .B0(n705), .C0(n704), .Y(n2892) );
  NAND2X1 U1248 ( .A(n156), .B(n170), .Y(n705) );
  NAND2X1 U1249 ( .A(N798), .B(n199), .Y(n704) );
  OAI211X1 U1250 ( .A0(n286), .A1(n710), .B0(n709), .C0(n708), .Y(n2893) );
  INVX1 U1251 ( .A(next_A[2]), .Y(n710) );
  NAND2X1 U1252 ( .A(N797), .B(n201), .Y(n709) );
  OAI211X1 U1253 ( .A0(n291), .A1(n714), .B0(n713), .C0(n712), .Y(n2894) );
  OR3XL U1254 ( .A(n1849), .B(n390), .C(n389), .Y(n1456) );
  NAND2BX1 U1255 ( .AN(n581), .B(n580), .Y(n2829) );
  OAI21XL U1256 ( .A0(n799), .A1(n175), .B0(n677), .Y(n581) );
  XOR3X2 U1257 ( .A(n139), .B(n150), .C(n132), .Y(f3_A_32[7]) );
  XOR3X2 U1258 ( .A(n141), .B(n152), .C(n133), .Y(f3_A_32[5]) );
  XOR3X2 U1259 ( .A(n156), .B(n145), .C(n137), .Y(f3_A_32[1]) );
  XOR3X2 U1260 ( .A(n138), .B(n149), .C(n131), .Y(f3_A_32[8]) );
  XOR3X2 U1261 ( .A(n66), .B(n146), .C(n136), .Y(f3_A_32[11]) );
  XOR3X2 U1262 ( .A(n142), .B(n153), .C(n134), .Y(f3_A_32[4]) );
  XOR3X2 U1263 ( .A(SHA256_result[224]), .B(n147), .C(n137), .Y(f3_A_32[10])
         );
  XOR3X2 U1264 ( .A(n156), .B(n144), .C(n134), .Y(f3_A_32[13]) );
  OAI21XL U1265 ( .A0(n163), .A1(n78), .B0(n1785), .Y(n2830) );
  AOI22X1 U1266 ( .A0(N828), .A1(n200), .B0(n66), .B1(n269), .Y(n1785) );
  OAI21XL U1267 ( .A0(n166), .A1(n823), .B0(n1760), .Y(n2805) );
  AOI22X1 U1268 ( .A0(N853), .A1(n205), .B0(n134), .B1(n270), .Y(n1760) );
  OAI21XL U1269 ( .A0(n166), .A1(n816), .B0(n1767), .Y(n2812) );
  AOI22X1 U1270 ( .A0(N846), .A1(n197), .B0(n140), .B1(n269), .Y(n1767) );
  OAI21XL U1271 ( .A0(n166), .A1(n811), .B0(n1772), .Y(n2817) );
  AOI22X1 U1272 ( .A0(N841), .A1(n199), .B0(n145), .B1(n269), .Y(n1772) );
  OAI21XL U1273 ( .A0(n166), .A1(n809), .B0(n1774), .Y(n2819) );
  OAI21XL U1274 ( .A0(n165), .A1(n805), .B0(n1778), .Y(n2823) );
  OAI21XL U1275 ( .A0(n165), .A1(n803), .B0(n1780), .Y(n2825) );
  OAI21XL U1276 ( .A0(n165), .A1(n802), .B0(n1781), .Y(n2826) );
  OAI21XL U1277 ( .A0(n165), .A1(n801), .B0(n1782), .Y(n2827) );
  AOI22X1 U1278 ( .A0(N831), .A1(n199), .B0(n155), .B1(n269), .Y(n1782) );
  OAI21XL U1279 ( .A0(n166), .A1(n820), .B0(n1763), .Y(n2808) );
  AOI22X1 U1280 ( .A0(N850), .A1(n206), .B0(n137), .B1(n269), .Y(n1763) );
  OAI21XL U1281 ( .A0(n166), .A1(n817), .B0(n1766), .Y(n2811) );
  AOI22X1 U1282 ( .A0(N847), .A1(n717), .B0(n139), .B1(n269), .Y(n1766) );
  OAI21XL U1283 ( .A0(n165), .A1(n800), .B0(n1783), .Y(n2828) );
  NAND3BX1 U1284 ( .AN(n574), .B(n573), .C(n572), .Y(n2806) );
  OAI21XL U1285 ( .A0(n822), .A1(n175), .B0(n677), .Y(n574) );
  NAND2BX1 U1286 ( .AN(n325), .B(n135), .Y(n573) );
  NAND2X1 U1287 ( .A(N852), .B(n200), .Y(n572) );
  NAND3BX1 U1288 ( .AN(n577), .B(n576), .C(n575), .Y(n2807) );
  OAI21XL U1289 ( .A0(n821), .A1(n175), .B0(n677), .Y(n577) );
  NAND2X1 U1290 ( .A(N851), .B(n195), .Y(n575) );
  NAND2BX1 U1291 ( .AN(n325), .B(n136), .Y(n576) );
  NAND3BX1 U1292 ( .AN(n396), .B(n395), .C(n394), .Y(n2475) );
  NAND2BX1 U1293 ( .AN(n944), .B(n400), .Y(n394) );
  OAI21XL U1294 ( .A0(n265), .A1(n443), .B0(n677), .Y(n396) );
  NAND3BX1 U1295 ( .AN(n399), .B(n398), .C(n397), .Y(n2476) );
  NAND2BX1 U1296 ( .AN(n943), .B(n400), .Y(n397) );
  NAND2BX1 U1297 ( .AN(n49), .B(N1022), .Y(n398) );
  OAI21XL U1298 ( .A0(n265), .A1(n444), .B0(n677), .Y(n399) );
  NAND3BX1 U1299 ( .AN(n403), .B(n402), .C(n401), .Y(n2479) );
  NAND2BX1 U1300 ( .AN(n940), .B(n400), .Y(n401) );
  OAI21XL U1301 ( .A0(n277), .A1(n81), .B0(n677), .Y(n403) );
  NAND2BX1 U1302 ( .AN(n554), .B(n553), .Y(n2763) );
  OAI21XL U1303 ( .A0(n860), .A1(n175), .B0(n677), .Y(n554) );
  NAND2BX1 U1304 ( .AN(n556), .B(n555), .Y(n2765) );
  OAI21XL U1305 ( .A0(n858), .A1(n175), .B0(n677), .Y(n556) );
  NAND2BX1 U1306 ( .AN(n579), .B(n578), .Y(n2809) );
  OAI21XL U1307 ( .A0(n819), .A1(n175), .B0(n677), .Y(n579) );
  OAI2BB1X1 U1308 ( .A0N(N806), .A1N(n195), .B0(n676), .Y(n2884) );
  AOI2BB2X1 U1309 ( .B0(n170), .B1(n148), .A0N(n279), .A1N(n675), .Y(n676) );
  INVXL U1310 ( .A(next_A[11]), .Y(n675) );
  NAND2X1 U1311 ( .A(n719), .B(n718), .Y(n2895) );
  NAND2X1 U1312 ( .A(n679), .B(n678), .Y(n2885) );
  AOI21X1 U1313 ( .A0(n183), .A1(n149), .B0(n128), .Y(n678) );
  AOI22XL U1314 ( .A0(next_A[10]), .A1(n269), .B0(N805), .B1(n196), .Y(n679)
         );
  INVX1 U1315 ( .A(n703), .Y(n174) );
  XOR3X2 U1316 ( .A(n155), .B(n143), .C(n133), .Y(f3_A_32[14]) );
  XOR3X2 U1317 ( .A(n140), .B(n152), .C(n131), .Y(f3_A_32[17]) );
  XOR3X2 U1318 ( .A(SHA256_result[224]), .B(n150), .C(n138), .Y(f3_A_32[19])
         );
  XOR3X2 U1319 ( .A(n141), .B(n153), .C(n132), .Y(f3_A_32[16]) );
  XOR3X2 U1320 ( .A(n157), .B(n145), .C(n135), .Y(f3_A_32[12]) );
  NOR2X1 U1321 ( .A(round[2]), .B(round[3]), .Y(n2378) );
  AOI31X1 U1322 ( .A0(n2343), .A1(n2344), .A2(n2345), .B0(n233), .Y(N2956) );
  AOI2BB2X1 U1323 ( .B0(n2277), .B1(n346), .A0N(n797), .A1N(n2349), .Y(n2343)
         );
  AOI211X1 U1324 ( .A0(n2209), .A1(n343), .B0(n2346), .C0(n2347), .Y(n2345) );
  AOI31X1 U1325 ( .A0(n2327), .A1(n2328), .A2(n2329), .B0(n233), .Y(N2958) );
  NOR3BX1 U1326 ( .AN(n2333), .B(n2225), .C(n2231), .Y(n2328) );
  AOI211X1 U1327 ( .A0(n2334), .A1(n2312), .B0(n2335), .C0(n2152), .Y(n2327)
         );
  AOI211X1 U1328 ( .A0(n2209), .A1(n1393), .B0(n2330), .C0(n2331), .Y(n2329)
         );
  AOI31X1 U1329 ( .A0(n2270), .A1(n2271), .A2(n2272), .B0(n234), .Y(N2964) );
  AOI211X1 U1330 ( .A0(n2209), .A1(n1393), .B0(n2273), .C0(n2158), .Y(n2272)
         );
  AOI211X1 U1331 ( .A0(n31), .A1(n2275), .B0(n2124), .C0(n2198), .Y(n2271) );
  AOI31X1 U1332 ( .A0(n2387), .A1(n2388), .A2(n2389), .B0(n233), .Y(N2950) );
  AOI221X1 U1333 ( .A0(n2283), .A1(n159), .B0(n2234), .B1(n1396), .C0(n2380), 
        .Y(n2387) );
  NOR4BX1 U1334 ( .AN(n2390), .B(n2162), .C(n2247), .D(n2314), .Y(n2389) );
  AOI31X1 U1335 ( .A0(n2239), .A1(n748), .A2(n2240), .B0(n234), .Y(N2967) );
  AOI222X1 U1336 ( .A0(n2249), .A1(n1396), .B0(n41), .B1(n2251), .C0(n2139), 
        .C1(n2252), .Y(n2239) );
  INVX1 U1337 ( .A(n2245), .Y(n748) );
  AOI211X1 U1338 ( .A0(n2121), .A1(n114), .B0(n2242), .C0(n2243), .Y(n2240) );
  AOI31X1 U1339 ( .A0(n2316), .A1(n2317), .A2(n2318), .B0(n233), .Y(N2959) );
  AOI222X1 U1340 ( .A0(n2325), .A1(n1396), .B0(n2176), .B1(n161), .C0(n2305), 
        .C1(n2326), .Y(n2316) );
  AOI211X1 U1341 ( .A0(n160), .A1(n2319), .B0(n2320), .C0(n2321), .Y(n2318) );
  AOI31X1 U1342 ( .A0(n2405), .A1(n2406), .A2(n2407), .B0(n233), .Y(N2947) );
  NOR3X1 U1343 ( .A(n2136), .B(n2177), .C(n782), .Y(n2406) );
  AOI211X1 U1344 ( .A0(n2221), .A1(n41), .B0(n2408), .C0(n2331), .Y(n2407) );
  AOI31X1 U1345 ( .A0(n2125), .A1(n2126), .A2(n2127), .B0(n234), .Y(N2976) );
  AOI22X1 U1346 ( .A0(n2138), .A1(n2139), .B0(n2140), .B1(n346), .Y(n2125) );
  AOI222X1 U1347 ( .A0(n2134), .A1(n159), .B0(n2135), .B1(n2136), .C0(n2137), 
        .C1(round[1]), .Y(n2126) );
  AOI211X1 U1348 ( .A0(n2128), .A1(n112), .B0(n2130), .C0(n2131), .Y(n2127) );
  AOI31X1 U1349 ( .A0(n2260), .A1(n2261), .A2(n2262), .B0(n234), .Y(N2965) );
  AOI222X1 U1350 ( .A0(n114), .A1(n2251), .B0(n2267), .B1(n1393), .C0(n2268), 
        .C1(n2226), .Y(n2261) );
  NOR4BX1 U1351 ( .AN(n2263), .B(n2174), .C(n2264), .D(n2140), .Y(n2262) );
  INVX1 U1352 ( .A(output_enable), .Y(n387) );
  AOI31X1 U1353 ( .A0(n2381), .A1(n2382), .A2(n2383), .B0(n233), .Y(N2951) );
  NOR4BX1 U1354 ( .AN(n778), .B(n2209), .C(n2384), .D(n2177), .Y(n2383) );
  AOI221X1 U1355 ( .A0(n2325), .A1(n1393), .B0(n2294), .B1(round[1]), .C0(
        n2386), .Y(n2381) );
  AOI31X1 U1356 ( .A0(n2203), .A1(n2204), .A2(n2205), .B0(n234), .Y(N2970) );
  AOI2BB2X1 U1357 ( .B0(n347), .B1(n2209), .A0N(n2210), .A1N(n346), .Y(n2203)
         );
  AOI211X1 U1358 ( .A0(n2206), .A1(n1396), .B0(n2207), .C0(n2208), .Y(n2205)
         );
  AOI31X1 U1359 ( .A0(n2351), .A1(n2352), .A2(n2353), .B0(n233), .Y(N2955) );
  NOR4BX1 U1360 ( .AN(n2166), .B(n2314), .C(n2354), .D(n2355), .Y(n2353) );
  AOI22X1 U1361 ( .A0(n2174), .A1(n161), .B0(n41), .B1(n2356), .Y(n2352) );
  NOR2X1 U1362 ( .A(n2297), .B(n2347), .Y(n2351) );
  AOI31X1 U1363 ( .A0(n2211), .A1(n2212), .A2(n2213), .B0(n234), .Y(N2969) );
  NOR3X1 U1364 ( .A(n2224), .B(n2162), .C(n2225), .Y(n2212) );
  AOI31X1 U1365 ( .A0(n2307), .A1(n2308), .A2(n2309), .B0(n233), .Y(N2960) );
  NOR4BX1 U1366 ( .AN(n2310), .B(n2311), .C(n2312), .D(n2225), .Y(n2309) );
  AOI31X1 U1367 ( .A0(n2288), .A1(n2289), .A2(n2290), .B0(n234), .Y(N2962) );
  NOR4BX1 U1368 ( .AN(n2165), .B(n2291), .C(n2292), .D(n2293), .Y(n2290) );
  AOI211X1 U1369 ( .A0(n2161), .A1(n2138), .B0(n2295), .C0(n2296), .Y(n2289)
         );
  AOI21X1 U1370 ( .A0(n2198), .A1(n343), .B0(n2297), .Y(n2288) );
  AOI31X1 U1371 ( .A0(n2153), .A1(n2154), .A2(n2155), .B0(n234), .Y(N2974) );
  NOR3BX1 U1372 ( .AN(n2160), .B(n2161), .C(n2162), .Y(n2154) );
  NOR3BX1 U1373 ( .AN(n2156), .B(n2157), .C(n2158), .Y(n2155) );
  AOI31X1 U1374 ( .A0(n2410), .A1(n2411), .A2(n2412), .B0(n233), .Y(N2946) );
  AOI222X1 U1375 ( .A0(n41), .A1(n2220), .B0(n2350), .B1(n2139), .C0(n2175), 
        .C1(round[3]), .Y(n2410) );
  AND4X2 U1376 ( .A(n2413), .B(n768), .C(n2165), .D(n2132), .Y(n2412) );
  XOR3X2 U1377 ( .A(n155), .B(n146), .C(n135), .Y(f3_A_32[23]) );
  XOR3X2 U1378 ( .A(n157), .B(n148), .C(n137), .Y(f3_A_32[21]) );
  XOR3X2 U1379 ( .A(n156), .B(n147), .C(n136), .Y(f3_A_32[22]) );
  AOI21X1 U1380 ( .A0(n2374), .A1(n2375), .B0(n233), .Y(N2952) );
  AOI211X1 U1381 ( .A0(n2323), .A1(round[3]), .B0(n2379), .C0(n2380), .Y(n2374) );
  AOI211X1 U1382 ( .A0(n2363), .A1(round[1]), .B0(n2376), .C0(n2377), .Y(n2375) );
  OAI222XL U1383 ( .A0(n1396), .A1(n780), .B0(n159), .B1(n2149), .C0(n2138), 
        .C1(n791), .Y(n2379) );
  INVX1 U1384 ( .A(n130), .Y(n234) );
  INVX1 U1385 ( .A(n1978), .Y(n253) );
  XOR3X2 U1386 ( .A(n154), .B(n145), .C(n134), .Y(f3_A_32[24]) );
  XOR3X2 U1387 ( .A(n142), .B(n151), .C(n132), .Y(f3_A_32[27]) );
  XOR3X2 U1388 ( .A(n144), .B(n153), .C(n133), .Y(f3_A_32[25]) );
  INVX1 U1389 ( .A(n2140), .Y(n753) );
  OAI211X1 U1390 ( .A0(round[2]), .A1(n753), .B0(n2210), .C0(n2233), .Y(n2331)
         );
  NOR2X1 U1391 ( .A(n793), .B(n343), .Y(n2342) );
  INVX1 U1392 ( .A(n2315), .Y(n762) );
  NAND3X1 U1393 ( .A(n749), .B(n2133), .C(n2156), .Y(n2297) );
  NOR2X1 U1394 ( .A(n343), .B(n785), .Y(n2322) );
  XOR3X2 U1395 ( .A(n141), .B(n150), .C(n131), .Y(f3_A_32[28]) );
  XOR3X2 U1396 ( .A(n158), .B(n148), .C(n139), .Y(f3_A_32[30]) );
  OAI2BB1X1 U1397 ( .A0N(n160), .A1N(n2302), .B0(n759), .Y(n2282) );
  INVX1 U1398 ( .A(n2139), .Y(n796) );
  INVX1 U1399 ( .A(n2226), .Y(n794) );
  OAI2BB1X1 U1400 ( .A0N(round[1]), .A1N(n2304), .B0(n2403), .Y(n2402) );
  AOI31X1 U1401 ( .A0(n776), .A1(n790), .A2(n2274), .B0(n161), .Y(n2404) );
  NOR3X1 U1402 ( .A(n346), .B(n161), .C(n794), .Y(n2314) );
  NOR2X1 U1403 ( .A(n159), .B(n160), .Y(n2305) );
  OAI222XL U1404 ( .A0(n769), .A1(n783), .B0(n2313), .B1(n756), .C0(n31), .C1(
        n750), .Y(n2311) );
  NOR2X1 U1405 ( .A(n2136), .B(n2305), .Y(n2313) );
  OAI222XL U1406 ( .A0(n159), .A1(n755), .B0(n781), .B1(n760), .C0(round[1]), 
        .C1(n2159), .Y(n2157) );
  NOR3X1 U1407 ( .A(n347), .B(round[2]), .C(n791), .Y(n2312) );
  OAI222XL U1408 ( .A0(n161), .A1(n2372), .B0(n765), .B1(n780), .C0(round[1]), 
        .C1(n772), .Y(n2368) );
  NOR2X1 U1409 ( .A(n2166), .B(round[2]), .Y(n2225) );
  OAI222XL U1410 ( .A0(n127), .A1(n2173), .B0(n2396), .B1(n784), .C0(n2409), 
        .C1(n765), .Y(n2408) );
  INVX1 U1411 ( .A(n2267), .Y(n784) );
  NOR3X1 U1412 ( .A(n2232), .B(n31), .C(n2324), .Y(n2409) );
  NOR2X1 U1413 ( .A(n2175), .B(n2177), .Y(n2244) );
  OAI31X1 U1414 ( .A0(n764), .A1(n160), .A2(round[3]), .B0(n2265), .Y(n2264)
         );
  AOI31X1 U1415 ( .A0(n765), .A1(n796), .A2(n41), .B0(n2266), .Y(n2265) );
  NOR2X1 U1416 ( .A(n781), .B(round[3]), .Y(n2176) );
  NOR3X1 U1417 ( .A(n161), .B(n159), .C(n793), .Y(n2293) );
  NAND2X1 U1418 ( .A(n2398), .B(n161), .Y(n2159) );
  NOR2X1 U1419 ( .A(n756), .B(round[2]), .Y(n2221) );
  NOR2X1 U1420 ( .A(n765), .B(round[2]), .Y(n2220) );
  NOR2X1 U1421 ( .A(n777), .B(round[2]), .Y(n2137) );
  OAI221XL U1422 ( .A0(n777), .A1(n2149), .B0(n765), .B1(n778), .C0(n2332), 
        .Y(n2330) );
  OAI21XL U1423 ( .A0(n2183), .A1(n2191), .B0(n32), .Y(n2332) );
  NOR2X1 U1424 ( .A(n777), .B(round[3]), .Y(n2189) );
  OAI211X1 U1426 ( .A0(n159), .A1(n764), .B0(n746), .C0(n758), .Y(n2201) );
  OAI22X1 U1427 ( .A0(n343), .A1(n789), .B0(n775), .B1(n127), .Y(n2347) );
  NOR3X1 U1428 ( .A(n343), .B(n159), .C(n796), .Y(n2373) );
  AOI221X1 U1429 ( .A0(n747), .A1(n159), .B0(n160), .B1(round[1]), .C0(n2350), 
        .Y(n2349) );
  NAND2X1 U1430 ( .A(n112), .B(n2139), .Y(n2149) );
  INVX1 U1431 ( .A(n31), .Y(n781) );
  NOR2X1 U1432 ( .A(n788), .B(round[3]), .Y(n2398) );
  AOI211X1 U1433 ( .A0(n160), .A1(n2257), .B0(n2177), .C0(n2144), .Y(n2256) );
  OAI21XL U1434 ( .A0(n347), .A1(n794), .B0(n760), .Y(n2257) );
  NOR2X1 U1435 ( .A(n2274), .B(n769), .Y(n2231) );
  AOI31X1 U1436 ( .A0(n774), .A1(n780), .A2(n2173), .B0(n769), .Y(n2172) );
  INVX1 U1437 ( .A(n2136), .Y(n780) );
  NOR2X1 U1438 ( .A(n777), .B(n343), .Y(n2252) );
  NOR2X1 U1439 ( .A(n756), .B(n159), .Y(n2258) );
  OAI211X1 U1440 ( .A0(n159), .A1(round[2]), .B0(n776), .C0(n786), .Y(n2285)
         );
  INVX1 U1441 ( .A(n2128), .Y(n786) );
  NOR2X1 U1442 ( .A(n343), .B(n791), .Y(n2248) );
  NAND2X1 U1443 ( .A(n2248), .B(round[3]), .Y(n2165) );
  OAI211X1 U1444 ( .A0(n769), .A1(n775), .B0(n766), .C0(n2133), .Y(n2130) );
  NOR2X1 U1445 ( .A(n794), .B(n160), .Y(n2195) );
  OAI211X1 U1446 ( .A0(n2341), .A1(n1396), .B0(n2160), .C0(n770), .Y(n2339) );
  AOI21X1 U1447 ( .A0(n31), .A1(n793), .B0(n2267), .Y(n2341) );
  OAI2BB2X1 U1448 ( .B0(n347), .B1(n2274), .A0N(n1396), .A1N(n2144), .Y(n2158)
         );
  NOR2X1 U1449 ( .A(n796), .B(n161), .Y(n2286) );
  NOR2X1 U1450 ( .A(n796), .B(n160), .Y(n2232) );
  OAI21XL U1451 ( .A0(n161), .A1(n797), .B0(n764), .Y(n2326) );
  OAI22X1 U1452 ( .A0(n1985), .A1(n901), .B0(n1984), .B1(n550), .Y(n386) );
  OAI22X1 U1453 ( .A0(n895), .A1(n1984), .B0(n907), .B1(n1985), .Y(n2037) );
  OAI22X1 U1454 ( .A0(n896), .A1(n1984), .B0(n908), .B1(n1985), .Y(n2033) );
  OAI22X1 U1455 ( .A0(n897), .A1(n1984), .B0(n909), .B1(n1985), .Y(n2029) );
  OAI22X1 U1456 ( .A0(n898), .A1(n1984), .B0(n910), .B1(n1985), .Y(n2025) );
  OAI22X1 U1457 ( .A0(n1985), .A1(n442), .B0(n246), .B1(n531), .Y(n358) );
  OAI21XL U1458 ( .A0(n159), .A1(n795), .B0(n2166), .Y(n2116) );
  OAI22X1 U1459 ( .A0(n889), .A1(n1984), .B0(n905), .B1(n244), .Y(n2061) );
  OAI22X1 U1460 ( .A0(n894), .A1(n1984), .B0(n906), .B1(n244), .Y(n2041) );
  OAI22X1 U1461 ( .A0(n1985), .A1(n904), .B0(n246), .B1(n506), .Y(n370) );
  INVX1 U1462 ( .A(n2323), .Y(n745) );
  NAND2BX1 U1463 ( .AN(n2173), .B(n112), .Y(n2263) );
  OAI22X1 U1464 ( .A0(n1985), .A1(n902), .B0(n246), .B1(n524), .Y(n362) );
  OAI22X1 U1465 ( .A0(n1985), .A1(n903), .B0(n246), .B1(n510), .Y(n368) );
  OAI22X1 U1466 ( .A0(n1985), .A1(n912), .B0(n1984), .B1(n440), .Y(n384) );
  NOR3X1 U1467 ( .A(n793), .B(n161), .C(n781), .Y(n2186) );
  INVX1 U1468 ( .A(n2234), .Y(n779) );
  NAND2X1 U1469 ( .A(n2144), .B(n161), .Y(n2333) );
  NAND2X1 U1470 ( .A(n2226), .B(n114), .Y(n2132) );
  NAND2X1 U1471 ( .A(n2121), .B(n31), .Y(n2372) );
  NOR2X1 U1472 ( .A(n789), .B(round[3]), .Y(n2150) );
  NOR2X1 U1473 ( .A(n2159), .B(round[2]), .Y(n2294) );
  AOI21X1 U1474 ( .A0(n2133), .A1(n786), .B0(n1396), .Y(n2361) );
  NAND3BX1 U1475 ( .AN(n2150), .B(n785), .C(n2269), .Y(n2215) );
  NAND3X1 U1476 ( .A(round[3]), .B(n1396), .C(n31), .Y(n2269) );
  CLKINVX3 U1477 ( .A(n1393), .Y(n347) );
  NAND3X1 U1478 ( .A(n752), .B(n2200), .C(n2385), .Y(n2384) );
  OAI21XL U1479 ( .A0(n2315), .A1(n2283), .B0(n159), .Y(n2385) );
  INVX1 U1480 ( .A(n2287), .Y(n775) );
  OAI221XL U1481 ( .A0(round[1]), .A1(n2146), .B0(round[2]), .B1(n757), .C0(
        n2147), .Y(n2145) );
  OAI21XL U1482 ( .A0(n2148), .A1(n782), .B0(n161), .Y(n2147) );
  OAI21XL U1483 ( .A0(n2118), .A1(n159), .B0(n2119), .Y(n2117) );
  OAI21XL U1484 ( .A0(n116), .A1(n2121), .B0(n2122), .Y(n2119) );
  AOI2BB1X1 U1485 ( .A0N(n2144), .A1N(n2176), .B0(n769), .Y(n2355) );
  AOI21X1 U1486 ( .A0(n2166), .A1(n780), .B0(n161), .Y(n2163) );
  AOI21X1 U1487 ( .A0(n2199), .A1(n786), .B0(n343), .Y(n2335) );
  AOI21X1 U1488 ( .A0(n753), .A1(n751), .B0(round[2]), .Y(n2208) );
  INVX1 U1489 ( .A(n2202), .Y(n773) );
  INVX1 U1490 ( .A(n2206), .Y(n783) );
  NAND3BX1 U1491 ( .AN(n2198), .B(n2199), .C(n2200), .Y(n2196) );
  NAND3X1 U1492 ( .A(n2216), .B(n2217), .C(n2218), .Y(n2214) );
  OAI21XL U1493 ( .A0(n2221), .A1(n116), .B0(n31), .Y(n2216) );
  OAI21XL U1494 ( .A0(n2219), .A1(n2220), .B0(n160), .Y(n2218) );
  OAI21XL U1495 ( .A0(n2128), .A1(n2174), .B0(n2138), .Y(n2217) );
  AOI2BB1X1 U1496 ( .A0N(n2174), .A1N(n2161), .B0(n161), .Y(n2414) );
  AOI2BB1X1 U1497 ( .A0N(n2144), .A1N(n2324), .B0(n347), .Y(n2377) );
  XOR3X2 U1498 ( .A(n66), .B(n147), .C(n138), .Y(f3_A_32[31]) );
  OR2X2 U1499 ( .A(n343), .B(n347), .Y(n127) );
  INVX1 U1500 ( .A(n127), .Y(n2138) );
  INVX1 U1501 ( .A(n41), .Y(n777) );
  NOR3X1 U1502 ( .A(n765), .B(n159), .C(round[3]), .Y(n2354) );
  NAND2X1 U1503 ( .A(n114), .B(n343), .Y(n2223) );
  OAI21XL U1504 ( .A0(n159), .A1(n345), .B0(n2223), .Y(n2364) );
  INVX1 U1505 ( .A(n1984), .Y(n247) );
  NOR2X1 U1506 ( .A(n160), .B(n769), .Y(n2397) );
  INVX1 U1507 ( .A(n33), .Y(n239) );
  INVX1 U1508 ( .A(n34), .Y(n254) );
  INVX1 U1509 ( .A(n1986), .Y(n243) );
  INVX1 U1510 ( .A(n1982), .Y(n250) );
  INVX1 U1511 ( .A(n35), .Y(n237) );
  INVX1 U1512 ( .A(n134), .Y(n630) );
  INVX1 U1513 ( .A(n137), .Y(n642) );
  INVX1 U1514 ( .A(n136), .Y(n638) );
  INVX1 U1515 ( .A(n148), .Y(n728) );
  INVX1 U1516 ( .A(n152), .Y(n724) );
  INVX1 U1517 ( .A(n142), .Y(n734) );
  INVX1 U1518 ( .A(n138), .Y(n738) );
  INVX1 U1519 ( .A(n141), .Y(n735) );
  INVX1 U1520 ( .A(n146), .Y(n730) );
  INVX1 U1521 ( .A(n149), .Y(n727) );
  INVX1 U1522 ( .A(n150), .Y(n726) );
  INVX1 U1523 ( .A(n143), .Y(n733) );
  INVX1 U1524 ( .A(n144), .Y(n732) );
  INVX1 U1525 ( .A(n132), .Y(n741) );
  INVX1 U1526 ( .A(n133), .Y(n739) );
  INVX1 U1527 ( .A(n158), .Y(n720) );
  INVX1 U1528 ( .A(n157), .Y(n707) );
  NAND2X1 U1529 ( .A(H4[29]), .B(n219), .Y(n451) );
  INVX1 U1530 ( .A(inner_busy), .Y(n348) );
  OAI211XL U1531 ( .A0(n23), .A1(n445), .B0(n56), .C0(n1609), .Y(n2668) );
  OAI211X1 U1532 ( .A0(n21), .A1(n531), .B0(n57), .C0(n1592), .Y(n2634) );
  NAND2X1 U1533 ( .A(H4[4]), .B(n215), .Y(n1592) );
  OAI211X1 U1534 ( .A0(n21), .A1(n535), .B0(n62), .C0(n1593), .Y(n2635) );
  NAND2X1 U1535 ( .A(H4[3]), .B(n215), .Y(n1593) );
  OAI211X1 U1536 ( .A0(n20), .A1(n72), .B0(n57), .C0(n1594), .Y(n2636) );
  NAND2X1 U1537 ( .A(H4[2]), .B(n215), .Y(n1594) );
  OAI211X1 U1538 ( .A0(n22), .A1(n935), .B0(n57), .C0(n1524), .Y(n2514) );
  OAI211X1 U1539 ( .A0(n19), .A1(n934), .B0(n61), .C0(n1525), .Y(n2515) );
  NAND2X1 U1540 ( .A(H6[27]), .B(n223), .Y(n1525) );
  OAI211X1 U1541 ( .A0(n24), .A1(n932), .B0(n55), .C0(n1527), .Y(n2517) );
  NAND2X1 U1542 ( .A(H6[25]), .B(n223), .Y(n1527) );
  OAI211X1 U1543 ( .A0(n19), .A1(n931), .B0(n58), .C0(n1528), .Y(n2518) );
  NAND2X1 U1544 ( .A(H6[24]), .B(n223), .Y(n1528) );
  OAI211X1 U1545 ( .A0(n21), .A1(n930), .B0(n59), .C0(n1529), .Y(n2519) );
  NAND2X1 U1546 ( .A(H6[23]), .B(n223), .Y(n1529) );
  OAI211X1 U1547 ( .A0(n18), .A1(n922), .B0(n58), .C0(n1532), .Y(n2527) );
  NAND2X1 U1548 ( .A(H6[15]), .B(n222), .Y(n1532) );
  OAI211X1 U1549 ( .A0(n20), .A1(n921), .B0(n60), .C0(n1533), .Y(n2528) );
  NAND2X1 U1550 ( .A(H6[14]), .B(n222), .Y(n1533) );
  OAI211X1 U1551 ( .A0(n20), .A1(n890), .B0(n60), .C0(n1587), .Y(n2624) );
  NAND2X1 U1552 ( .A(H4[14]), .B(n216), .Y(n1587) );
  OAI211X1 U1553 ( .A0(n21), .A1(n900), .B0(n61), .C0(n1583), .Y(n2614) );
  NAND2X1 U1554 ( .A(H4[24]), .B(n216), .Y(n1583) );
  OAI211X1 U1555 ( .A0(n21), .A1(n894), .B0(n60), .C0(n1585), .Y(n2620) );
  NAND2X1 U1556 ( .A(H4[18]), .B(n216), .Y(n1585) );
  OAI211X1 U1557 ( .A0(n20), .A1(n70), .B0(n60), .C0(n1596), .Y(n2638) );
  NAND2X1 U1558 ( .A(H4[0]), .B(n215), .Y(n1596) );
  OAI211X1 U1559 ( .A0(n21), .A1(n819), .B0(n58), .C0(n1793), .Y(n2841) );
  NAND2X1 U1560 ( .A(H1[22]), .B(n214), .Y(n1793) );
  OAI211X1 U1561 ( .A0(n22), .A1(n906), .B0(n58), .C0(n1602), .Y(n2652) );
  NAND2X1 U1562 ( .A(H5[18]), .B(n215), .Y(n1602) );
  OAI211X1 U1563 ( .A0(n18), .A1(n905), .B0(n57), .C0(n1605), .Y(n2657) );
  NAND2X1 U1564 ( .A(H5[13]), .B(n214), .Y(n1605) );
  OAI211X1 U1565 ( .A0(n18), .A1(n542), .B0(n58), .C0(n1595), .Y(n2637) );
  NAND2X1 U1566 ( .A(H4[1]), .B(n215), .Y(n1595) );
  OAI211X1 U1567 ( .A0(n22), .A1(n888), .B0(n58), .C0(n1588), .Y(n2626) );
  NAND2X1 U1568 ( .A(H4[12]), .B(n216), .Y(n1588) );
  OAI211X1 U1569 ( .A0(n17), .A1(n84), .B0(n54), .C0(n1591), .Y(n2633) );
  NAND2X1 U1570 ( .A(H4[5]), .B(n216), .Y(n1591) );
  NAND2X1 U1571 ( .A(H5[3]), .B(n214), .Y(n1608) );
  OAI211X1 U1572 ( .A0(n19), .A1(n1140), .B0(n58), .C0(n1598), .Y(n2642) );
  NAND2X1 U1573 ( .A(H5[28]), .B(n215), .Y(n1598) );
  OAI211X1 U1574 ( .A0(n18), .A1(n1141), .B0(n54), .C0(n1599), .Y(n2643) );
  NAND2X1 U1575 ( .A(H5[27]), .B(n215), .Y(n1599) );
  OAI211X1 U1576 ( .A0(n18), .A1(n1143), .B0(n58), .C0(n1600), .Y(n2645) );
  NAND2X1 U1577 ( .A(H5[25]), .B(n215), .Y(n1600) );
  OAI211X1 U1578 ( .A0(n19), .A1(n1157), .B0(n56), .C0(n1606), .Y(n2659) );
  NAND2X1 U1579 ( .A(H5[11]), .B(n214), .Y(n1606) );
  NAND2X1 U1580 ( .A(H4[9]), .B(n216), .Y(n1589) );
  NAND2X1 U1581 ( .A(H4[6]), .B(n216), .Y(n1590) );
  OAI211X1 U1582 ( .A0(n23), .A1(n933), .B0(n57), .C0(n1526), .Y(n2516) );
  NAND2X1 U1583 ( .A(H6[26]), .B(n223), .Y(n1526) );
  OAI211X1 U1584 ( .A0(n24), .A1(n924), .B0(n60), .C0(n1530), .Y(n2525) );
  NAND2X1 U1585 ( .A(H6[17]), .B(n222), .Y(n1530) );
  OAI211X1 U1586 ( .A0(n20), .A1(n923), .B0(n55), .C0(n1531), .Y(n2526) );
  NAND2X1 U1587 ( .A(H6[16]), .B(n222), .Y(n1531) );
  OAI211X1 U1588 ( .A0(n21), .A1(n919), .B0(n62), .C0(n1534), .Y(n2530) );
  NAND2X1 U1589 ( .A(H6[12]), .B(n221), .Y(n1534) );
  OAI211X1 U1590 ( .A0(n24), .A1(n826), .B0(n59), .C0(n1788), .Y(n2834) );
  NAND2X1 U1591 ( .A(H1[29]), .B(n214), .Y(n1788) );
  OAI211X1 U1592 ( .A0(n20), .A1(n825), .B0(n54), .C0(n1789), .Y(n2835) );
  NAND2X1 U1593 ( .A(H1[28]), .B(n214), .Y(n1789) );
  OAI211X1 U1594 ( .A0(n24), .A1(n824), .B0(n60), .C0(n1790), .Y(n2836) );
  NAND2X1 U1595 ( .A(H1[27]), .B(n214), .Y(n1790) );
  OAI211X1 U1596 ( .A0(n21), .A1(n818), .B0(n57), .C0(n1794), .Y(n2842) );
  NAND2X1 U1597 ( .A(H1[21]), .B(n214), .Y(n1794) );
  OAI211X1 U1598 ( .A0(n24), .A1(n815), .B0(n55), .C0(n1795), .Y(n2845) );
  NAND2X1 U1599 ( .A(H1[18]), .B(n213), .Y(n1795) );
  OAI211X1 U1600 ( .A0(n22), .A1(n814), .B0(n57), .C0(n1796), .Y(n2846) );
  NAND2X1 U1601 ( .A(H1[17]), .B(n213), .Y(n1796) );
  OAI211X1 U1602 ( .A0(n23), .A1(n812), .B0(n57), .C0(n1798), .Y(n2848) );
  NAND2X1 U1603 ( .A(H1[15]), .B(n213), .Y(n1798) );
  OAI211X1 U1604 ( .A0(n18), .A1(n810), .B0(n55), .C0(n1799), .Y(n2850) );
  NAND2X1 U1605 ( .A(H1[13]), .B(n213), .Y(n1799) );
  OAI211X1 U1606 ( .A0(n24), .A1(n893), .B0(n57), .C0(n1586), .Y(n2621) );
  NAND2X1 U1607 ( .A(H4[17]), .B(n216), .Y(n1586) );
  NAND2X1 U1608 ( .A(H4[28]), .B(n216), .Y(n1582) );
  OAI211X1 U1609 ( .A0(n22), .A1(n895), .B0(n57), .C0(n1584), .Y(n2619) );
  NAND2X1 U1610 ( .A(H4[19]), .B(n216), .Y(n1584) );
  OAI211X1 U1611 ( .A0(n19), .A1(n853), .B0(n56), .C0(n1543), .Y(n2546) );
  NAND2X1 U1612 ( .A(H2[29]), .B(n220), .Y(n1543) );
  OAI211X1 U1613 ( .A0(n20), .A1(n850), .B0(n54), .C0(n1546), .Y(n2549) );
  NAND2X1 U1614 ( .A(H2[26]), .B(n219), .Y(n1546) );
  OAI211X1 U1615 ( .A0(n18), .A1(n846), .B0(n61), .C0(n1547), .Y(n2553) );
  NAND2X1 U1616 ( .A(H2[22]), .B(n219), .Y(n1547) );
  OAI211X1 U1617 ( .A0(n17), .A1(n843), .B0(n56), .C0(n1549), .Y(n2556) );
  NAND2X1 U1618 ( .A(H2[19]), .B(n219), .Y(n1549) );
  OAI211X1 U1619 ( .A0(n24), .A1(n842), .B0(n62), .C0(n1550), .Y(n2557) );
  NAND2X1 U1620 ( .A(H2[18]), .B(n219), .Y(n1550) );
  OAI211X1 U1621 ( .A0(n19), .A1(n841), .B0(n60), .C0(n1551), .Y(n2558) );
  NAND2X1 U1622 ( .A(H2[17]), .B(n219), .Y(n1551) );
  OAI211X1 U1623 ( .A0(n18), .A1(n839), .B0(n60), .C0(n1552), .Y(n2560) );
  NAND2X1 U1624 ( .A(H2[15]), .B(n219), .Y(n1552) );
  OAI211X1 U1625 ( .A0(n17), .A1(n838), .B0(n54), .C0(n1553), .Y(n2561) );
  NAND2X1 U1626 ( .A(H2[14]), .B(n218), .Y(n1553) );
  OAI211X1 U1627 ( .A0(n24), .A1(n837), .B0(n62), .C0(n1554), .Y(n2562) );
  NAND2X1 U1628 ( .A(H2[13]), .B(n218), .Y(n1554) );
  OAI211X1 U1629 ( .A0(n22), .A1(n836), .B0(n60), .C0(n1555), .Y(n2563) );
  NAND2X1 U1630 ( .A(H2[12]), .B(n218), .Y(n1555) );
  NAND2X1 U1631 ( .A(H2[5]), .B(n218), .Y(n1559) );
  NAND2X1 U1632 ( .A(H2[4]), .B(n218), .Y(n1560) );
  NAND2X1 U1633 ( .A(H4[30]), .B(n216), .Y(n1581) );
  OAI211X1 U1634 ( .A0(n17), .A1(n1144), .B0(n58), .C0(n1601), .Y(n2646) );
  NAND2X1 U1635 ( .A(H5[24]), .B(n215), .Y(n1601) );
  OAI211X1 U1636 ( .A0(n23), .A1(n1152), .B0(n54), .C0(n1603), .Y(n2654) );
  NAND2X1 U1637 ( .A(H5[16]), .B(n215), .Y(n1603) );
  OAI211X1 U1638 ( .A0(n23), .A1(n1154), .B0(n55), .C0(n1604), .Y(n2656) );
  NAND2X1 U1639 ( .A(H5[14]), .B(n215), .Y(n1604) );
  OAI211X1 U1640 ( .A0(n24), .A1(n88), .B0(n56), .C0(n1805), .Y(n2863) );
  OAI211X1 U1641 ( .A0(n19), .A1(n822), .B0(n58), .C0(n1791), .Y(n2838) );
  NAND2X1 U1642 ( .A(H1[25]), .B(n214), .Y(n1791) );
  OAI211X1 U1643 ( .A0(n18), .A1(n821), .B0(n56), .C0(n1792), .Y(n2839) );
  NAND2X1 U1644 ( .A(H1[24]), .B(n214), .Y(n1792) );
  NAND2X1 U1645 ( .A(H1[2]), .B(n213), .Y(n1804) );
  OAI211X1 U1646 ( .A0(n21), .A1(n901), .B0(n62), .C0(n1597), .Y(n2639) );
  NAND2X1 U1647 ( .A(H5[31]), .B(n215), .Y(n1597) );
  NAND2X1 U1648 ( .A(n71), .B(n216), .Y(n1580) );
  OAI211X1 U1649 ( .A0(n17), .A1(n813), .B0(n62), .C0(n1797), .Y(n2847) );
  NAND2X1 U1650 ( .A(H1[16]), .B(n213), .Y(n1797) );
  NAND2X1 U1651 ( .A(H1[10]), .B(n213), .Y(n1801) );
  NAND2X1 U1652 ( .A(H1[31]), .B(n214), .Y(n1787) );
  OAI211X1 U1653 ( .A0(n18), .A1(n852), .B0(n57), .C0(n1544), .Y(n2547) );
  NAND2X1 U1654 ( .A(H2[28]), .B(n220), .Y(n1544) );
  OAI211X1 U1655 ( .A0(n19), .A1(n851), .B0(n61), .C0(n1545), .Y(n2548) );
  NAND2X1 U1656 ( .A(H2[27]), .B(n220), .Y(n1545) );
  OAI211X1 U1657 ( .A0(n22), .A1(n845), .B0(n62), .C0(n1548), .Y(n2554) );
  NAND2X1 U1658 ( .A(H2[21]), .B(n219), .Y(n1548) );
  NAND2X1 U1659 ( .A(H2[9]), .B(n218), .Y(n1556) );
  NAND2X1 U1660 ( .A(H2[6]), .B(n218), .Y(n1558) );
  OAI211X1 U1661 ( .A0(n19), .A1(n872), .B0(n54), .C0(n1571), .Y(n2591) );
  NAND2X1 U1662 ( .A(H3[15]), .B(n217), .Y(n1571) );
  OAI211X1 U1663 ( .A0(n20), .A1(n883), .B0(n58), .C0(n1564), .Y(n2580) );
  NAND2X1 U1664 ( .A(H3[26]), .B(n218), .Y(n1564) );
  OAI211X1 U1665 ( .A0(n24), .A1(n881), .B0(n59), .C0(n1565), .Y(n2582) );
  NAND2X1 U1666 ( .A(H3[24]), .B(n218), .Y(n1565) );
  OAI211X1 U1667 ( .A0(n21), .A1(n886), .B0(n61), .C0(n1563), .Y(n2577) );
  NAND2X1 U1668 ( .A(H3[29]), .B(n218), .Y(n1563) );
  OAI211X1 U1669 ( .A0(n21), .A1(n879), .B0(n62), .C0(n1566), .Y(n2584) );
  NAND2X1 U1670 ( .A(H3[22]), .B(n217), .Y(n1566) );
  OAI211X1 U1671 ( .A0(n19), .A1(n876), .B0(n55), .C0(n1567), .Y(n2587) );
  NAND2X1 U1672 ( .A(H3[19]), .B(n217), .Y(n1567) );
  OAI211X1 U1673 ( .A0(n23), .A1(n874), .B0(n61), .C0(n1569), .Y(n2589) );
  NAND2X1 U1674 ( .A(H3[17]), .B(n217), .Y(n1569) );
  OAI211X1 U1675 ( .A0(n18), .A1(n870), .B0(n60), .C0(n1573), .Y(n2593) );
  NAND2X1 U1676 ( .A(H3[13]), .B(n217), .Y(n1573) );
  OAI211X1 U1677 ( .A0(n20), .A1(n869), .B0(n61), .C0(n1574), .Y(n2594) );
  NAND2X1 U1678 ( .A(H3[12]), .B(n217), .Y(n1574) );
  NAND2X1 U1679 ( .A(H3[8]), .B(n217), .Y(n1576) );
  NAND2X1 U1680 ( .A(H3[5]), .B(n217), .Y(n1577) );
  NAND2X1 U1681 ( .A(H3[4]), .B(n217), .Y(n1578) );
  NAND2X1 U1682 ( .A(H3[31]), .B(n218), .Y(n1562) );
  OAI211X1 U1683 ( .A0(n20), .A1(n970), .B0(n61), .C0(n1438), .Y(n2417) );
  NAND2X1 U1684 ( .A(H7[30]), .B(n222), .Y(n1438) );
  OAI211X1 U1685 ( .A0(n20), .A1(n968), .B0(n55), .C0(n1439), .Y(n2419) );
  NAND2X1 U1686 ( .A(H7[28]), .B(n222), .Y(n1439) );
  OAI211X1 U1687 ( .A0(n17), .A1(n967), .B0(n56), .C0(n1440), .Y(n2420) );
  NAND2X1 U1688 ( .A(H7[27]), .B(n222), .Y(n1440) );
  OAI211X1 U1689 ( .A0(n20), .A1(n965), .B0(n54), .C0(n1441), .Y(n2422) );
  NAND2X1 U1690 ( .A(H7[25]), .B(n222), .Y(n1441) );
  OAI211X1 U1691 ( .A0(n19), .A1(n873), .B0(n56), .C0(n1570), .Y(n2590) );
  NAND2X1 U1692 ( .A(H3[16]), .B(n219), .Y(n1570) );
  OAI211X1 U1693 ( .A0(n17), .A1(n871), .B0(n62), .C0(n1572), .Y(n2592) );
  NAND2X1 U1694 ( .A(H3[14]), .B(n217), .Y(n1572) );
  OAI211X1 U1695 ( .A0(n19), .A1(n964), .B0(n60), .C0(n1442), .Y(n2423) );
  NAND2X1 U1696 ( .A(H7[24]), .B(n222), .Y(n1442) );
  OAI211X1 U1697 ( .A0(n22), .A1(n963), .B0(n55), .C0(n1443), .Y(n2424) );
  NAND2X1 U1698 ( .A(H7[23]), .B(n222), .Y(n1443) );
  OAI211X1 U1699 ( .A0(n22), .A1(n962), .B0(n59), .C0(n1444), .Y(n2425) );
  NAND2X1 U1700 ( .A(H7[22]), .B(n222), .Y(n1444) );
  OAI211X1 U1701 ( .A0(n23), .A1(n961), .B0(n54), .C0(n1445), .Y(n2426) );
  NAND2X1 U1702 ( .A(H7[21]), .B(n222), .Y(n1445) );
  OAI211X1 U1703 ( .A0(n18), .A1(n955), .B0(n55), .C0(n1446), .Y(n2432) );
  NAND2X1 U1704 ( .A(H7[15]), .B(n223), .Y(n1446) );
  OAI211X1 U1705 ( .A0(n19), .A1(n954), .B0(n56), .C0(n1447), .Y(n2433) );
  NAND2X1 U1706 ( .A(H7[14]), .B(n223), .Y(n1447) );
  OAI211X1 U1707 ( .A0(n24), .A1(n875), .B0(n56), .C0(n1568), .Y(n2588) );
  NAND2X1 U1708 ( .A(H3[18]), .B(n217), .Y(n1568) );
  OAI211X1 U1709 ( .A0(n18), .A1(n940), .B0(n56), .C0(n1453), .Y(n2447) );
  OAI211X1 U1710 ( .A0(n22), .A1(n742), .B0(n60), .C0(n1861), .Y(n2897) );
  INVX1 U1711 ( .A(n131), .Y(n742) );
  NAND2X1 U1712 ( .A(H0[30]), .B(n213), .Y(n1861) );
  OAI211X1 U1713 ( .A0(n24), .A1(n741), .B0(n62), .C0(n1862), .Y(n2898) );
  NAND2X1 U1714 ( .A(H0[29]), .B(n213), .Y(n1862) );
  OAI211X1 U1715 ( .A0(n21), .A1(n739), .B0(n60), .C0(n1863), .Y(n2900) );
  NAND2X1 U1716 ( .A(H0[27]), .B(n212), .Y(n1863) );
  OAI211X1 U1717 ( .A0(n21), .A1(n633), .B0(n57), .C0(n1864), .Y(n2902) );
  INVX1 U1718 ( .A(n135), .Y(n633) );
  NAND2X1 U1719 ( .A(H0[25]), .B(n212), .Y(n1864) );
  OAI211X1 U1720 ( .A0(n23), .A1(n736), .B0(n54), .C0(n1865), .Y(n2908) );
  INVX1 U1721 ( .A(n140), .Y(n736) );
  NAND2X1 U1722 ( .A(H0[19]), .B(n212), .Y(n1865) );
  OAI211X1 U1723 ( .A0(n23), .A1(n733), .B0(n61), .C0(n1866), .Y(n2911) );
  NAND2X1 U1724 ( .A(H0[16]), .B(n212), .Y(n1866) );
  OAI211X1 U1725 ( .A0(n23), .A1(n732), .B0(n60), .C0(n1867), .Y(n2912) );
  NAND2X1 U1726 ( .A(H0[15]), .B(n212), .Y(n1867) );
  OAI211X1 U1727 ( .A0(n22), .A1(n731), .B0(n61), .C0(n1868), .Y(n2913) );
  INVX1 U1728 ( .A(n145), .Y(n731) );
  NAND2X1 U1729 ( .A(H0[14]), .B(n212), .Y(n1868) );
  OAI211X1 U1730 ( .A0(n22), .A1(n730), .B0(n55), .C0(n1869), .Y(n2914) );
  NAND2X1 U1731 ( .A(H0[13]), .B(n212), .Y(n1869) );
  OAI211X1 U1732 ( .A0(n19), .A1(n727), .B0(n56), .C0(n1870), .Y(n2917) );
  NAND2X1 U1733 ( .A(H0[10]), .B(n212), .Y(n1870) );
  OAI211X1 U1734 ( .A0(n17), .A1(n726), .B0(n55), .C0(n1871), .Y(n2918) );
  NAND2X1 U1735 ( .A(H0[9]), .B(n212), .Y(n1871) );
  OAI211X1 U1736 ( .A0(n20), .A1(n723), .B0(n56), .C0(n1872), .Y(n2921) );
  INVX1 U1737 ( .A(n153), .Y(n723) );
  NAND2X1 U1738 ( .A(H0[6]), .B(n212), .Y(n1872) );
  OAI211X1 U1739 ( .A0(n20), .A1(n707), .B0(n57), .C0(n1874), .Y(n2925) );
  NAND2X1 U1740 ( .A(H0[2]), .B(n212), .Y(n1874) );
  OAI211X1 U1741 ( .A0(n23), .A1(n720), .B0(n54), .C0(n1876), .Y(n2927) );
  NAND2X1 U1742 ( .A(H0[0]), .B(n217), .Y(n1876) );
  INVXL U1743 ( .A(next_E[19]), .Y(n484) );
  OAI211X1 U1744 ( .A0(n284), .A1(n46), .B0(n486), .C0(n485), .Y(n2716) );
  OAI211X1 U1745 ( .A0(n286), .A1(n489), .B0(n488), .C0(n487), .Y(n2717) );
  INVXL U1746 ( .A(next_E[17]), .Y(n489) );
  NAND2X1 U1747 ( .A(N940), .B(n199), .Y(n487) );
  OAI211X1 U1748 ( .A0(n283), .A1(n496), .B0(n495), .C0(n494), .Y(n2720) );
  INVXL U1749 ( .A(next_E[14]), .Y(n496) );
  XOR3X2 U1750 ( .A(SHA256_result[109]), .B(n63), .C(SHA256_result[114]), .Y(
        f4_E_32[7]) );
  XOR3X2 U1751 ( .A(SHA256_result[116]), .B(SHA256_result[103]), .C(
        SHA256_result[121]), .Y(f4_E_32[14]) );
  OAI21XL U1752 ( .A0(n162), .A1(n912), .B0(n1611), .Y(n2672) );
  OAI21XL U1753 ( .A0(n744), .A1(n969), .B0(n1460), .Y(n2450) );
  AOI22X1 U1754 ( .A0(N1048), .A1(n203), .B0(SHA256_result[61]), .B1(n275), 
        .Y(n1460) );
  XOR3X2 U1755 ( .A(SHA256_result[114]), .B(SHA256_result[101]), .C(
        SHA256_result[119]), .Y(f4_E_32[12]) );
  XOR3X2 U1756 ( .A(SHA256_result[110]), .B(n67), .C(SHA256_result[115]), .Y(
        f4_E_32[8]) );
  XOR3X2 U1757 ( .A(SHA256_result[117]), .B(SHA256_result[104]), .C(
        SHA256_result[122]), .Y(f4_E_32[15]) );
  XOR3X2 U1758 ( .A(SHA256_result[115]), .B(SHA256_result[102]), .C(
        SHA256_result[120]), .Y(f4_E_32[13]) );
  XOR3X2 U1759 ( .A(SHA256_result[112]), .B(SHA256_result[99]), .C(
        SHA256_result[117]), .Y(f4_E_32[10]) );
  XOR3X2 U1760 ( .A(SHA256_result[111]), .B(SHA256_result[98]), .C(
        SHA256_result[116]), .Y(f4_E_32[9]) );
  OAI2BB2X1 U1761 ( .B0(n342), .B1(n898), .A0N(H4[22]), .A1N(n227), .Y(n2616)
         );
  OAI2BB2X1 U1762 ( .B0(n342), .B1(n889), .A0N(H4[13]), .A1N(n224), .Y(n2625)
         );
  OAI2BB2X1 U1763 ( .B0(n342), .B1(n743), .A0N(H0[31]), .A1N(n210), .Y(n2896)
         );
  OAI2BB2X1 U1764 ( .B0(n342), .B1(n740), .A0N(H0[28]), .A1N(n219), .Y(n2899)
         );
  OAI2BB2X1 U1765 ( .B0(n342), .B1(n892), .A0N(H4[16]), .A1N(n218), .Y(n2622)
         );
  OAI2BB2X1 U1766 ( .B0(n342), .B1(n910), .A0N(H5[22]), .A1N(n227), .Y(n2648)
         );
  OAI2BB2X1 U1767 ( .B0(n342), .B1(n909), .A0N(H5[21]), .A1N(n227), .Y(n2649)
         );
  OAI2BB2X1 U1768 ( .B0(n342), .B1(n908), .A0N(H5[20]), .A1N(n227), .Y(n2650)
         );
  OAI2BB2X1 U1769 ( .B0(n342), .B1(n907), .A0N(H5[19]), .A1N(n227), .Y(n2651)
         );
  OAI2BB2X1 U1770 ( .B0(n342), .B1(n912), .A0N(H5[30]), .A1N(n225), .Y(n2640)
         );
  OAI2BB2X1 U1771 ( .B0(n342), .B1(n899), .A0N(H4[23]), .A1N(n227), .Y(n2615)
         );
  OAI2BB2X1 U1772 ( .B0(n342), .B1(n78), .A0N(H1[1]), .A1N(n223), .Y(n2862) );
  OAI2BB2X1 U1773 ( .B0(n342), .B1(n823), .A0N(H1[26]), .A1N(n226), .Y(n2837)
         );
  OAI2BB2X1 U1774 ( .B0(n342), .B1(n816), .A0N(H1[19]), .A1N(n225), .Y(n2844)
         );
  OAI2BB2X1 U1775 ( .B0(n342), .B1(n811), .A0N(H1[14]), .A1N(n225), .Y(n2849)
         );
  OAI2BB2X1 U1776 ( .B0(n342), .B1(n809), .A0N(H1[12]), .A1N(n225), .Y(n2851)
         );
  OAI2BB2X1 U1777 ( .B0(n342), .B1(n855), .A0N(H2[31]), .A1N(n224), .Y(n2544)
         );
  OAI2BB2X1 U1778 ( .B0(n342), .B1(n848), .A0N(H2[24]), .A1N(n224), .Y(n2551)
         );
  OAI2BB2X1 U1779 ( .B0(n342), .B1(n840), .A0N(H2[16]), .A1N(n224), .Y(n2559)
         );
  OAI2BB2X1 U1780 ( .B0(n342), .B1(n834), .A0N(H2[10]), .A1N(n224), .Y(n2565)
         );
  OAI2BB2X1 U1781 ( .B0(n342), .B1(n929), .A0N(H6[22]), .A1N(n227), .Y(n2520)
         );
  OAI2BB2X1 U1782 ( .B0(n342), .B1(n928), .A0N(H6[21]), .A1N(n226), .Y(n2521)
         );
  OAI2BB2X1 U1783 ( .B0(n342), .B1(n937), .A0N(H6[30]), .A1N(n226), .Y(n2512)
         );
  OAI2BB2X1 U1784 ( .B0(n342), .B1(n897), .A0N(H4[21]), .A1N(n227), .Y(n2617)
         );
  OAI2BB2X1 U1785 ( .B0(n342), .B1(n896), .A0N(H4[20]), .A1N(n214), .Y(n2618)
         );
  OAI2BB2X1 U1786 ( .B0(n342), .B1(n891), .A0N(H4[15]), .A1N(n215), .Y(n2623)
         );
  OAI2BB2X1 U1787 ( .B0(n342), .B1(n1145), .A0N(H5[23]), .A1N(n227), .Y(n2647)
         );
  OAI2BB2X1 U1788 ( .B0(n342), .B1(n1151), .A0N(H5[17]), .A1N(n227), .Y(n2653)
         );
  OAI2BB2X1 U1789 ( .B0(n342), .B1(n1142), .A0N(H5[26]), .A1N(n227), .Y(n2644)
         );
  OAI21XL U1790 ( .A0(n342), .A1(n550), .B0(n549), .Y(n2607) );
  NAND2X1 U1791 ( .A(H4[31]), .B(n220), .Y(n549) );
  OAI2BB2X1 U1792 ( .B0(n342), .B1(n827), .A0N(H1[30]), .A1N(n226), .Y(n2833)
         );
  OAI2BB2X1 U1793 ( .B0(n342), .B1(n820), .A0N(H1[23]), .A1N(n225), .Y(n2840)
         );
  OAI2BB2X1 U1794 ( .B0(n342), .B1(n817), .A0N(H1[20]), .A1N(n225), .Y(n2843)
         );
  XOR3X2 U1795 ( .A(SHA256_result[127]), .B(SHA256_result[108]), .C(
        SHA256_result[113]), .Y(f4_E_32[6]) );
  OAI2BB2X1 U1796 ( .B0(n342), .B1(n885), .A0N(H3[28]), .A1N(n223), .Y(n2578)
         );
  OAI2BB2X1 U1797 ( .B0(n342), .B1(n884), .A0N(H3[27]), .A1N(n221), .Y(n2579)
         );
  OAI2BB2X1 U1798 ( .B0(n342), .B1(n854), .A0N(H2[30]), .A1N(n224), .Y(n2545)
         );
  OAI2BB2X1 U1799 ( .B0(n342), .B1(n849), .A0N(H2[25]), .A1N(n224), .Y(n2550)
         );
  OAI2BB2X1 U1800 ( .B0(n342), .B1(n847), .A0N(H2[23]), .A1N(n224), .Y(n2552)
         );
  OAI2BB2X1 U1801 ( .B0(n342), .B1(n844), .A0N(H2[20]), .A1N(n225), .Y(n2555)
         );
  OAI2BB2X1 U1802 ( .B0(n342), .B1(n835), .A0N(H2[11]), .A1N(n224), .Y(n2564)
         );
  OAI2BB2X1 U1803 ( .B0(n342), .B1(n831), .A0N(H2[7]), .A1N(n224), .Y(n2568)
         );
  OAI2BB2X1 U1804 ( .B0(n342), .B1(n877), .A0N(H3[20]), .A1N(n222), .Y(n2586)
         );
  OAI2BB2X1 U1805 ( .B0(n342), .B1(n878), .A0N(H3[21]), .A1N(n217), .Y(n2585)
         );
  OAI2BB2X1 U1806 ( .B0(n342), .B1(n927), .A0N(H6[20]), .A1N(n226), .Y(n2522)
         );
  OAI2BB2X1 U1807 ( .B0(n342), .B1(n926), .A0N(H6[19]), .A1N(n225), .Y(n2523)
         );
  OAI2BB2X1 U1808 ( .B0(n342), .B1(n925), .A0N(H6[18]), .A1N(n225), .Y(n2524)
         );
  OAI2BB2X1 U1809 ( .B0(n342), .B1(n920), .A0N(H6[13]), .A1N(n225), .Y(n2529)
         );
  OAI2BB2X1 U1810 ( .B0(n342), .B1(n938), .A0N(H6[31]), .A1N(n212), .Y(n2511)
         );
  OAI2BB2X1 U1811 ( .B0(n342), .B1(n936), .A0N(H6[29]), .A1N(n222), .Y(n2513)
         );
  OAI2BB2X1 U1812 ( .B0(n342), .B1(n887), .A0N(H3[30]), .A1N(n224), .Y(n2576)
         );
  OAI2BB2X1 U1813 ( .B0(n342), .B1(n859), .A0N(H3[2]), .A1N(n226), .Y(n2604)
         );
  OAI2BB2X1 U1814 ( .B0(n342), .B1(n911), .A0N(H5[29]), .A1N(n227), .Y(n2641)
         );
  OAI2BB2X1 U1815 ( .B0(n342), .B1(n966), .A0N(H7[26]), .A1N(n225), .Y(n2421)
         );
  OAI2BB2X1 U1816 ( .B0(n342), .B1(n942), .A0N(H7[2]), .A1N(n226), .Y(n2445)
         );
  OAI2BB2X1 U1817 ( .B0(n342), .B1(n882), .A0N(H3[25]), .A1N(n210), .Y(n2581)
         );
  OAI2BB2X1 U1818 ( .B0(n342), .B1(n880), .A0N(H3[23]), .A1N(n224), .Y(n2583)
         );
  OAI2BB2X1 U1819 ( .B0(n342), .B1(n960), .A0N(H7[20]), .A1N(n226), .Y(n2427)
         );
  OAI2BB2X1 U1820 ( .B0(n342), .B1(n959), .A0N(H7[19]), .A1N(n226), .Y(n2428)
         );
  OAI2BB2X1 U1821 ( .B0(n342), .B1(n958), .A0N(H7[18]), .A1N(n226), .Y(n2429)
         );
  OAI2BB2X1 U1822 ( .B0(n342), .B1(n957), .A0N(H7[17]), .A1N(n226), .Y(n2430)
         );
  OAI2BB2X1 U1823 ( .B0(n342), .B1(n956), .A0N(H7[16]), .A1N(n226), .Y(n2431)
         );
  OAI2BB2X1 U1824 ( .B0(n342), .B1(n953), .A0N(H7[13]), .A1N(n227), .Y(n2434)
         );
  OAI2BB2X1 U1825 ( .B0(n342), .B1(n952), .A0N(H7[12]), .A1N(n227), .Y(n2435)
         );
  OAI2BB2X1 U1826 ( .B0(n342), .B1(n939), .A0N(H7[31]), .A1N(n225), .Y(n2416)
         );
  OAI2BB2X1 U1827 ( .B0(n342), .B1(n969), .A0N(H7[29]), .A1N(n225), .Y(n2418)
         );
  OAI21XL U1828 ( .A0(n342), .A1(n464), .B0(n463), .Y(n2612) );
  NAND2X1 U1829 ( .A(H4[26]), .B(n220), .Y(n463) );
  OAI21XL U1830 ( .A0(n342), .A1(n460), .B0(n459), .Y(n2611) );
  NAND2X1 U1831 ( .A(H4[27]), .B(n219), .Y(n459) );
  OAI21XL U1832 ( .A0(n342), .A1(n468), .B0(n467), .Y(n2613) );
  NAND2X1 U1833 ( .A(H4[25]), .B(n220), .Y(n467) );
  OAI21XL U1834 ( .A0(n342), .A1(n520), .B0(n519), .Y(n2631) );
  NAND2X1 U1835 ( .A(H4[7]), .B(n220), .Y(n519) );
  OAI21XL U1836 ( .A0(n342), .A1(n502), .B0(n501), .Y(n2627) );
  NAND2X1 U1837 ( .A(H4[11]), .B(n220), .Y(n501) );
  OAI21XL U1838 ( .A0(n342), .A1(n646), .B0(n645), .Y(n2905) );
  NAND2X1 U1839 ( .A(H0[22]), .B(n221), .Y(n645) );
  OAI2BB2X1 U1840 ( .B0(n342), .B1(n728), .A0N(H0[11]), .A1N(n224), .Y(n2916)
         );
  OAI2BB2X1 U1841 ( .B0(n342), .B1(n724), .A0N(H0[7]), .A1N(n224), .Y(n2920)
         );
  OAI2BB2X1 U1842 ( .B0(n342), .B1(n734), .A0N(H0[17]), .A1N(n224), .Y(n2910)
         );
  INVX1 U1843 ( .A(n139), .Y(n737) );
  OAI2BB2X1 U1844 ( .B0(n342), .B1(n729), .A0N(H0[12]), .A1N(n224), .Y(n2915)
         );
  INVX1 U1845 ( .A(n147), .Y(n729) );
  OAI2BB2X1 U1846 ( .B0(n342), .B1(n725), .A0N(H0[8]), .A1N(n224), .Y(n2919)
         );
  INVX1 U1847 ( .A(n151), .Y(n725) );
  OAI21XL U1848 ( .A0(n342), .A1(n443), .B0(n406), .Y(n2538) );
  OAI21XL U1849 ( .A0(n342), .A1(n515), .B0(n514), .Y(n2630) );
  NAND2X1 U1850 ( .A(H4[8]), .B(n220), .Y(n514) );
  OAI21XL U1851 ( .A0(n342), .A1(n506), .B0(n505), .Y(n2628) );
  NAND2X1 U1852 ( .A(H4[10]), .B(n220), .Y(n505) );
  OAI21XL U1853 ( .A0(n165), .A1(n885), .B0(n1694), .Y(n2738) );
  AOI22X1 U1854 ( .A0(N919), .A1(n199), .B0(SHA256_result[188]), .B1(n271), 
        .Y(n1694) );
  XOR3X2 U1855 ( .A(SHA256_result[113]), .B(SHA256_result[100]), .C(
        SHA256_result[118]), .Y(f4_E_32[11]) );
  OAI21XL U1856 ( .A0(n342), .A1(n446), .B0(n411), .Y(n2540) );
  OAI21XL U1857 ( .A0(n342), .A1(n558), .B0(n557), .Y(n2572) );
  OAI21XL U1858 ( .A0(n342), .A1(n630), .B0(n629), .Y(n2901) );
  NAND2X1 U1859 ( .A(H0[26]), .B(n221), .Y(n629) );
  OAI21XL U1860 ( .A0(n342), .A1(n642), .B0(n641), .Y(n2904) );
  NAND2X1 U1861 ( .A(H0[23]), .B(n221), .Y(n641) );
  OAI21XL U1862 ( .A0(n342), .A1(n638), .B0(n637), .Y(n2903) );
  NAND2X1 U1863 ( .A(H0[24]), .B(n221), .Y(n637) );
  OAI21XL U1864 ( .A0(n342), .A1(n697), .B0(n696), .Y(n2923) );
  NAND2X1 U1865 ( .A(H0[4]), .B(n221), .Y(n696) );
  OAI21XL U1866 ( .A0(n342), .A1(n702), .B0(n701), .Y(n2924) );
  NAND2X1 U1867 ( .A(H0[3]), .B(n222), .Y(n701) );
  OAI21XL U1868 ( .A0(n342), .A1(n571), .B0(n570), .Y(n2799) );
  OAI21XL U1869 ( .A0(n342), .A1(n562), .B0(n561), .Y(n2573) );
  NAND3BX1 U1870 ( .AN(n420), .B(n419), .C(n418), .Y(n2674) );
  OAI21XL U1871 ( .A0(n1140), .A1(n175), .B0(n677), .Y(n420) );
  NAND2X1 U1872 ( .A(N983), .B(n195), .Y(n418) );
  AOI21X1 U1873 ( .A0(SHA256_result[126]), .A1(n180), .B0(n128), .Y(n450) );
  NAND2XL U1874 ( .A(n44), .B(n335), .Y(n449) );
  NAND2X1 U1875 ( .A(H0[5]), .B(n212), .Y(n1873) );
  INVX1 U1876 ( .A(n154), .Y(n692) );
  NAND2X1 U1877 ( .A(H0[1]), .B(n212), .Y(n1875) );
  NOR2X1 U1878 ( .A(n24), .B(n92), .Y(n711) );
  NAND2XL U1879 ( .A(next_E[28]), .B(n276), .Y(n457) );
  NAND3X1 U1880 ( .A(n473), .B(n472), .C(n471), .Y(n2710) );
  NAND2XL U1881 ( .A(next_E[24]), .B(n276), .Y(n472) );
  NAND2X1 U1882 ( .A(N947), .B(n199), .Y(n471) );
  AOI2BB2X1 U1883 ( .B0(n168), .B1(SHA256_result[111]), .A0N(n316), .A1N(n492), 
        .Y(n493) );
  INVXL U1884 ( .A(next_E[15]), .Y(n492) );
  OAI2BB1X1 U1885 ( .A0N(N944), .A1N(n205), .B0(n479), .Y(n2713) );
  INVXL U1886 ( .A(next_E[21]), .Y(n478) );
  OAI2BB1X1 U1887 ( .A0N(N943), .A1N(n721), .B0(n481), .Y(n2714) );
  INVXL U1888 ( .A(next_E[20]), .Y(n480) );
  OAI2BB1X1 U1889 ( .A0N(N939), .A1N(n206), .B0(n491), .Y(n2718) );
  INVXL U1890 ( .A(next_E[16]), .Y(n490) );
  OAI2BB1X1 U1891 ( .A0N(n90), .A1N(SHA256_result[224]), .B0(n615), .Y(
        f2_ABC_32[0]) );
  OAI21XL U1892 ( .A0(SHA256_result[224]), .A1(n90), .B0(SHA256_result[160]), 
        .Y(n615) );
  OAI221XL U1893 ( .A0(n303), .A1(n900), .B0(n194), .B1(n1144), .C0(n1617), 
        .Y(n2678) );
  OAI221XL U1894 ( .A0(n302), .A1(n892), .B0(n178), .B1(n1152), .C0(n1625), 
        .Y(n2686) );
  OAI221XL U1895 ( .A0(n302), .A1(n890), .B0(n178), .B1(n1154), .C0(n1627), 
        .Y(n2688) );
  OAI221XL U1896 ( .A0(n307), .A1(n1140), .B0(n193), .B1(n935), .C0(n1496), 
        .Y(n2483) );
  OAI221XL U1897 ( .A0(n306), .A1(n1141), .B0(n191), .B1(n934), .C0(n1497), 
        .Y(n2484) );
  OAI221XL U1898 ( .A0(n306), .A1(n1143), .B0(n190), .B1(n932), .C0(n1499), 
        .Y(n2486) );
  OAI221XL U1899 ( .A0(n305), .A1(n1144), .B0(n192), .B1(n931), .C0(n1500), 
        .Y(n2487) );
  OAI221XL U1900 ( .A0(n305), .A1(n1145), .B0(n194), .B1(n930), .C0(n1501), 
        .Y(n2488) );
  OAI221XL U1901 ( .A0(n306), .A1(n1142), .B0(n194), .B1(n933), .C0(n1498), 
        .Y(n2485) );
  OAI221XL U1902 ( .A0(n305), .A1(n1151), .B0(n193), .B1(n924), .C0(n1507), 
        .Y(n2494) );
  AOI21X1 U1903 ( .A0(N1004), .A1(n199), .B0(n258), .Y(n1507) );
  OAI221XL U1904 ( .A0(n304), .A1(n1152), .B0(n190), .B1(n923), .C0(n1508), 
        .Y(n2495) );
  AOI21X1 U1905 ( .A0(N1003), .A1(n200), .B0(n258), .Y(n1508) );
  OAI221XL U1906 ( .A0(n303), .A1(n1161), .B0(n194), .B1(n914), .C0(n1517), 
        .Y(n2504) );
  NAND2XL U1907 ( .A(SHA256_result[34]), .B(n170), .Y(n413) );
  NAND2X1 U1908 ( .A(N989), .B(n198), .Y(n412) );
  OAI211X1 U1909 ( .A0(n78), .A1(n321), .B0(n567), .C0(n566), .Y(n2797) );
  OAI211X1 U1910 ( .A0(n284), .A1(n531), .B0(n433), .C0(n432), .Y(n2698) );
  OAI211X1 U1911 ( .A0(n285), .A1(n72), .B0(n437), .C0(n436), .Y(n2700) );
  NAND2X1 U1912 ( .A(N957), .B(n204), .Y(n437) );
  AOI21XL U1913 ( .A0(SHA256_result[66]), .A1(n180), .B0(n260), .Y(n436) );
  OAI211X1 U1914 ( .A0(n1163), .A1(n320), .B0(n405), .C0(n404), .Y(n2506) );
  NAND2X1 U1915 ( .A(N992), .B(n200), .Y(n405) );
  OAI211X1 U1916 ( .A0(n1167), .A1(n321), .B0(n415), .C0(n414), .Y(n2510) );
  OAI211X1 U1917 ( .A0(n1165), .A1(n322), .B0(n410), .C0(n409), .Y(n2508) );
  AOI21XL U1918 ( .A0(SHA256_result[35]), .A1(n179), .B0(n261), .Y(n409) );
  OAI211X1 U1919 ( .A0(n288), .A1(n509), .B0(n508), .C0(n507), .Y(n2724) );
  INVX1 U1920 ( .A(next_E[10]), .Y(n509) );
  NAND2X1 U1921 ( .A(SHA256_result[106]), .B(n170), .Y(n508) );
  NAND2X1 U1922 ( .A(N933), .B(n203), .Y(n507) );
  OAI211X1 U1923 ( .A0(n285), .A1(n513), .B0(n512), .C0(n511), .Y(n2725) );
  NAND2X1 U1924 ( .A(N932), .B(n204), .Y(n512) );
  AOI21XL U1925 ( .A0(SHA256_result[105]), .A1(n181), .B0(n128), .Y(n511) );
  OAI211X1 U1926 ( .A0(n288), .A1(n518), .B0(n517), .C0(n516), .Y(n2726) );
  NAND2XL U1927 ( .A(SHA256_result[104]), .B(n168), .Y(n517) );
  NAND2X1 U1928 ( .A(N931), .B(n206), .Y(n516) );
  OAI211X1 U1929 ( .A0(n284), .A1(n523), .B0(n522), .C0(n521), .Y(n2727) );
  NAND2XL U1930 ( .A(SHA256_result[103]), .B(n171), .Y(n522) );
  NAND2X1 U1931 ( .A(N930), .B(n721), .Y(n521) );
  OAI211X1 U1932 ( .A0(n289), .A1(n527), .B0(n526), .C0(n525), .Y(n2728) );
  NAND2X1 U1933 ( .A(N929), .B(n717), .Y(n526) );
  AOI21XL U1934 ( .A0(SHA256_result[102]), .A1(n181), .B0(n260), .Y(n525) );
  OAI211X1 U1935 ( .A0(n282), .A1(n530), .B0(n529), .C0(n528), .Y(n2729) );
  OAI211X1 U1936 ( .A0(n290), .A1(n534), .B0(n533), .C0(n532), .Y(n2730) );
  NAND2X1 U1937 ( .A(N927), .B(n196), .Y(n533) );
  OAI211X1 U1938 ( .A0(n286), .A1(n538), .B0(n537), .C0(n536), .Y(n2731) );
  INVX1 U1939 ( .A(next_E[3]), .Y(n538) );
  NAND2X1 U1940 ( .A(N926), .B(n204), .Y(n537) );
  AOI21XL U1941 ( .A0(SHA256_result[99]), .A1(n184), .B0(n128), .Y(n536) );
  OAI211X1 U1942 ( .A0(n290), .A1(n541), .B0(n540), .C0(n539), .Y(n2732) );
  NAND2X1 U1943 ( .A(N925), .B(n200), .Y(n540) );
  AOI21XL U1944 ( .A0(SHA256_result[98]), .A1(n180), .B0(n257), .Y(n539) );
  OAI211X1 U1945 ( .A0(n285), .A1(n545), .B0(n544), .C0(n543), .Y(n2733) );
  NAND2X1 U1946 ( .A(N924), .B(n198), .Y(n544) );
  AOI21XL U1947 ( .A0(n67), .A1(n181), .B0(n128), .Y(n543) );
  OAI211X1 U1948 ( .A0(n290), .A1(n548), .B0(n547), .C0(n546), .Y(n2734) );
  INVX1 U1949 ( .A(next_E[0]), .Y(n548) );
  NAND2X1 U1950 ( .A(N923), .B(n197), .Y(n547) );
  AOI21XL U1951 ( .A0(n63), .A1(n180), .B0(n258), .Y(n546) );
  OAI211X1 U1952 ( .A0(n287), .A1(n800), .B0(n560), .C0(n559), .Y(n2795) );
  OAI211X1 U1953 ( .A0(n291), .A1(n799), .B0(n564), .C0(n563), .Y(n2796) );
  OAI211X1 U1954 ( .A0(n291), .A1(n88), .B0(n569), .C0(n568), .Y(n2798) );
  NAND2X1 U1955 ( .A(N859), .B(n204), .Y(n568) );
  OAI21XL U1956 ( .A0(n162), .A1(n928), .B0(n1503), .Y(n2490) );
  OAI21XL U1957 ( .A0(n162), .A1(n927), .B0(n1504), .Y(n2491) );
  OAI21XL U1958 ( .A0(n163), .A1(n926), .B0(n1505), .Y(n2492) );
  OAI21XL U1959 ( .A0(n163), .A1(n925), .B0(n1506), .Y(n2493) );
  OAI21XL U1960 ( .A0(n163), .A1(n920), .B0(n1511), .Y(n2498) );
  OAI21XL U1961 ( .A0(n163), .A1(n917), .B0(n1514), .Y(n2501) );
  OAI21XL U1962 ( .A0(n163), .A1(n916), .B0(n1515), .Y(n2502) );
  OAI21XL U1963 ( .A0(n163), .A1(n913), .B0(n1518), .Y(n2505) );
  OAI21XL U1964 ( .A0(n162), .A1(n1142), .B0(n1615), .Y(n2676) );
  AOI22X1 U1965 ( .A0(N981), .A1(n203), .B0(SHA256_result[122]), .B1(n273), 
        .Y(n1615) );
  OAI21XL U1966 ( .A0(n162), .A1(n1145), .B0(n1618), .Y(n2679) );
  OAI21XL U1967 ( .A0(n162), .A1(n910), .B0(n1619), .Y(n2680) );
  OAI21XL U1968 ( .A0(n744), .A1(n966), .B0(n1463), .Y(n2453) );
  AOI22X1 U1969 ( .A0(N1045), .A1(n204), .B0(SHA256_result[58]), .B1(n275), 
        .Y(n1463) );
  OAI21XL U1970 ( .A0(n744), .A1(n960), .B0(n1469), .Y(n2459) );
  OAI21XL U1971 ( .A0(n744), .A1(n959), .B0(n1470), .Y(n2460) );
  OAI21XL U1972 ( .A0(n744), .A1(n958), .B0(n1471), .Y(n2461) );
  OAI21XL U1973 ( .A0(n744), .A1(n957), .B0(n1472), .Y(n2462) );
  OAI2BB1X1 U1974 ( .A0N(SHA256_result[199]), .A1N(n152), .B0(n608), .Y(
        f2_ABC_32[7]) );
  OAI21XL U1975 ( .A0(SHA256_result[199]), .A1(n152), .B0(SHA256_result[167]), 
        .Y(n608) );
  OAI2BB1X1 U1976 ( .A0N(SHA256_result[201]), .A1N(n150), .B0(n606), .Y(
        f2_ABC_32[9]) );
  OAI2BB1X1 U1977 ( .A0N(SHA256_result[198]), .A1N(n153), .B0(n609), .Y(
        f2_ABC_32[6]) );
  OAI21XL U1978 ( .A0(SHA256_result[198]), .A1(n153), .B0(SHA256_result[166]), 
        .Y(n609) );
  OAI2BB1X1 U1979 ( .A0N(SHA256_result[203]), .A1N(n148), .B0(n604), .Y(
        f2_ABC_32[11]) );
  OAI21XL U1980 ( .A0(SHA256_result[203]), .A1(n148), .B0(SHA256_result[171]), 
        .Y(n604) );
  OAI2BB1X1 U1981 ( .A0N(SHA256_result[197]), .A1N(n154), .B0(n610), .Y(
        f2_ABC_32[5]) );
  OAI21XL U1982 ( .A0(SHA256_result[197]), .A1(n154), .B0(SHA256_result[165]), 
        .Y(n610) );
  OAI21XL U1983 ( .A0(SHA256_result[200]), .A1(n151), .B0(SHA256_result[168]), 
        .Y(n607) );
  OAI21XL U1984 ( .A0(SHA256_result[196]), .A1(n155), .B0(SHA256_result[164]), 
        .Y(n611) );
  OAI2BB1X1 U1985 ( .A0N(SHA256_result[202]), .A1N(n149), .B0(n605), .Y(
        f2_ABC_32[10]) );
  NAND2BX1 U1986 ( .AN(n428), .B(n427), .Y(n2691) );
  OAI21XL U1987 ( .A0(n1157), .A1(n175), .B0(n677), .Y(n428) );
  XOR3X2 U1988 ( .A(SHA256_result[110]), .B(n63), .C(SHA256_result[123]), .Y(
        f4_E_32[21]) );
  XOR3X2 U1989 ( .A(SHA256_result[111]), .B(n67), .C(SHA256_result[124]), .Y(
        f4_E_32[22]) );
  XOR3X2 U1990 ( .A(SHA256_result[121]), .B(SHA256_result[108]), .C(
        SHA256_result[126]), .Y(f4_E_32[19]) );
  XOR3X2 U1991 ( .A(SHA256_result[118]), .B(SHA256_result[105]), .C(
        SHA256_result[123]), .Y(f4_E_32[16]) );
  XOR3X2 U1992 ( .A(SHA256_result[119]), .B(SHA256_result[106]), .C(
        SHA256_result[124]), .Y(f4_E_32[17]) );
  XOR3X2 U1993 ( .A(SHA256_result[246]), .B(n148), .C(n25), .Y(f3_A_32[9]) );
  MX2X1 U1994 ( .A(SHA256_result[53]), .B(SHA256_result[85]), .S0(
        SHA256_result[117]), .Y(f1_EFG_32[21]) );
  MX2X1 U1995 ( .A(SHA256_result[50]), .B(SHA256_result[82]), .S0(
        SHA256_result[114]), .Y(f1_EFG_32[18]) );
  XOR3X2 U1996 ( .A(SHA256_result[106]), .B(SHA256_result[101]), .C(
        SHA256_result[120]), .Y(f4_E_32[31]) );
  OAI21XL U1997 ( .A0(n162), .A1(n909), .B0(n1620), .Y(n2681) );
  OAI21XL U1998 ( .A0(n164), .A1(n908), .B0(n1621), .Y(n2682) );
  OAI21XL U1999 ( .A0(n164), .A1(n907), .B0(n1622), .Y(n2683) );
  OAI21XL U2000 ( .A0(n164), .A1(n904), .B0(n1631), .Y(n2692) );
  AOI22X1 U2001 ( .A0(N965), .A1(n206), .B0(SHA256_result[106]), .B1(n272), 
        .Y(n1631) );
  OAI21XL U2002 ( .A0(n163), .A1(n903), .B0(n1632), .Y(n2693) );
  AOI22XL U2003 ( .A0(N964), .A1(n199), .B0(SHA256_result[105]), .B1(n272), 
        .Y(n1632) );
  OAI21XL U2004 ( .A0(n163), .A1(n902), .B0(n1635), .Y(n2696) );
  OAI21XL U2006 ( .A0(n163), .A1(n1163), .B0(n1636), .Y(n2697) );
  OAI21XL U2007 ( .A0(n163), .A1(n1167), .B0(n1640), .Y(n2701) );
  AOI22XL U2008 ( .A0(N956), .A1(n205), .B0(n67), .B1(n272), .Y(n1640) );
  OAI21XL U2009 ( .A0(n164), .A1(n1151), .B0(n1624), .Y(n2685) );
  OAI21XL U2010 ( .A0(n164), .A1(n1156), .B0(n1629), .Y(n2690) );
  AOI22XL U2011 ( .A0(N967), .A1(n202), .B0(SHA256_result[108]), .B1(n272), 
        .Y(n1629) );
  OAI21XL U2012 ( .A0(n165), .A1(n1168), .B0(n1641), .Y(n2702) );
  OAI21XL U2013 ( .A0(n165), .A1(n848), .B0(n1730), .Y(n2774) );
  AOI22X1 U2014 ( .A0(N883), .A1(n197), .B0(SHA256_result[216]), .B1(n270), 
        .Y(n1730) );
  OAI21XL U2015 ( .A0(n162), .A1(n840), .B0(n1738), .Y(n2782) );
  OAI21XL U2016 ( .A0(n165), .A1(n834), .B0(n1744), .Y(n2788) );
  OAI21XL U2017 ( .A0(n162), .A1(n929), .B0(n1502), .Y(n2489) );
  OAI21XL U2018 ( .A0(n162), .A1(n884), .B0(n1695), .Y(n2739) );
  AOI22X1 U2019 ( .A0(N918), .A1(n197), .B0(SHA256_result[187]), .B1(n271), 
        .Y(n1695) );
  OAI21XL U2020 ( .A0(n165), .A1(n849), .B0(n1729), .Y(n2773) );
  AOI22X1 U2021 ( .A0(N884), .A1(n201), .B0(SHA256_result[217]), .B1(n270), 
        .Y(n1729) );
  OAI21XL U2022 ( .A0(n165), .A1(n847), .B0(n1731), .Y(n2775) );
  OAI21XL U2023 ( .A0(n162), .A1(n844), .B0(n1734), .Y(n2778) );
  OAI21XL U2024 ( .A0(n165), .A1(n835), .B0(n1743), .Y(n2787) );
  AOI22X1 U2025 ( .A0(N870), .A1(n197), .B0(SHA256_result[203]), .B1(n270), 
        .Y(n1743) );
  OAI21XL U2026 ( .A0(n165), .A1(n831), .B0(n1747), .Y(n2791) );
  OAI21XL U2027 ( .A0(n164), .A1(n877), .B0(n1702), .Y(n2746) );
  OAI21XL U2028 ( .A0(n162), .A1(n878), .B0(n1701), .Y(n2745) );
  OAI21XL U2029 ( .A0(n164), .A1(n868), .B0(n1711), .Y(n2755) );
  OAI21XL U2030 ( .A0(n164), .A1(n866), .B0(n1713), .Y(n2757) );
  OAI21XL U2031 ( .A0(n164), .A1(n864), .B0(n1715), .Y(n2759) );
  OAI21XL U2032 ( .A0(n164), .A1(n863), .B0(n1716), .Y(n2760) );
  OAI21XL U2033 ( .A0(n165), .A1(n859), .B0(n1720), .Y(n2764) );
  AOI22XL U2034 ( .A0(N893), .A1(n195), .B0(SHA256_result[162]), .B1(n271), 
        .Y(n1720) );
  OAI21XL U2035 ( .A0(n165), .A1(n857), .B0(n1722), .Y(n2766) );
  OAI21XL U2036 ( .A0(n744), .A1(n949), .B0(n1480), .Y(n2470) );
  OAI21XL U2037 ( .A0(n744), .A1(n947), .B0(n1482), .Y(n2472) );
  AOI22X1 U2038 ( .A0(N1026), .A1(n196), .B0(SHA256_result[39]), .B1(n274), 
        .Y(n1482) );
  OAI21XL U2039 ( .A0(n744), .A1(n946), .B0(n1483), .Y(n2473) );
  OAI21XL U2040 ( .A0(n744), .A1(n945), .B0(n1484), .Y(n2474) );
  OAI21XL U2041 ( .A0(n744), .A1(n942), .B0(n1487), .Y(n2477) );
  AOI22XL U2042 ( .A0(N1021), .A1(n203), .B0(SHA256_result[34]), .B1(n274), 
        .Y(n1487) );
  OAI21XL U2043 ( .A0(n744), .A1(n941), .B0(n1488), .Y(n2478) );
  OAI21XL U2044 ( .A0(n165), .A1(n882), .B0(n1697), .Y(n2741) );
  AOI22X1 U2045 ( .A0(N916), .A1(n205), .B0(SHA256_result[185]), .B1(n271), 
        .Y(n1697) );
  OAI21XL U2046 ( .A0(n162), .A1(n880), .B0(n1699), .Y(n2743) );
  AOI22X1 U2047 ( .A0(N914), .A1(n206), .B0(SHA256_result[183]), .B1(n271), 
        .Y(n1699) );
  OAI21XL U2048 ( .A0(n744), .A1(n956), .B0(n1473), .Y(n2463) );
  OAI21XL U2049 ( .A0(n744), .A1(n953), .B0(n1476), .Y(n2466) );
  OAI21XL U2050 ( .A0(n744), .A1(n952), .B0(n1477), .Y(n2467) );
  NAND3BX1 U2051 ( .AN(n423), .B(n422), .C(n421), .Y(n2675) );
  OAI21XL U2052 ( .A0(n1141), .A1(n175), .B0(n677), .Y(n423) );
  NAND2X1 U2053 ( .A(N982), .B(n197), .Y(n421) );
  NAND3BX1 U2054 ( .AN(n426), .B(n425), .C(n424), .Y(n2677) );
  OAI21XL U2055 ( .A0(n1143), .A1(n175), .B0(n677), .Y(n426) );
  OAI2BB1X1 U2056 ( .A0N(N934), .A1N(n199), .B0(n504), .Y(n2723) );
  INVXL U2057 ( .A(next_E[11]), .Y(n503) );
  NAND2X1 U2058 ( .A(n500), .B(n499), .Y(n2722) );
  AOI21XL U2059 ( .A0(n183), .A1(SHA256_result[108]), .B0(n261), .Y(n499) );
  NAND2BX1 U2060 ( .AN(n430), .B(n429), .Y(n2695) );
  OAI21XL U2061 ( .A0(n1161), .A1(n175), .B0(n677), .Y(n430) );
  NAND2BX1 U2062 ( .AN(n435), .B(n434), .Y(n2699) );
  OAI21XL U2063 ( .A0(n1165), .A1(n175), .B0(n677), .Y(n435) );
  OAI2BB1X1 U2064 ( .A0N(N936), .A1N(n195), .B0(n498), .Y(n2721) );
  AOI2BB2XL U2065 ( .B0(n168), .B1(SHA256_result[109]), .A0N(n323), .A1N(n497), 
        .Y(n498) );
  INVXL U2066 ( .A(next_E[13]), .Y(n497) );
  NAND2BX1 U2067 ( .AN(n583), .B(n582), .Y(n2831) );
  OAI2BB1X1 U2068 ( .A0N(SHA256_result[206]), .A1N(n145), .B0(n601), .Y(
        f2_ABC_32[14]) );
  OAI21XL U2069 ( .A0(SHA256_result[206]), .A1(n145), .B0(SHA256_result[174]), 
        .Y(n601) );
  OAI2BB1X1 U2070 ( .A0N(SHA256_result[209]), .A1N(n142), .B0(n598), .Y(
        f2_ABC_32[17]) );
  OAI21XL U2071 ( .A0(SHA256_result[209]), .A1(n142), .B0(SHA256_result[177]), 
        .Y(n598) );
  OAI2BB1X1 U2072 ( .A0N(SHA256_result[207]), .A1N(n144), .B0(n600), .Y(
        f2_ABC_32[15]) );
  OAI21XL U2073 ( .A0(SHA256_result[207]), .A1(n144), .B0(SHA256_result[175]), 
        .Y(n600) );
  OAI2BB1X1 U2074 ( .A0N(SHA256_result[210]), .A1N(n141), .B0(n597), .Y(
        f2_ABC_32[18]) );
  OAI21XL U2075 ( .A0(SHA256_result[210]), .A1(n141), .B0(SHA256_result[178]), 
        .Y(n597) );
  OAI2BB1X1 U2076 ( .A0N(SHA256_result[204]), .A1N(n147), .B0(n603), .Y(
        f2_ABC_32[12]) );
  OAI21XL U2077 ( .A0(SHA256_result[204]), .A1(n147), .B0(SHA256_result[172]), 
        .Y(n603) );
  OAI2BB1X1 U2078 ( .A0N(SHA256_result[205]), .A1N(n146), .B0(n602), .Y(
        f2_ABC_32[13]) );
  OAI21XL U2079 ( .A0(SHA256_result[205]), .A1(n146), .B0(SHA256_result[173]), 
        .Y(n602) );
  XOR3X2 U2080 ( .A(SHA256_result[101]), .B(n63), .C(SHA256_result[115]), .Y(
        f4_E_32[26]) );
  XOR3X2 U2081 ( .A(SHA256_result[113]), .B(SHA256_result[99]), .C(
        SHA256_result[126]), .Y(f4_E_32[24]) );
  XOR3X2 U2082 ( .A(SHA256_result[127]), .B(SHA256_result[109]), .C(
        SHA256_result[122]), .Y(f4_E_32[20]) );
  XOR3X2 U2083 ( .A(n154), .B(n142), .C(SHA256_result[252]), .Y(f3_A_32[15])
         );
  MX2X1 U2084 ( .A(SHA256_result[52]), .B(SHA256_result[84]), .S0(
        SHA256_result[116]), .Y(f1_EFG_32[20]) );
  XOR3X2 U2085 ( .A(n139), .B(n151), .C(n25), .Y(f3_A_32[18]) );
  MX2X1 U2086 ( .A(SHA256_result[54]), .B(SHA256_result[86]), .S0(
        SHA256_result[118]), .Y(f1_EFG_32[22]) );
  INVX1 U2087 ( .A(n1489), .Y(n744) );
  OAI21XL U2088 ( .A0(first_block), .A1(n1490), .B0(n1491), .Y(n1489) );
  INVX1 U2089 ( .A(SHA256_result[56]), .Y(n931) );
  INVX1 U2090 ( .A(SHA256_result[57]), .Y(n932) );
  INVX1 U2091 ( .A(SHA256_result[59]), .Y(n934) );
  AOI31X1 U2092 ( .A0(n2399), .A1(n2400), .A2(n2401), .B0(n233), .Y(N2948) );
  AND3X2 U2093 ( .A(n2165), .B(n2133), .C(n785), .Y(n2400) );
  AOI211X1 U2094 ( .A0(n2248), .A1(n1388), .B0(n2402), .C0(n2116), .Y(n2401)
         );
  AOI31X1 U2095 ( .A0(n2365), .A1(n2366), .A2(n2367), .B0(n233), .Y(N2953) );
  NOR3X1 U2096 ( .A(n2224), .B(n2249), .C(n2191), .Y(n2366) );
  AOI211X1 U2097 ( .A0(n2268), .A1(n1388), .B0(n2368), .C0(n2369), .Y(n2367)
         );
  AOI31X1 U2098 ( .A0(n2278), .A1(n2279), .A2(n2280), .B0(n234), .Y(N2963) );
  AOI211X1 U2099 ( .A0(n2220), .A1(n1370), .B0(n2281), .C0(n2282), .Y(n2280)
         );
  AOI31X1 U2100 ( .A0(n2141), .A1(n2142), .A2(n2143), .B0(n234), .Y(N2975) );
  AOI31X1 U2101 ( .A0(n777), .A1(n1383), .A2(n2135), .B0(n2152), .Y(n2141) );
  NOR3BX1 U2102 ( .AN(n2149), .B(n2150), .C(n2151), .Y(n2142) );
  AOI211X1 U2103 ( .A0(n2144), .A1(n112), .B0(n2145), .C0(n767), .Y(n2143) );
  AOI31X1 U2104 ( .A0(n2058), .A1(n2059), .A2(n2060), .B0(n252), .Y(N3060) );
  AOI31X1 U2105 ( .A0(n2038), .A1(n2039), .A2(n2040), .B0(n252), .Y(N3065) );
  AOI31X1 U2106 ( .A0(n2034), .A1(n2035), .A2(n2036), .B0(n252), .Y(N3066) );
  AOI22X1 U2107 ( .A0(n241), .A1(SHA256_result[147]), .B0(n240), .B1(
        SHA256_result[179]), .Y(n2035) );
  AOI31X1 U2108 ( .A0(n2030), .A1(n2031), .A2(n2032), .B0(n252), .Y(N3067) );
  AOI22X1 U2109 ( .A0(n241), .A1(SHA256_result[148]), .B0(n240), .B1(
        SHA256_result[180]), .Y(n2031) );
  AOI31X1 U2110 ( .A0(n2062), .A1(n2063), .A2(n2064), .B0(n252), .Y(N3059) );
  AOI31X1 U2111 ( .A0(n2046), .A1(n2047), .A2(n2048), .B0(n252), .Y(N3063) );
  AOI31X1 U2112 ( .A0(n2042), .A1(n2043), .A2(n2044), .B0(n252), .Y(N3064) );
  AOI31X1 U2113 ( .A0(n2026), .A1(n2027), .A2(n2028), .B0(n252), .Y(N3068) );
  AOI22X1 U2114 ( .A0(n241), .A1(SHA256_result[149]), .B0(n240), .B1(
        SHA256_result[181]), .Y(n2027) );
  AOI31X1 U2115 ( .A0(n2022), .A1(n2023), .A2(n2024), .B0(n252), .Y(N3069) );
  AOI22X1 U2116 ( .A0(n241), .A1(SHA256_result[150]), .B0(n240), .B1(
        SHA256_result[182]), .Y(n2023) );
  AOI31X1 U2117 ( .A0(n2054), .A1(n2055), .A2(n2056), .B0(n252), .Y(N3061) );
  AOI31X1 U2118 ( .A0(n2050), .A1(n2051), .A2(n2052), .B0(n252), .Y(N3062) );
  AOI31X1 U2119 ( .A0(n2018), .A1(n2019), .A2(n2020), .B0(n252), .Y(N3070) );
  AOI22X1 U2120 ( .A0(n241), .A1(SHA256_result[151]), .B0(n240), .B1(
        SHA256_result[183]), .Y(n2019) );
  AOI31X1 U2121 ( .A0(n2014), .A1(n2015), .A2(n2016), .B0(n251), .Y(N3071) );
  AOI22X1 U2122 ( .A0(n242), .A1(SHA256_result[152]), .B0(n239), .B1(
        SHA256_result[184]), .Y(n2015) );
  AOI31X1 U2123 ( .A0(n2110), .A1(n2111), .A2(n2112), .B0(n251), .Y(N3047) );
  AOI31X1 U2124 ( .A0(n2336), .A1(n2337), .A2(n2338), .B0(n233), .Y(N2957) );
  AOI2BB2X1 U2125 ( .B0(n2137), .B1(n343), .A0N(n2146), .A1N(n769), .Y(n2336)
         );
  AOI22X1 U2126 ( .A0(n2258), .A1(n1383), .B0(n2189), .B1(n347), .Y(n2337) );
  AOI31X1 U2127 ( .A0(n2106), .A1(n2107), .A2(n2108), .B0(n251), .Y(N3048) );
  AOI211XL U2128 ( .A0(n249), .A1(n75), .B0(n352), .C0(n351), .Y(n2108) );
  AOI31X1 U2129 ( .A0(n2090), .A1(n2091), .A2(n2092), .B0(n251), .Y(N3052) );
  AOI31X1 U2130 ( .A0(n2102), .A1(n2103), .A2(n2104), .B0(n251), .Y(N3049) );
  AOI211XL U2131 ( .A0(n248), .A1(SHA256_result[34]), .B0(n354), .C0(n353), 
        .Y(n2104) );
  AOI31X1 U2132 ( .A0(n2192), .A1(n2193), .A2(n2194), .B0(n234), .Y(N2971) );
  AOI2BB2X1 U2133 ( .B0(n2176), .B1(n113), .A0N(n2184), .A1N(n346), .Y(n2192)
         );
  AOI22X1 U2134 ( .A0(n2201), .A1(n1383), .B0(n2202), .B1(n2138), .Y(n2193) );
  AOI211X1 U2135 ( .A0(n2195), .A1(n1396), .B0(n2196), .C0(n2197), .Y(n2194)
         );
  AOI31X1 U2136 ( .A0(n2086), .A1(n2087), .A2(n2088), .B0(n251), .Y(N3053) );
  AOI31X1 U2137 ( .A0(n2074), .A1(n2075), .A2(n2076), .B0(n251), .Y(N3056) );
  AOI31X1 U2138 ( .A0(n1979), .A1(n1980), .A2(n1981), .B0(n252), .Y(N3078) );
  AOI22X1 U2139 ( .A0(n242), .A1(SHA256_result[159]), .B0(n240), .B1(
        SHA256_result[191]), .Y(n1980) );
  AOI211X1 U2140 ( .A0(n248), .A1(SHA256_result[63]), .B0(n386), .C0(n385), 
        .Y(n1981) );
  AOI31X1 U2141 ( .A0(n1994), .A1(n1995), .A2(n1996), .B0(n1978), .Y(N3076) );
  AOI22X1 U2142 ( .A0(n242), .A1(SHA256_result[157]), .B0(n239), .B1(
        SHA256_result[189]), .Y(n1995) );
  AOI211X1 U2143 ( .A0(n248), .A1(SHA256_result[61]), .B0(n382), .C0(n381), 
        .Y(n1996) );
  AOI31X1 U2144 ( .A0(n2098), .A1(n2099), .A2(n2100), .B0(n251), .Y(N3050) );
  AOI211XL U2145 ( .A0(n1982), .A1(SHA256_result[35]), .B0(n356), .C0(n355), 
        .Y(n2100) );
  AOI31X1 U2146 ( .A0(n2082), .A1(n2083), .A2(n2084), .B0(n251), .Y(N3054) );
  AOI31X1 U2147 ( .A0(n2006), .A1(n2007), .A2(n2008), .B0(n1978), .Y(N3073) );
  AOI22X1 U2148 ( .A0(n242), .A1(SHA256_result[154]), .B0(n240), .B1(
        SHA256_result[186]), .Y(n2007) );
  AOI211X1 U2149 ( .A0(n248), .A1(SHA256_result[58]), .B0(n376), .C0(n375), 
        .Y(n2008) );
  AOI31X1 U2150 ( .A0(n2094), .A1(n2095), .A2(n2096), .B0(n251), .Y(N3051) );
  AOI31X1 U2151 ( .A0(n2070), .A1(n2071), .A2(n2072), .B0(n251), .Y(N3057) );
  AOI31X1 U2152 ( .A0(n1990), .A1(n1991), .A2(n1992), .B0(n1978), .Y(N3077) );
  AOI22X1 U2153 ( .A0(n242), .A1(SHA256_result[158]), .B0(n239), .B1(
        SHA256_result[190]), .Y(n1991) );
  AOI211X1 U2154 ( .A0(n248), .A1(SHA256_result[62]), .B0(n384), .C0(n383), 
        .Y(n1992) );
  AOI31X1 U2155 ( .A0(n2391), .A1(n2392), .A2(n2393), .B0(n233), .Y(N2949) );
  AOI32X1 U2156 ( .A0(n343), .A1(n1388), .A2(n2305), .B0(n112), .B1(n2398), 
        .Y(n2391) );
  AOI211X1 U2157 ( .A0(n2322), .A1(n1393), .B0(n2394), .C0(n2386), .Y(n2393)
         );
  AOI31X1 U2158 ( .A0(n2078), .A1(n2079), .A2(n2080), .B0(n251), .Y(N3055) );
  AOI31X1 U2159 ( .A0(n2066), .A1(n2067), .A2(n2068), .B0(n251), .Y(N3058) );
  AOI31X1 U2160 ( .A0(n2010), .A1(n2011), .A2(n2012), .B0(n1978), .Y(N3072) );
  AOI22X1 U2161 ( .A0(n242), .A1(SHA256_result[153]), .B0(n240), .B1(
        SHA256_result[185]), .Y(n2011) );
  AOI31X1 U2162 ( .A0(n2002), .A1(n2003), .A2(n2004), .B0(n1978), .Y(N3074) );
  AOI22X1 U2163 ( .A0(n242), .A1(SHA256_result[155]), .B0(n239), .B1(
        SHA256_result[187]), .Y(n2003) );
  AOI211X1 U2164 ( .A0(n248), .A1(SHA256_result[59]), .B0(n378), .C0(n377), 
        .Y(n2004) );
  AOI31X1 U2165 ( .A0(n1998), .A1(n1999), .A2(n2000), .B0(n1978), .Y(N3075) );
  AOI22X1 U2166 ( .A0(n242), .A1(SHA256_result[156]), .B0(n240), .B1(
        SHA256_result[188]), .Y(n1999) );
  AOI211X1 U2167 ( .A0(n248), .A1(SHA256_result[60]), .B0(n380), .C0(n379), 
        .Y(n2000) );
  AOI31X1 U2168 ( .A0(n2178), .A1(n2179), .A2(n2180), .B0(n234), .Y(N2972) );
  NOR3BX1 U2169 ( .AN(n2181), .B(n2182), .C(n2183), .Y(n2180) );
  AOI21X1 U2170 ( .A0(n2187), .A1(n159), .B0(n767), .Y(n2178) );
  AOI31X1 U2171 ( .A0(n2357), .A1(n2358), .A2(n2359), .B0(n233), .Y(N2954) );
  AOI222X1 U2172 ( .A0(n2363), .A1(n2283), .B0(n2364), .B1(n1388), .C0(n2286), 
        .C1(n41), .Y(n2358) );
  NOR4BX1 U2173 ( .AN(n772), .B(n2360), .C(n2361), .D(n2362), .Y(n2359) );
  AOI31X1 U2174 ( .A0(n2167), .A1(n2168), .A2(n2169), .B0(n234), .Y(N2973) );
  AOI222X1 U2175 ( .A0(n2175), .A1(n1383), .B0(n2124), .B1(n1370), .C0(n2176), 
        .C1(n1393), .Y(n2168) );
  NOR3X1 U2176 ( .A(n2170), .B(n2171), .C(n2172), .Y(n2169) );
  AOI31X1 U2177 ( .A0(n2227), .A1(n2228), .A2(n2229), .B0(n234), .Y(N2968) );
  AOI22X1 U2178 ( .A0(n2238), .A1(n1370), .B0(n2138), .B1(n2136), .Y(n2227) );
  NOR3X1 U2179 ( .A(n2230), .B(n2231), .C(n2171), .Y(n2229) );
  AOI211X1 U2180 ( .A0(n2139), .A1(n2235), .B0(n2236), .C0(n2237), .Y(n2228)
         );
  AOI31X1 U2181 ( .A0(n2253), .A1(n2254), .A2(n2255), .B0(n234), .Y(N2966) );
  AOI222X1 U2182 ( .A0(n2136), .A1(n756), .B0(n2232), .B1(n765), .C0(n2258), 
        .C1(n1383), .Y(n2254) );
  AND4X2 U2183 ( .A(n2256), .B(n789), .C(n2159), .D(n778), .Y(n2255) );
  INVX1 U2184 ( .A(SHA256_result[58]), .Y(n933) );
  OAI2BB1X1 U2185 ( .A0N(SHA256_result[214]), .A1N(SHA256_result[246]), .B0(
        n593), .Y(f2_ABC_32[22]) );
  OAI21XL U2186 ( .A0(SHA256_result[214]), .A1(SHA256_result[246]), .B0(
        SHA256_result[182]), .Y(n593) );
  OAI2BB1X1 U2187 ( .A0N(SHA256_result[212]), .A1N(n139), .B0(n595), .Y(
        f2_ABC_32[20]) );
  OAI21XL U2188 ( .A0(SHA256_result[212]), .A1(n139), .B0(SHA256_result[180]), 
        .Y(n595) );
  OAI2BB1X1 U2189 ( .A0N(SHA256_result[213]), .A1N(n138), .B0(n594), .Y(
        f2_ABC_32[21]) );
  OAI21XL U2190 ( .A0(SHA256_result[213]), .A1(n138), .B0(SHA256_result[181]), 
        .Y(n594) );
  OAI2BB1X1 U2191 ( .A0N(SHA256_result[211]), .A1N(n140), .B0(n596), .Y(
        f2_ABC_32[19]) );
  OAI21XL U2192 ( .A0(SHA256_result[211]), .A1(n140), .B0(SHA256_result[179]), 
        .Y(n596) );
  OAI2BB1X1 U2193 ( .A0N(SHA256_result[208]), .A1N(n143), .B0(n599), .Y(
        f2_ABC_32[16]) );
  OAI21XL U2194 ( .A0(SHA256_result[208]), .A1(n143), .B0(SHA256_result[176]), 
        .Y(n599) );
  XOR3X2 U2195 ( .A(SHA256_result[102]), .B(n67), .C(SHA256_result[116]), .Y(
        f4_E_32[27]) );
  XOR3X2 U2196 ( .A(SHA256_result[127]), .B(SHA256_result[100]), .C(
        SHA256_result[114]), .Y(f4_E_32[25]) );
  XOR3X2 U2197 ( .A(SHA256_result[104]), .B(SHA256_result[99]), .C(
        SHA256_result[118]), .Y(f4_E_32[29]) );
  XOR3X2 U2198 ( .A(SHA256_result[103]), .B(SHA256_result[98]), .C(
        SHA256_result[117]), .Y(f4_E_32[28]) );
  XOR3X2 U2199 ( .A(n66), .B(n149), .C(SHA256_result[246]), .Y(f3_A_32[20]) );
  NAND2X1 U2200 ( .A(n253), .B(read_counter[0]), .Y(N3079) );
  NAND3BX1 U2201 ( .AN(n255), .B(n1976), .C(n253), .Y(N3081) );
  OAI2BB1X1 U2202 ( .A0N(n972), .A1N(N3079), .B0(read_counter[2]), .Y(n1976)
         );
  NAND2X1 U2203 ( .A(n253), .B(n1977), .Y(N3080) );
  XNOR2X1 U2204 ( .A(n972), .B(read_counter[0]), .Y(n1977) );
  INVX1 U2205 ( .A(SHA256_result[60]), .Y(n935) );
  OAI2BB1X1 U2206 ( .A0N(SHA256_result[215]), .A1N(n137), .B0(n592), .Y(
        f2_ABC_32[23]) );
  OAI21XL U2207 ( .A0(SHA256_result[215]), .A1(n137), .B0(SHA256_result[183]), 
        .Y(n592) );
  OAI2BB1X1 U2208 ( .A0N(SHA256_result[217]), .A1N(n135), .B0(n590), .Y(
        f2_ABC_32[25]) );
  OAI21XL U2209 ( .A0(SHA256_result[217]), .A1(n135), .B0(SHA256_result[185]), 
        .Y(n590) );
  OAI2BB1X1 U2210 ( .A0N(SHA256_result[216]), .A1N(n136), .B0(n591), .Y(
        f2_ABC_32[24]) );
  OAI21XL U2211 ( .A0(SHA256_result[216]), .A1(n136), .B0(SHA256_result[184]), 
        .Y(n591) );
  OAI2BB1X1 U2212 ( .A0N(SHA256_result[218]), .A1N(n134), .B0(n589), .Y(
        f2_ABC_32[26]) );
  OAI21XL U2213 ( .A0(SHA256_result[218]), .A1(n134), .B0(SHA256_result[186]), 
        .Y(n589) );
  XOR3X2 U2214 ( .A(SHA256_result[105]), .B(SHA256_result[100]), .C(
        SHA256_result[119]), .Y(f4_E_32[30]) );
  MX2X1 U2215 ( .A(SHA256_result[62]), .B(SHA256_result[94]), .S0(
        SHA256_result[126]), .Y(f1_EFG_32[30]) );
  XOR3X2 U2216 ( .A(n143), .B(n152), .C(SHA256_result[252]), .Y(f3_A_32[26])
         );
  NOR2X1 U2217 ( .A(n1383), .B(n1388), .Y(n2226) );
  NOR2X1 U2218 ( .A(n768), .B(n1370), .Y(n2191) );
  AOI211X1 U2219 ( .A0(n747), .A1(n1383), .B0(n2259), .C0(n2247), .Y(n2395) );
  OAI2BB1X1 U2220 ( .A0N(SHA256_result[220]), .A1N(SHA256_result[252]), .B0(
        n587), .Y(f2_ABC_32[28]) );
  OAI21XL U2221 ( .A0(SHA256_result[220]), .A1(SHA256_result[252]), .B0(
        SHA256_result[188]), .Y(n587) );
  OAI2BB1X1 U2222 ( .A0N(SHA256_result[219]), .A1N(n133), .B0(n588), .Y(
        f2_ABC_32[27]) );
  OAI21XL U2223 ( .A0(SHA256_result[219]), .A1(n133), .B0(SHA256_result[187]), 
        .Y(n588) );
  OAI2BB1X1 U2224 ( .A0N(SHA256_result[222]), .A1N(n131), .B0(n585), .Y(
        f2_ABC_32[30]) );
  OAI21XL U2225 ( .A0(SHA256_result[222]), .A1(n131), .B0(SHA256_result[190]), 
        .Y(n585) );
  OAI2BB1X1 U2226 ( .A0N(SHA256_result[221]), .A1N(n132), .B0(n586), .Y(
        f2_ABC_32[29]) );
  OAI21XL U2227 ( .A0(SHA256_result[221]), .A1(n132), .B0(SHA256_result[189]), 
        .Y(n586) );
  INVX1 U2228 ( .A(n2188), .Y(n767) );
  AOI221X1 U2229 ( .A0(n345), .A1(n2189), .B0(n1388), .B1(n2190), .C0(n2191), 
        .Y(n2188) );
  XOR3X2 U2230 ( .A(n140), .B(n149), .C(n25), .Y(f3_A_32[29]) );
  MX2X1 U2231 ( .A(SHA256_result[63]), .B(SHA256_result[95]), .S0(
        SHA256_result[127]), .Y(f1_EFG_32[31]) );
  NOR2X1 U2232 ( .A(n781), .B(n1388), .Y(n2136) );
  NOR2X1 U2233 ( .A(n788), .B(n1388), .Y(n2144) );
  OAI222XL U2234 ( .A0(n757), .A1(n1388), .B0(n2246), .B1(n160), .C0(n774), 
        .C1(n1393), .Y(n2245) );
  AOI211X1 U2235 ( .A0(n1383), .A1(n2138), .B0(n2219), .C0(n2247), .Y(n2246)
         );
  OAI222XL U2236 ( .A0(n797), .A1(n127), .B0(n1393), .B1(n773), .C0(n1388), 
        .C1(n755), .Y(n2281) );
  OAI221XL U2237 ( .A0(n794), .A1(n1393), .B0(n1388), .B1(n756), .C0(n2184), 
        .Y(n2319) );
  NOR2X1 U2238 ( .A(n765), .B(n1388), .Y(n2315) );
  INVX1 U2239 ( .A(read_counter[2]), .Y(n973) );
  NOR2X1 U2240 ( .A(n1383), .B(n347), .Y(n2121) );
  NOR2X1 U2241 ( .A(n777), .B(n1388), .Y(n2202) );
  OAI31X1 U2242 ( .A0(n769), .A1(n791), .A2(n1383), .B0(n2210), .Y(n2284) );
  NOR2X1 U2243 ( .A(n788), .B(n1383), .Y(n2128) );
  NOR2X1 U2244 ( .A(n1383), .B(n346), .Y(n2324) );
  NAND2X1 U2245 ( .A(n782), .B(n1388), .Y(n2133) );
  NAND2X1 U2246 ( .A(n114), .B(n1383), .Y(n2173) );
  NOR2X1 U2247 ( .A(n764), .B(n1383), .Y(n2124) );
  NOR2X1 U2248 ( .A(n2166), .B(n1388), .Y(n2198) );
  NOR2X1 U2249 ( .A(n777), .B(n1383), .Y(n2287) );
  NOR2X1 U2250 ( .A(n127), .B(n1388), .Y(n2185) );
  NAND2X1 U2251 ( .A(n31), .B(n1388), .Y(n2274) );
  NOR2X1 U2252 ( .A(n796), .B(n1370), .Y(n2267) );
  NOR2X1 U2253 ( .A(n765), .B(n1383), .Y(n2302) );
  INVX1 U2254 ( .A(read_counter[0]), .Y(n971) );
  AOI31X1 U2255 ( .A0(n1388), .A1(n1370), .A2(n2138), .B0(n2231), .Y(n2310) );
  AOI21X1 U2256 ( .A0(n2165), .A1(n758), .B0(n1388), .Y(n2164) );
  AOI21X1 U2257 ( .A0(n753), .A1(n2181), .B0(n1388), .Y(n2295) );
  OAI22X1 U2258 ( .A0(n1142), .A1(n1985), .B0(n1984), .B1(n464), .Y(n376) );
  OAI22X1 U2259 ( .A0(n1141), .A1(n1985), .B0(n1984), .B1(n460), .Y(n378) );
  OAI22X1 U2260 ( .A0(n1143), .A1(n244), .B0(n246), .B1(n468), .Y(n374) );
  OAI22X1 U2261 ( .A0(n900), .A1(n246), .B0(n1144), .B1(n244), .Y(n2017) );
  OAI22X1 U2262 ( .A0(n1140), .A1(n1985), .B0(n1984), .B1(n455), .Y(n380) );
  NAND3X1 U2263 ( .A(n971), .B(n973), .C(read_counter[1]), .Y(n1985) );
  NAND3X1 U2264 ( .A(read_counter[0]), .B(n973), .C(read_counter[1]), .Y(n1984) );
  OAI21XL U2265 ( .A0(round[3]), .A1(n2370), .B0(n2371), .Y(n2369) );
  AOI22X1 U2266 ( .A0(n765), .A1(n1370), .B0(n2135), .B1(n159), .Y(n2370) );
  OAI21XL U2267 ( .A0(n2183), .A1(n2326), .B0(n346), .Y(n2371) );
  BUFX3 U2268 ( .A(round[4]), .Y(n159) );
  OAI2BB1X1 U2269 ( .A0N(SHA256_result[223]), .A1N(n25), .B0(n584), .Y(
        f2_ABC_32[31]) );
  OAI21XL U2270 ( .A0(SHA256_result[223]), .A1(n25), .B0(SHA256_result[191]), 
        .Y(n584) );
  NOR2X1 U2271 ( .A(n1388), .B(n346), .Y(n2363) );
  NOR3X1 U2272 ( .A(read_counter[0]), .B(read_counter[1]), .C(n973), .Y(n1986)
         );
  NOR3X1 U2273 ( .A(read_counter[1]), .B(read_counter[2]), .C(n971), .Y(n1982)
         );
  NOR3X1 U2274 ( .A(n756), .B(n1383), .C(n1370), .Y(n2237) );
  INVXL U2275 ( .A(SHA256_result[103]), .Y(n520) );
  INVXL U2276 ( .A(SHA256_result[109]), .Y(n889) );
  INVXL U2277 ( .A(SHA256_result[99]), .Y(n535) );
  INVXL U2278 ( .A(SHA256_result[110]), .Y(n890) );
  INVXL U2279 ( .A(SHA256_result[104]), .Y(n515) );
  INVXL U2280 ( .A(n67), .Y(n542) );
  INVXL U2281 ( .A(SHA256_result[108]), .Y(n888) );
  INVXL U2282 ( .A(SHA256_result[102]), .Y(n524) );
  INVXL U2283 ( .A(SHA256_result[105]), .Y(n510) );
  AND2X2 U2284 ( .A(n255), .B(SHA256_result[25]), .Y(n373) );
  AND2X2 U2285 ( .A(n255), .B(SHA256_result[26]), .Y(n375) );
  AND2X2 U2286 ( .A(n255), .B(SHA256_result[27]), .Y(n377) );
  AND2X2 U2287 ( .A(n255), .B(SHA256_result[28]), .Y(n379) );
  AND2X2 U2288 ( .A(n255), .B(SHA256_result[30]), .Y(n383) );
  AND2X2 U2289 ( .A(n255), .B(SHA256_result[31]), .Y(n385) );
  AND2X2 U2290 ( .A(n255), .B(SHA256_result[29]), .Y(n381) );
  INVX1 U2291 ( .A(SHA256_result[94]), .Y(n912) );
  INVX1 U2292 ( .A(SHA256_result[218]), .Y(n823) );
  INVX1 U2293 ( .A(SHA256_result[211]), .Y(n816) );
  INVX1 U2294 ( .A(SHA256_result[191]), .Y(n855) );
  INVX1 U2295 ( .A(SHA256_result[184]), .Y(n848) );
  INVX1 U2296 ( .A(SHA256_result[214]), .Y(n819) );
  INVX1 U2297 ( .A(SHA256_result[222]), .Y(n827) );
  INVX1 U2298 ( .A(SHA256_result[215]), .Y(n820) );
  INVX1 U2299 ( .A(SHA256_result[212]), .Y(n817) );
  INVX1 U2300 ( .A(SHA256_result[221]), .Y(n826) );
  INVX1 U2301 ( .A(SHA256_result[220]), .Y(n825) );
  INVX1 U2302 ( .A(SHA256_result[219]), .Y(n824) );
  INVX1 U2303 ( .A(SHA256_result[213]), .Y(n818) );
  INVX1 U2304 ( .A(SHA256_result[156]), .Y(n885) );
  INVX1 U2305 ( .A(SHA256_result[155]), .Y(n884) );
  INVX1 U2306 ( .A(SHA256_result[190]), .Y(n854) );
  INVX1 U2307 ( .A(SHA256_result[185]), .Y(n849) );
  INVX1 U2308 ( .A(SHA256_result[183]), .Y(n847) );
  INVX1 U2309 ( .A(SHA256_result[180]), .Y(n844) );
  INVX1 U2310 ( .A(SHA256_result[189]), .Y(n853) );
  INVX1 U2311 ( .A(SHA256_result[186]), .Y(n850) );
  INVX1 U2312 ( .A(SHA256_result[182]), .Y(n846) );
  INVX1 U2313 ( .A(SHA256_result[179]), .Y(n843) );
  INVX1 U2314 ( .A(SHA256_result[148]), .Y(n877) );
  INVX1 U2315 ( .A(SHA256_result[149]), .Y(n878) );
  INVX1 U2316 ( .A(SHA256_result[63]), .Y(n938) );
  INVX1 U2317 ( .A(SHA256_result[61]), .Y(n936) );
  INVX1 U2318 ( .A(SHA256_result[158]), .Y(n887) );
  INVX1 U2319 ( .A(SHA256_result[139]), .Y(n868) );
  INVX1 U2320 ( .A(SHA256_result[137]), .Y(n866) );
  INVX1 U2321 ( .A(SHA256_result[135]), .Y(n864) );
  INVX1 U2322 ( .A(SHA256_result[134]), .Y(n863) );
  INVX1 U2323 ( .A(SHA256_result[130]), .Y(n859) );
  INVX1 U2324 ( .A(SHA256_result[93]), .Y(n911) );
  INVX1 U2325 ( .A(SHA256_result[153]), .Y(n882) );
  INVX1 U2326 ( .A(SHA256_result[151]), .Y(n880) );
  INVX1 U2327 ( .A(SHA256_result[26]), .Y(n966) );
  INVX1 U2328 ( .A(SHA256_result[31]), .Y(n939) );
  INVX1 U2329 ( .A(SHA256_result[217]), .Y(n822) );
  INVX1 U2330 ( .A(SHA256_result[216]), .Y(n821) );
  INVX1 U2331 ( .A(SHA256_result[29]), .Y(n969) );
  INVX1 U2332 ( .A(SHA256_result[95]), .Y(n901) );
  INVX1 U2333 ( .A(SHA256_result[131]), .Y(n860) );
  INVX1 U2334 ( .A(SHA256_result[223]), .Y(n798) );
  INVX1 U2335 ( .A(SHA256_result[188]), .Y(n852) );
  INVX1 U2336 ( .A(SHA256_result[187]), .Y(n851) );
  INVX1 U2337 ( .A(SHA256_result[181]), .Y(n845) );
  INVX1 U2338 ( .A(SHA256_result[143]), .Y(n872) );
  INVX1 U2339 ( .A(SHA256_result[154]), .Y(n883) );
  INVX1 U2340 ( .A(SHA256_result[152]), .Y(n881) );
  INVX1 U2341 ( .A(SHA256_result[157]), .Y(n886) );
  INVX1 U2342 ( .A(SHA256_result[150]), .Y(n879) );
  INVX1 U2343 ( .A(SHA256_result[147]), .Y(n876) );
  INVX1 U2344 ( .A(SHA256_result[145]), .Y(n874) );
  INVX1 U2345 ( .A(SHA256_result[141]), .Y(n870) );
  INVX1 U2346 ( .A(SHA256_result[140]), .Y(n869) );
  INVX1 U2347 ( .A(SHA256_result[138]), .Y(n867) );
  INVX1 U2348 ( .A(SHA256_result[136]), .Y(n865) );
  INVX1 U2349 ( .A(SHA256_result[133]), .Y(n862) );
  INVX1 U2350 ( .A(SHA256_result[132]), .Y(n861) );
  INVX1 U2351 ( .A(SHA256_result[159]), .Y(n856) );
  INVX1 U2352 ( .A(SHA256_result[144]), .Y(n873) );
  INVX1 U2353 ( .A(SHA256_result[142]), .Y(n871) );
  INVX1 U2354 ( .A(SHA256_result[30]), .Y(n970) );
  INVX1 U2355 ( .A(SHA256_result[28]), .Y(n968) );
  INVX1 U2356 ( .A(SHA256_result[27]), .Y(n967) );
  INVX1 U2357 ( .A(SHA256_result[25]), .Y(n965) );
  INVX1 U2358 ( .A(SHA256_result[24]), .Y(n964) );
  INVX1 U2359 ( .A(SHA256_result[23]), .Y(n963) );
  INVX1 U2360 ( .A(SHA256_result[22]), .Y(n962) );
  INVX1 U2361 ( .A(SHA256_result[146]), .Y(n875) );
  AOI21XL U2362 ( .A0(next_E[23]), .A1(n276), .B0(n474), .Y(n475) );
  AOI21XL U2363 ( .A0(next_E[22]), .A1(n275), .B0(n476), .Y(n477) );
  NAND2XL U2364 ( .A(next_A[29]), .B(n276), .Y(n622) );
  AOI21XL U2365 ( .A0(next_E[29]), .A1(n276), .B0(n453), .Y(n454) );
  INVXL U2366 ( .A(next_A[18]), .Y(n656) );
  INVXL U2367 ( .A(next_A[19]), .Y(n655) );
  XOR3X2 U2368 ( .A(SHA256_result[111]), .B(SHA256_result[106]), .C(
        SHA256_result[125]), .Y(f4_E_32[4]) );
  XOR3X2 U2369 ( .A(SHA256_result[120]), .B(SHA256_result[107]), .C(n51), .Y(
        f4_E_32[18]) );
  XOR3X2 U2370 ( .A(SHA256_result[112]), .B(SHA256_result[98]), .C(n51), .Y(
        f4_E_32[23]) );
  OAI21XL U2371 ( .A0(n162), .A1(n911), .B0(n1612), .Y(n2673) );
  NOR2X1 U2372 ( .A(n166), .B(n452), .Y(n453) );
  OAI21XL U2373 ( .A0(n342), .A1(n452), .B0(n451), .Y(n2609) );
  OAI22X1 U2374 ( .A0(n1985), .A1(n911), .B0(n1984), .B1(n452), .Y(n382) );
  INVXL U2375 ( .A(n43), .Y(n651) );
  AOI21XL U2376 ( .A0(next_E[25]), .A1(n276), .B0(n469), .Y(n470) );
  AOI21XL U2377 ( .A0(next_E[26]), .A1(n276), .B0(n465), .Y(n466) );
  NAND2XL U2378 ( .A(next_A[27]), .B(n276), .Y(n627) );
  AOI21XL U2379 ( .A0(next_A[23]), .A1(n275), .B0(n643), .Y(n644) );
  NAND2XL U2380 ( .A(next_A[25]), .B(n276), .Y(n635) );
  AOI21XL U2381 ( .A0(next_A[26]), .A1(n275), .B0(n631), .Y(n632) );
  MX2X4 U2382 ( .A(n50), .B(SHA256_result[70]), .S0(SHA256_result[102]), .Y(
        f1_EFG_32[6]) );
  MXI2X4 U2383 ( .A(n447), .B(n1167), .S0(n67), .Y(f1_EFG_32[1]) );
  XOR3X4 U2384 ( .A(SHA256_result[109]), .B(SHA256_result[104]), .C(
        SHA256_result[123]), .Y(f4_E_32[2]) );
endmodule


module controller_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module controller ( clk, reset, first_block, last_block, output_enable, busy, 
        inner_busy );
  input clk, reset, first_block, last_block;
  output output_enable, busy, inner_busy;
  wire   N11, N24, N25, N26, N27, N28, N29, N30, N47, N48, N49, n12, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n9, n10, n11, n13;
  wire   [1:0] state;
  wire   [6:0] counter1;
  wire   [2:0] counter2;

  CLKINVX4 U24 ( .A(reset), .Y(n12) );
  controller_DW01_inc_0 add_82 ( .A(counter1), .SUM({N30, N29, N28, N27, N26, 
        N25, N24}) );
  DFFHQX1 counter2_reg_2_ ( .D(N49), .CK(clk), .Q(counter2[2]) );
  DFFHQX1 counter2_reg_0_ ( .D(N47), .CK(clk), .Q(counter2[0]) );
  DFFHQX1 counter2_reg_1_ ( .D(N48), .CK(clk), .Q(counter2[1]) );
  DFFTRX1 counter1_reg_6_ ( .D(N30), .RN(n19), .CK(clk), .Q(counter1[6]) );
  DFFTRX1 counter1_reg_5_ ( .D(N29), .RN(n19), .CK(clk), .Q(counter1[5]) );
  DFFTRX1 counter1_reg_4_ ( .D(N28), .RN(n19), .CK(clk), .Q(counter1[4]) );
  DFFTRX1 counter1_reg_3_ ( .D(N27), .RN(n19), .CK(clk), .Q(counter1[3]) );
  DFFTRX1 counter1_reg_2_ ( .D(N26), .RN(n19), .CK(clk), .Q(counter1[2]) );
  DFFTRX1 counter1_reg_1_ ( .D(N25), .RN(n19), .CK(clk), .Q(counter1[1]) );
  DFFTRX1 counter1_reg_0_ ( .D(N24), .RN(n19), .CK(clk), .Q(counter1[0]) );
  DFFHQX1 state_reg_1_ ( .D(N11), .CK(clk), .Q(state[1]) );
  DFFTRX1 state_reg_0_ ( .D(n12), .RN(n10), .CK(clk), .Q(state[0]) );
  NOR2BX2 U3 ( .AN(state[1]), .B(state[0]), .Y(output_enable) );
  NOR2BX1 U4 ( .AN(state[0]), .B(state[1]), .Y(inner_busy) );
  NOR2XL U5 ( .A(state[1]), .B(state[0]), .Y(n14) );
  NAND2XL U6 ( .A(output_enable), .B(n12), .Y(n17) );
  NAND3XL U7 ( .A(n9), .B(n12), .C(inner_busy), .Y(n21) );
  AOI22XL U8 ( .A0(first_block), .A1(n14), .B0(inner_busy), .B1(n22), .Y(n23)
         );
  INVX1 U9 ( .A(n14), .Y(busy) );
  INVX1 U10 ( .A(n22), .Y(n9) );
  AOI211X1 U11 ( .A0(n13), .A1(n20), .B0(n9), .C0(reset), .Y(n19) );
  INVX1 U12 ( .A(last_block), .Y(n13) );
  INVX1 U13 ( .A(n23), .Y(n10) );
  OAI211X1 U14 ( .A0(counter2[2]), .A1(n17), .B0(n21), .C0(n15), .Y(N11) );
  AOI2BB1X1 U15 ( .A0N(counter2[1]), .A1N(n17), .B0(N47), .Y(n15) );
  NOR2X1 U16 ( .A(n17), .B(counter2[0]), .Y(N47) );
  OAI21XL U17 ( .A0(n15), .A1(n11), .B0(n16), .Y(N49) );
  NAND4BXL U18 ( .AN(n17), .B(counter2[1]), .C(counter2[0]), .D(n11), .Y(n16)
         );
  INVX1 U19 ( .A(counter2[2]), .Y(n11) );
  NOR2X1 U20 ( .A(n18), .B(n17), .Y(N48) );
  XNOR2X1 U21 ( .A(counter2[0]), .B(counter2[1]), .Y(n18) );
  NAND2X1 U22 ( .A(counter1[6]), .B(n20), .Y(n22) );
  NOR4X1 U23 ( .A(counter1[2]), .B(counter1[1]), .C(counter1[0]), .D(n24), .Y(
        n20) );
  OR3XL U25 ( .A(counter1[5]), .B(counter1[4]), .C(counter1[3]), .Y(n24) );
endmodule


module top ( clk, reset, data, write_enable, last_block, first_block, busy, 
        digest, output_enable );
  input [31:0] data;
  output [31:0] digest;
  input clk, reset, write_enable, last_block, first_block;
  output busy, output_enable;
  wire   inner_busy;
  wire   [31:0] Wt;

  message_schedule our_message_schedule ( .clk(clk), .reset(reset), .data(data), .write_enable(write_enable), .inner_busy(inner_busy), .Wt(Wt) );
  hash_core our_hash_core ( .clk(clk), .reset(reset), .Wt(Wt), .inner_busy(
        inner_busy), .first_block(first_block), .output_enable(output_enable), 
        .digest(digest) );
  controller our_controller ( .clk(clk), .reset(reset), .first_block(
        first_block), .last_block(last_block), .output_enable(output_enable), 
        .busy(busy), .inner_busy(inner_busy) );
endmodule


module sha256_chip ( clk, reset, data, write_enable, last_block, first_block, 
        busy, digest, output_enable );
  input [31:0] data;
  output [31:0] digest;
  input clk, reset, write_enable, last_block, first_block;
  output busy, output_enable;
  wire   net_clk, net_reset, net_write_enable, net_last_block, net_first_block,
         net_busy, net_output_enable;
  wire   [31:0] net_data;
  wire   [31:0] net_digest;

  PIW PIW_clk ( .PAD(clk), .C(net_clk) );
  PIW PIW_reset ( .PAD(reset), .C(net_reset) );
  PIW PIW_data0 ( .PAD(data[0]), .C(net_data[0]) );
  PIW PIW_data1 ( .PAD(data[1]), .C(net_data[1]) );
  PIW PIW_data2 ( .PAD(data[2]), .C(net_data[2]) );
  PIW PIW_data3 ( .PAD(data[3]), .C(net_data[3]) );
  PIW PIW_data4 ( .PAD(data[4]), .C(net_data[4]) );
  PIW PIW_data5 ( .PAD(data[5]), .C(net_data[5]) );
  PIW PIW_data6 ( .PAD(data[6]), .C(net_data[6]) );
  PIW PIW_data7 ( .PAD(data[7]), .C(net_data[7]) );
  PIW PIW_data8 ( .PAD(data[8]), .C(net_data[8]) );
  PIW PIW_data9 ( .PAD(data[9]), .C(net_data[9]) );
  PIW PIW_data10 ( .PAD(data[10]), .C(net_data[10]) );
  PIW PIW_data11 ( .PAD(data[11]), .C(net_data[11]) );
  PIW PIW_data12 ( .PAD(data[12]), .C(net_data[12]) );
  PIW PIW_data13 ( .PAD(data[13]), .C(net_data[13]) );
  PIW PIW_data14 ( .PAD(data[14]), .C(net_data[14]) );
  PIW PIW_data15 ( .PAD(data[15]), .C(net_data[15]) );
  PIW PIW_data16 ( .PAD(data[16]), .C(net_data[16]) );
  PIW PIW_data17 ( .PAD(data[17]), .C(net_data[17]) );
  PIW PIW_data18 ( .PAD(data[18]), .C(net_data[18]) );
  PIW PIW_data19 ( .PAD(data[19]), .C(net_data[19]) );
  PIW PIW_data20 ( .PAD(data[20]), .C(net_data[20]) );
  PIW PIW_data21 ( .PAD(data[21]), .C(net_data[21]) );
  PIW PIW_data22 ( .PAD(data[22]), .C(net_data[22]) );
  PIW PIW_data23 ( .PAD(data[23]), .C(net_data[23]) );
  PIW PIW_data24 ( .PAD(data[24]), .C(net_data[24]) );
  PIW PIW_data25 ( .PAD(data[25]), .C(net_data[25]) );
  PIW PIW_data26 ( .PAD(data[26]), .C(net_data[26]) );
  PIW PIW_data27 ( .PAD(data[27]), .C(net_data[27]) );
  PIW PIW_data28 ( .PAD(data[28]), .C(net_data[28]) );
  PIW PIW_data29 ( .PAD(data[29]), .C(net_data[29]) );
  PIW PIW_data30 ( .PAD(data[30]), .C(net_data[30]) );
  PIW PIW_data31 ( .PAD(data[31]), .C(net_data[31]) );
  PIW PIW_write_enable ( .PAD(write_enable), .C(net_write_enable) );
  PIW PIW_last_block ( .PAD(last_block), .C(net_last_block) );
  PIW PIW_first_block ( .PAD(first_block), .C(net_first_block) );
  PO8W PO8W_busy ( .I(net_busy), .PAD(busy) );
  PO8W PO8W_digest0 ( .I(net_digest[0]), .PAD(digest[0]) );
  PO8W PO8W_digest1 ( .I(net_digest[1]), .PAD(digest[1]) );
  PO8W PO8W_digest2 ( .I(net_digest[2]), .PAD(digest[2]) );
  PO8W PO8W_digest3 ( .I(net_digest[3]), .PAD(digest[3]) );
  PO8W PO8W_digest4 ( .I(net_digest[4]), .PAD(digest[4]) );
  PO8W PO8W_digest5 ( .I(net_digest[5]), .PAD(digest[5]) );
  PO8W PO8W_digest6 ( .I(net_digest[6]), .PAD(digest[6]) );
  PO8W PO8W_digest7 ( .I(net_digest[7]), .PAD(digest[7]) );
  PO8W PO8W_digest8 ( .I(net_digest[8]), .PAD(digest[8]) );
  PO8W PO8W_digest9 ( .I(net_digest[9]), .PAD(digest[9]) );
  PO8W PO8W_digest10 ( .I(net_digest[10]), .PAD(digest[10]) );
  PO8W PO8W_digest11 ( .I(net_digest[11]), .PAD(digest[11]) );
  PO8W PO8W_digest12 ( .I(net_digest[12]), .PAD(digest[12]) );
  PO8W PO8W_digest13 ( .I(net_digest[13]), .PAD(digest[13]) );
  PO8W PO8W_digest14 ( .I(net_digest[14]), .PAD(digest[14]) );
  PO8W PO8W_digest15 ( .I(net_digest[15]), .PAD(digest[15]) );
  PO8W PO8W_digest16 ( .I(net_digest[16]), .PAD(digest[16]) );
  PO8W PO8W_digest17 ( .I(net_digest[17]), .PAD(digest[17]) );
  PO8W PO8W_digest18 ( .I(net_digest[18]), .PAD(digest[18]) );
  PO8W PO8W_digest19 ( .I(net_digest[19]), .PAD(digest[19]) );
  PO8W PO8W_digest20 ( .I(net_digest[20]), .PAD(digest[20]) );
  PO8W PO8W_digest21 ( .I(net_digest[21]), .PAD(digest[21]) );
  PO8W PO8W_digest22 ( .I(net_digest[22]), .PAD(digest[22]) );
  PO8W PO8W_digest23 ( .I(net_digest[23]), .PAD(digest[23]) );
  PO8W PO8W_digest24 ( .I(net_digest[24]), .PAD(digest[24]) );
  PO8W PO8W_digest25 ( .I(net_digest[25]), .PAD(digest[25]) );
  PO8W PO8W_digest26 ( .I(net_digest[26]), .PAD(digest[26]) );
  PO8W PO8W_digest27 ( .I(net_digest[27]), .PAD(digest[27]) );
  PO8W PO8W_digest28 ( .I(net_digest[28]), .PAD(digest[28]) );
  PO8W PO8W_digest29 ( .I(net_digest[29]), .PAD(digest[29]) );
  PO8W PO8W_digest30 ( .I(net_digest[30]), .PAD(digest[30]) );
  PO8W PO8W_digest31 ( .I(net_digest[31]), .PAD(digest[31]) );
  PO8W PO8W_output_enable ( .I(net_output_enable), .PAD(output_enable) );
  top inst_top ( .clk(net_clk), .reset(net_reset), .data(net_data), 
        .write_enable(net_write_enable), .last_block(net_last_block), 
        .first_block(net_first_block), .busy(net_busy), .digest(net_digest), 
        .output_enable(net_output_enable) );
endmodule


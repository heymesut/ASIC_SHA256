
module message_schedule_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module message_schedule_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module message_schedule_DW01_add_19 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221;

  AOI21X2 U2 ( .A0(n169), .A1(n174), .B0(n175), .Y(n172) );
  OAI21X2 U3 ( .A0(n217), .A1(n218), .B0(n41), .Y(n174) );
  NOR2X1 U4 ( .A(n193), .B(n168), .Y(n4) );
  NAND2X1 U5 ( .A(n98), .B(n106), .Y(n119) );
  INVX4 U6 ( .A(n176), .Y(n175) );
  CLKINVX3 U7 ( .A(n83), .Y(n81) );
  NAND3BX1 U8 ( .AN(n105), .B(n111), .C(n112), .Y(n99) );
  OAI21X4 U9 ( .A0(n172), .A1(n168), .B0(n173), .Y(n171) );
  NOR2X1 U10 ( .A(A[30]), .B(B[30]), .Y(n10) );
  NAND2X4 U11 ( .A(n89), .B(n79), .Y(n87) );
  NAND2X1 U12 ( .A(B[25]), .B(A[25]), .Y(n79) );
  OAI2BB1X2 U13 ( .A0N(n152), .A1N(n133), .B0(n140), .Y(n149) );
  NAND4BBX2 U14 ( .AN(n32), .BN(n12), .C(n30), .D(n24), .Y(n177) );
  OR2X4 U15 ( .A(A[19]), .B(B[19]), .Y(n142) );
  NAND4BBX2 U16 ( .AN(n20), .BN(n16), .C(n197), .D(n196), .Y(n168) );
  INVX1 U17 ( .A(n213), .Y(n32) );
  INVX1 U18 ( .A(n198), .Y(n16) );
  INVX1 U19 ( .A(n118), .Y(n105) );
  INVX1 U20 ( .A(n148), .Y(n130) );
  NAND3X1 U21 ( .A(n213), .B(n30), .C(n214), .Y(n212) );
  INVX1 U22 ( .A(n133), .Y(n138) );
  AOI21X2 U23 ( .A0(n159), .A1(n160), .B0(n161), .Y(n158) );
  INVX1 U24 ( .A(n162), .Y(n161) );
  OR2X2 U25 ( .A(A[3]), .B(B[3]), .Y(n216) );
  OAI2BB1X2 U26 ( .A0N(n194), .A1N(n195), .B0(n196), .Y(n173) );
  OAI2BB1X1 U27 ( .A0N(n211), .A1N(n212), .B0(n24), .Y(n176) );
  NOR2X1 U28 ( .A(A[25]), .B(B[25]), .Y(n77) );
  OAI21X1 U29 ( .A0(n51), .A1(n52), .B0(n53), .Y(n50) );
  NAND3BX2 U30 ( .AN(n127), .B(n128), .C(n129), .Y(n126) );
  NOR2BX2 U31 ( .AN(n200), .B(n201), .Y(n194) );
  CLKINVX3 U32 ( .A(n202), .Y(n201) );
  OR2X4 U33 ( .A(A[23]), .B(B[23]), .Y(n112) );
  NAND2XL U34 ( .A(B[15]), .B(A[15]), .Y(n162) );
  AOI21X2 U35 ( .A0(n101), .A1(n102), .B0(n103), .Y(n100) );
  NAND2X1 U36 ( .A(B[14]), .B(A[14]), .Y(n165) );
  NAND2X4 U37 ( .A(B[5]), .B(A[5]), .Y(n33) );
  NAND2X4 U38 ( .A(n121), .B(n122), .Y(n98) );
  NOR2X2 U39 ( .A(n109), .B(n110), .Y(n101) );
  CLKINVX3 U40 ( .A(n112), .Y(n109) );
  INVX3 U41 ( .A(n179), .Y(n167) );
  OAI21X2 U42 ( .A0(n183), .A1(n167), .B0(n165), .Y(n181) );
  NOR2X2 U43 ( .A(n36), .B(n177), .Y(n6) );
  OR2X4 U44 ( .A(A[11]), .B(B[11]), .Y(n196) );
  XNOR2X4 U45 ( .A(n7), .B(n66), .Y(SUM[29]) );
  NAND2X4 U46 ( .A(n54), .B(n1), .Y(n56) );
  OR2X4 U47 ( .A(n6), .B(n175), .Y(n17) );
  INVX8 U48 ( .A(n68), .Y(n58) );
  NAND2X4 U49 ( .A(B[7]), .B(A[7]), .Y(n23) );
  NOR2BX1 U50 ( .AN(n162), .B(n166), .Y(n182) );
  INVX2 U51 ( .A(n180), .Y(n166) );
  NAND4BX1 U52 ( .AN(n11), .B(n178), .C(n179), .D(n180), .Y(n170) );
  OAI211X2 U53 ( .A0(n11), .A1(n163), .B0(n164), .C0(n165), .Y(n160) );
  XOR2X2 U54 ( .A(n181), .B(n182), .Y(SUM[15]) );
  NAND2BX4 U55 ( .AN(n170), .B(n171), .Y(n157) );
  AOI21X4 U56 ( .A0(n48), .A1(n49), .B0(n50), .Y(n47) );
  OAI21X2 U57 ( .A0(n57), .A1(n58), .B0(n59), .Y(n49) );
  OR2X4 U58 ( .A(A[15]), .B(B[15]), .Y(n180) );
  XNOR3X4 U59 ( .A(B[30]), .B(A[30]), .C(n9), .Y(SUM[30]) );
  NAND2XL U60 ( .A(n196), .B(n202), .Y(n204) );
  NAND2X2 U61 ( .A(B[11]), .B(A[11]), .Y(n202) );
  NOR2X4 U62 ( .A(n166), .B(n167), .Y(n159) );
  NAND2X1 U63 ( .A(B[27]), .B(A[27]), .Y(n76) );
  NAND3BX1 U64 ( .AN(n77), .B(n83), .C(n82), .Y(n71) );
  NAND2X4 U65 ( .A(n157), .B(n158), .Y(n128) );
  XNOR2X4 U66 ( .A(n8), .B(n84), .Y(SUM[27]) );
  NOR2BX2 U67 ( .AN(n82), .B(n81), .Y(n73) );
  OR2X4 U68 ( .A(A[27]), .B(B[27]), .Y(n82) );
  OAI21X4 U69 ( .A0(n189), .A1(n190), .B0(n163), .Y(n187) );
  INVX4 U70 ( .A(n191), .Y(n190) );
  INVX4 U71 ( .A(n184), .Y(n183) );
  NAND2X2 U72 ( .A(n90), .B(n91), .Y(n89) );
  OAI21X4 U73 ( .A0(n115), .A1(n110), .B0(n108), .Y(n113) );
  INVX2 U74 ( .A(n116), .Y(n115) );
  XOR2X4 U75 ( .A(n113), .B(n114), .Y(SUM[23]) );
  OAI21X4 U76 ( .A0(n70), .A1(n71), .B0(n72), .Y(n68) );
  AOI21X2 U77 ( .A0(n73), .A1(n74), .B0(n75), .Y(n72) );
  XOR2X4 U78 ( .A(n46), .B(n47), .Y(SUM[31]) );
  NAND2X2 U79 ( .A(n70), .B(n93), .Y(n91) );
  NAND2X4 U80 ( .A(n94), .B(n95), .Y(n70) );
  INVXL U81 ( .A(n30), .Y(n26) );
  OR2X4 U82 ( .A(A[6]), .B(B[6]), .Y(n30) );
  NAND2X2 U83 ( .A(B[6]), .B(A[6]), .Y(n27) );
  NAND2XL U84 ( .A(B[18]), .B(A[18]), .Y(n141) );
  OAI21X4 U85 ( .A0(n57), .A1(n58), .B0(n59), .Y(n1) );
  INVX1 U86 ( .A(n174), .Y(n36) );
  OR2X2 U87 ( .A(n4), .B(n5), .Y(n191) );
  NAND2XL U88 ( .A(n17), .B(n203), .Y(n210) );
  NAND2XL U89 ( .A(B[13]), .B(A[13]), .Y(n164) );
  XOR2X1 U90 ( .A(n191), .B(n192), .Y(SUM[12]) );
  NOR2X1 U91 ( .A(n186), .B(n11), .Y(n2) );
  INVXL U92 ( .A(n164), .Y(n3) );
  OR2X2 U93 ( .A(n2), .B(n3), .Y(n184) );
  INVXL U94 ( .A(n173), .Y(n5) );
  INVX1 U95 ( .A(n17), .Y(n193) );
  OR2X2 U96 ( .A(A[7]), .B(B[7]), .Y(n24) );
  NAND2X1 U97 ( .A(B[8]), .B(A[8]), .Y(n19) );
  NAND2X1 U98 ( .A(B[22]), .B(A[22]), .Y(n108) );
  OR2X2 U99 ( .A(A[8]), .B(B[8]), .Y(n203) );
  NOR2BXL U100 ( .AN(n104), .B(n109), .Y(n114) );
  XOR2XL U101 ( .A(n69), .B(n58), .Y(SUM[28]) );
  NOR2X2 U102 ( .A(A[13]), .B(B[13]), .Y(n11) );
  OR2X4 U103 ( .A(A[26]), .B(B[26]), .Y(n83) );
  NAND2X1 U104 ( .A(B[4]), .B(A[4]), .Y(n37) );
  NAND2XL U105 ( .A(B[26]), .B(A[26]), .Y(n80) );
  OR2XL U106 ( .A(A[2]), .B(B[2]), .Y(n62) );
  OR2X1 U107 ( .A(A[12]), .B(B[12]), .Y(n178) );
  NAND2XL U108 ( .A(B[28]), .B(A[28]), .Y(n59) );
  CLKINVX2 U109 ( .A(n177), .Y(n169) );
  OAI21X4 U110 ( .A0(n98), .A1(n99), .B0(n100), .Y(n94) );
  INVX1 U111 ( .A(n60), .Y(n57) );
  NAND2X1 U112 ( .A(n15), .B(n19), .Y(n199) );
  OAI2BB1X1 U113 ( .A0N(n118), .A1N(n119), .B0(n107), .Y(n116) );
  NAND2X1 U114 ( .A(n33), .B(n37), .Y(n214) );
  INVX1 U115 ( .A(n142), .Y(n131) );
  NAND2X1 U116 ( .A(B[10]), .B(A[10]), .Y(n200) );
  NOR2X1 U117 ( .A(A[4]), .B(B[4]), .Y(n12) );
  NOR2X1 U118 ( .A(A[30]), .B(B[30]), .Y(n51) );
  NAND2X1 U119 ( .A(B[12]), .B(A[12]), .Y(n163) );
  NAND2X1 U120 ( .A(B[2]), .B(A[2]), .Y(n44) );
  NAND2X1 U121 ( .A(A[24]), .B(B[24]), .Y(n78) );
  NAND2X2 U122 ( .A(n125), .B(n126), .Y(n121) );
  INVX2 U123 ( .A(n111), .Y(n110) );
  NOR2BXL U124 ( .AN(n85), .B(n81), .Y(n88) );
  NOR2BXL U125 ( .AN(n79), .B(n77), .Y(n92) );
  NAND2XL U126 ( .A(n59), .B(n60), .Y(n69) );
  NAND2X1 U127 ( .A(n59), .B(n67), .Y(n7) );
  NAND2X1 U128 ( .A(n85), .B(n86), .Y(n8) );
  NAND2XL U129 ( .A(n68), .B(n60), .Y(n67) );
  NAND2XL U130 ( .A(n128), .B(n132), .Y(n154) );
  NOR2BXL U131 ( .AN(n141), .B(n130), .Y(n151) );
  INVXL U132 ( .A(n95), .Y(n97) );
  NOR2BXL U133 ( .AN(n165), .B(n167), .Y(n185) );
  NOR2BXL U134 ( .AN(n108), .B(n110), .Y(n117) );
  NOR2BXL U135 ( .AN(n107), .B(n105), .Y(n120) );
  NAND2XL U136 ( .A(n137), .B(n142), .Y(n146) );
  AOI21XL U137 ( .A0(n148), .A1(n149), .B0(n150), .Y(n147) );
  NAND2XL U138 ( .A(n132), .B(n133), .Y(n127) );
  INVXL U139 ( .A(n132), .Y(n156) );
  NOR2BXL U140 ( .AN(n140), .B(n138), .Y(n153) );
  AOI21XL U141 ( .A0(n197), .A1(n206), .B0(n207), .Y(n205) );
  NOR2BXL U142 ( .AN(n15), .B(n16), .Y(n14) );
  AND2X1 U143 ( .A(n200), .B(n197), .Y(n208) );
  NOR2BXL U144 ( .AN(n163), .B(n189), .Y(n192) );
  NOR2BXL U145 ( .AN(n19), .B(n20), .Y(n18) );
  NOR2BXL U146 ( .AN(n65), .B(n144), .Y(n143) );
  AND2X1 U147 ( .A(n41), .B(n216), .Y(n40) );
  AND2X2 U148 ( .A(n55), .B(n56), .Y(n9) );
  NAND2XL U149 ( .A(B[19]), .B(A[19]), .Y(n137) );
  NAND2XL U150 ( .A(B[23]), .B(A[23]), .Y(n104) );
  NAND2XL U151 ( .A(B[21]), .B(A[21]), .Y(n107) );
  NAND2XL U152 ( .A(B[17]), .B(A[17]), .Y(n140) );
  NAND2XL U153 ( .A(B[1]), .B(A[1]), .Y(n65) );
  NAND2XL U154 ( .A(A[29]), .B(B[29]), .Y(n52) );
  NAND2XL U155 ( .A(B[30]), .B(A[30]), .Y(n53) );
  NAND2XL U156 ( .A(B[3]), .B(A[3]), .Y(n41) );
  OR2XL U157 ( .A(A[20]), .B(B[20]), .Y(n122) );
  NOR2BX1 U158 ( .AN(n54), .B(n10), .Y(n48) );
  NAND2XL U159 ( .A(B[29]), .B(A[29]), .Y(n55) );
  NAND2XL U160 ( .A(B[24]), .B(A[24]), .Y(n93) );
  NAND2XL U161 ( .A(B[26]), .B(A[26]), .Y(n85) );
  INVXL U162 ( .A(n145), .Y(n64) );
  AND2X1 U163 ( .A(n145), .B(n221), .Y(SUM[0]) );
  OR2XL U164 ( .A(A[0]), .B(B[0]), .Y(n221) );
  NOR2X1 U165 ( .A(n131), .B(n130), .Y(n134) );
  NOR2X1 U166 ( .A(n130), .B(n131), .Y(n129) );
  OAI211X1 U167 ( .A0(n105), .A1(n106), .B0(n107), .C0(n108), .Y(n102) );
  INVX1 U168 ( .A(n104), .Y(n103) );
  OAI211X1 U169 ( .A0(n77), .A1(n78), .B0(n79), .C0(n80), .Y(n74) );
  AOI21X1 U170 ( .A0(n134), .A1(n135), .B0(n136), .Y(n125) );
  OAI211X1 U171 ( .A0(n138), .A1(n139), .B0(n140), .C0(n141), .Y(n135) );
  NAND3X1 U172 ( .A(n197), .B(n198), .C(n199), .Y(n195) );
  NOR2BX1 U173 ( .AN(n27), .B(n215), .Y(n211) );
  XOR2X1 U174 ( .A(n91), .B(n92), .Y(SUM[25]) );
  XOR2X1 U175 ( .A(n87), .B(n88), .Y(SUM[26]) );
  NAND2X1 U176 ( .A(n76), .B(n82), .Y(n84) );
  NAND2X1 U177 ( .A(n54), .B(n55), .Y(n66) );
  NAND2X1 U178 ( .A(n87), .B(n83), .Y(n86) );
  INVX1 U179 ( .A(n137), .Y(n136) );
  INVX1 U180 ( .A(n23), .Y(n215) );
  OAI21XL U181 ( .A0(n209), .A1(n16), .B0(n15), .Y(n206) );
  INVX1 U182 ( .A(n13), .Y(n209) );
  INVX1 U183 ( .A(n187), .Y(n186) );
  NAND2X1 U184 ( .A(n62), .B(n216), .Y(n218) );
  NOR2X1 U185 ( .A(n219), .B(n220), .Y(n217) );
  INVX1 U186 ( .A(n44), .Y(n219) );
  INVX1 U187 ( .A(n63), .Y(n144) );
  INVX1 U188 ( .A(n203), .Y(n20) );
  NAND2X1 U189 ( .A(n210), .B(n19), .Y(n13) );
  NAND2X1 U190 ( .A(n154), .B(n139), .Y(n152) );
  XOR2X1 U191 ( .A(n149), .B(n151), .Y(SUM[18]) );
  XOR2X1 U192 ( .A(n94), .B(n96), .Y(SUM[24]) );
  NOR2BX1 U193 ( .AN(n93), .B(n97), .Y(n96) );
  XOR2X1 U194 ( .A(n184), .B(n185), .Y(SUM[14]) );
  XOR2X1 U195 ( .A(n187), .B(n188), .Y(SUM[13]) );
  NOR2BX1 U196 ( .AN(n164), .B(n11), .Y(n188) );
  XOR2X1 U197 ( .A(n128), .B(n155), .Y(SUM[16]) );
  NOR2BX1 U198 ( .AN(n139), .B(n156), .Y(n155) );
  XOR2X1 U199 ( .A(n204), .B(n205), .Y(SUM[11]) );
  INVX1 U200 ( .A(n200), .Y(n207) );
  XOR2X1 U201 ( .A(n146), .B(n147), .Y(SUM[19]) );
  INVX1 U202 ( .A(n141), .Y(n150) );
  XOR2X1 U203 ( .A(n152), .B(n153), .Y(SUM[17]) );
  XOR2X1 U204 ( .A(n116), .B(n117), .Y(SUM[22]) );
  XOR2X1 U205 ( .A(n119), .B(n120), .Y(SUM[21]) );
  XOR2X1 U206 ( .A(n121), .B(n123), .Y(SUM[20]) );
  NOR2BX1 U207 ( .AN(n106), .B(n124), .Y(n123) );
  INVX1 U208 ( .A(n122), .Y(n124) );
  INVX1 U209 ( .A(n76), .Y(n75) );
  OAI21XL U210 ( .A0(n12), .A1(n36), .B0(n37), .Y(n34) );
  OAI21XL U211 ( .A0(n31), .A1(n32), .B0(n33), .Y(n28) );
  INVX1 U212 ( .A(n34), .Y(n31) );
  INVX1 U213 ( .A(n178), .Y(n189) );
  NOR2BX1 U214 ( .AN(n27), .B(n26), .Y(n29) );
  OAI21XL U215 ( .A0(n25), .A1(n26), .B0(n27), .Y(n21) );
  INVX1 U216 ( .A(n28), .Y(n25) );
  AND2X2 U217 ( .A(n23), .B(n24), .Y(n22) );
  INVX1 U218 ( .A(n62), .Y(n43) );
  NOR2BX1 U219 ( .AN(n37), .B(n12), .Y(n38) );
  NOR2BX1 U220 ( .AN(n33), .B(n32), .Y(n35) );
  NOR2BX1 U221 ( .AN(n44), .B(n43), .Y(n61) );
  OAI21XL U222 ( .A0(n42), .A1(n43), .B0(n44), .Y(n39) );
  INVX1 U223 ( .A(n45), .Y(n42) );
  OAI2BB1X1 U224 ( .A0N(n63), .A1N(n64), .B0(n65), .Y(n45) );
  OR2X2 U225 ( .A(A[10]), .B(B[10]), .Y(n197) );
  NAND2X1 U226 ( .A(B[9]), .B(A[9]), .Y(n15) );
  OR2X2 U227 ( .A(A[14]), .B(B[14]), .Y(n179) );
  OR2X2 U228 ( .A(A[18]), .B(B[18]), .Y(n148) );
  OR2X2 U229 ( .A(A[17]), .B(B[17]), .Y(n133) );
  OR2X2 U230 ( .A(A[5]), .B(B[5]), .Y(n213) );
  OR2X2 U231 ( .A(A[9]), .B(B[9]), .Y(n198) );
  OR2X2 U232 ( .A(A[22]), .B(B[22]), .Y(n111) );
  OR2X2 U233 ( .A(A[21]), .B(B[21]), .Y(n118) );
  NAND2X1 U234 ( .A(B[20]), .B(A[20]), .Y(n106) );
  NAND2X1 U235 ( .A(B[16]), .B(A[16]), .Y(n139) );
  OR2X2 U236 ( .A(A[29]), .B(B[29]), .Y(n54) );
  OR2X2 U237 ( .A(A[16]), .B(B[16]), .Y(n132) );
  OR2X2 U238 ( .A(A[28]), .B(B[28]), .Y(n60) );
  OAI21XL U239 ( .A0(n144), .A1(n145), .B0(n65), .Y(n220) );
  OR2X2 U240 ( .A(A[25]), .B(B[25]), .Y(n90) );
  OR2X2 U241 ( .A(A[24]), .B(B[24]), .Y(n95) );
  OR2X2 U242 ( .A(A[1]), .B(B[1]), .Y(n63) );
  XOR2X1 U243 ( .A(n206), .B(n208), .Y(SUM[10]) );
  NAND2X1 U244 ( .A(B[0]), .B(A[0]), .Y(n145) );
  XOR2X1 U245 ( .A(n64), .B(n143), .Y(SUM[1]) );
  XOR2X1 U246 ( .A(n45), .B(n61), .Y(SUM[2]) );
  XOR2X1 U247 ( .A(n39), .B(n40), .Y(SUM[3]) );
  XOR2X1 U248 ( .A(n174), .B(n38), .Y(SUM[4]) );
  XOR2X1 U249 ( .A(n34), .B(n35), .Y(SUM[5]) );
  XOR2X1 U250 ( .A(n28), .B(n29), .Y(SUM[6]) );
  XOR2X1 U251 ( .A(n21), .B(n22), .Y(SUM[7]) );
  XOR2X1 U252 ( .A(n17), .B(n18), .Y(SUM[8]) );
  XOR2X1 U253 ( .A(n13), .B(n14), .Y(SUM[9]) );
  XNOR2X1 U254 ( .A(B[31]), .B(A[31]), .Y(n46) );
endmodule


module message_schedule_DW01_add_22 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n228, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227;

  CLKINVX3 U2 ( .A(n224), .Y(n43) );
  NAND2X2 U3 ( .A(n36), .B(n37), .Y(n34) );
  NAND2X2 U4 ( .A(n222), .B(n223), .Y(n171) );
  OAI21X1 U5 ( .A0(n155), .A1(n156), .B0(n157), .Y(n154) );
  NAND2X2 U6 ( .A(B[13]), .B(A[13]), .Y(n162) );
  NAND2X2 U7 ( .A(B[8]), .B(A[8]), .Y(n22) );
  XOR2X2 U8 ( .A(n141), .B(n142), .Y(SUM[19]) );
  BUFX4 U9 ( .A(n228), .Y(SUM[5]) );
  NOR2X2 U10 ( .A(n12), .B(n7), .Y(n208) );
  NOR2X2 U11 ( .A(n7), .B(n214), .Y(n4) );
  NOR2X4 U12 ( .A(A[9]), .B(B[9]), .Y(n7) );
  NOR2X2 U13 ( .A(n43), .B(n13), .Y(n223) );
  NOR2X1 U14 ( .A(n11), .B(n30), .Y(n227) );
  AOI2BB1X2 U15 ( .A0N(n11), .A1N(n28), .B0(n221), .Y(n220) );
  NOR2X2 U16 ( .A(n163), .B(n181), .Y(n177) );
  OAI21XL U17 ( .A0(n98), .A1(n109), .B0(n110), .Y(n108) );
  NOR2X1 U18 ( .A(n176), .B(n10), .Y(n201) );
  INVX1 U19 ( .A(n116), .Y(n98) );
  INVX1 U20 ( .A(n107), .Y(n99) );
  INVX2 U21 ( .A(n212), .Y(n211) );
  OR2X2 U22 ( .A(A[3]), .B(B[3]), .Y(n224) );
  OAI21XL U23 ( .A0(n135), .A1(n136), .B0(n137), .Y(n134) );
  OR2X2 U24 ( .A(A[6]), .B(B[6]), .Y(n26) );
  NOR2X2 U25 ( .A(A[7]), .B(B[7]), .Y(n11) );
  INVX1 U26 ( .A(n9), .Y(n2) );
  INVX4 U27 ( .A(n26), .Y(n30) );
  NAND2X2 U28 ( .A(n93), .B(n94), .Y(n89) );
  AOI21X1 U29 ( .A0(n173), .A1(n174), .B0(n175), .Y(n151) );
  NAND2X1 U30 ( .A(n62), .B(n63), .Y(n56) );
  OAI21XL U31 ( .A0(n163), .A1(n190), .B0(n162), .Y(n188) );
  NAND2X2 U32 ( .A(n3), .B(n205), .Y(n209) );
  NOR2BX1 U33 ( .AN(n60), .B(n139), .Y(n138) );
  NAND2X1 U34 ( .A(n50), .B(n51), .Y(n49) );
  XOR2X2 U35 ( .A(n50), .B(n52), .Y(SUM[30]) );
  INVX1 U36 ( .A(n167), .Y(n200) );
  INVX1 U37 ( .A(n128), .Y(n135) );
  INVX4 U38 ( .A(n20), .Y(n215) );
  NOR3X2 U39 ( .A(n176), .B(n166), .C(n10), .Y(n175) );
  NAND2X4 U40 ( .A(n177), .B(n178), .Y(n166) );
  OAI2BB1X1 U41 ( .A0N(n145), .A1N(n124), .B0(n133), .Y(n141) );
  OAI2BB1X2 U42 ( .A0N(n147), .A1N(n128), .B0(n137), .Y(n145) );
  XOR2X2 U43 ( .A(n182), .B(n183), .Y(SUM[15]) );
  XOR2X2 U44 ( .A(n188), .B(n189), .Y(SUM[14]) );
  NOR2BXL U45 ( .AN(n42), .B(n43), .Y(n41) );
  NOR2X1 U46 ( .A(n166), .B(n167), .Y(n169) );
  XOR2X2 U47 ( .A(n27), .B(n29), .Y(SUM[6]) );
  OAI2BB1X2 U48 ( .A0N(n32), .A1N(n2), .B0(n31), .Y(n27) );
  NAND2X4 U49 ( .A(n121), .B(n122), .Y(n97) );
  NAND4BX4 U50 ( .AN(n123), .B(n124), .C(n125), .D(n126), .Y(n122) );
  OAI2BB1X4 U51 ( .A0N(n198), .A1N(n36), .B0(n199), .Y(n192) );
  XOR2X4 U52 ( .A(n82), .B(n83), .Y(SUM[27]) );
  OAI21X4 U53 ( .A0(n84), .A1(n74), .B0(n73), .Y(n82) );
  INVX4 U54 ( .A(n85), .Y(n84) );
  NAND3X2 U55 ( .A(n95), .B(n96), .C(n97), .Y(n94) );
  NOR2X2 U56 ( .A(n167), .B(n166), .Y(n173) );
  NAND3BX2 U57 ( .AN(n165), .B(n168), .C(n169), .Y(n152) );
  NAND2X2 U58 ( .A(B[1]), .B(A[1]), .Y(n60) );
  INVX4 U59 ( .A(n17), .Y(n214) );
  NOR2BXL U60 ( .AN(n19), .B(n7), .Y(n18) );
  OAI2BB1X4 U61 ( .A0N(n195), .A1N(n192), .B0(n191), .Y(n187) );
  NOR2X1 U62 ( .A(n7), .B(n8), .Y(n202) );
  NOR2BXL U63 ( .AN(n31), .B(n9), .Y(n33) );
  AOI21X2 U64 ( .A0(n31), .A1(n35), .B0(n9), .Y(n218) );
  NAND2X2 U65 ( .A(B[5]), .B(A[5]), .Y(n31) );
  XOR2X4 U66 ( .A(n23), .B(n24), .Y(SUM[7]) );
  NOR2X4 U67 ( .A(A[10]), .B(B[10]), .Y(n8) );
  OAI2BB1X4 U68 ( .A0N(n127), .A1N(n126), .B0(n136), .Y(n147) );
  NAND3X4 U69 ( .A(n151), .B(n152), .C(n153), .Y(n126) );
  AOI21X2 U70 ( .A0(n161), .A1(n162), .B0(n163), .Y(n160) );
  INVX2 U71 ( .A(n186), .Y(n163) );
  NOR2X2 U72 ( .A(A[2]), .B(B[2]), .Y(n13) );
  INVX2 U73 ( .A(n58), .Y(n139) );
  OAI21X4 U74 ( .A0(n16), .A1(n54), .B0(n55), .Y(n50) );
  AOI21X4 U75 ( .A0(n202), .A1(n203), .B0(n204), .Y(n176) );
  NAND2X2 U76 ( .A(n226), .B(n227), .Y(n165) );
  XOR2X2 U77 ( .A(n111), .B(n112), .Y(SUM[23]) );
  OAI21X2 U78 ( .A0(n113), .A1(n99), .B0(n106), .Y(n111) );
  NAND2X2 U79 ( .A(n19), .B(n22), .Y(n203) );
  CLKINVX2 U80 ( .A(n19), .Y(n5) );
  NAND2X1 U81 ( .A(B[9]), .B(A[9]), .Y(n19) );
  NAND2X2 U82 ( .A(n207), .B(n208), .Y(n167) );
  NAND2X2 U83 ( .A(n34), .B(n35), .Y(n32) );
  NOR2X2 U84 ( .A(n9), .B(n39), .Y(n226) );
  XOR2X2 U85 ( .A(n212), .B(n213), .Y(SUM[10]) );
  NAND2XL U86 ( .A(B[7]), .B(A[7]), .Y(n25) );
  OR2X1 U87 ( .A(A[16]), .B(B[16]), .Y(n127) );
  NAND2XL U88 ( .A(B[18]), .B(A[18]), .Y(n133) );
  NOR2X2 U89 ( .A(A[5]), .B(B[5]), .Y(n9) );
  OR2X4 U90 ( .A(n211), .B(n8), .Y(n3) );
  NAND2X2 U91 ( .A(B[10]), .B(A[10]), .Y(n205) );
  XOR2X4 U92 ( .A(n209), .B(n210), .Y(SUM[11]) );
  OR2X2 U93 ( .A(n4), .B(n5), .Y(n212) );
  OAI2BB1X4 U94 ( .A0N(n218), .A1N(n219), .B0(n220), .Y(n174) );
  NOR2XL U95 ( .A(n11), .B(n30), .Y(n219) );
  INVX2 U96 ( .A(n195), .Y(n181) );
  NOR2X2 U97 ( .A(A[8]), .B(B[8]), .Y(n12) );
  OAI2BB1X2 U98 ( .A0N(n26), .A1N(n27), .B0(n28), .Y(n23) );
  NAND2XL U99 ( .A(B[21]), .B(A[21]), .Y(n110) );
  NAND2XL U100 ( .A(B[19]), .B(A[19]), .Y(n131) );
  NOR2X1 U101 ( .A(n179), .B(n180), .Y(n178) );
  NAND2XL U102 ( .A(n158), .B(n159), .Y(n156) );
  NOR2BX1 U103 ( .AN(n162), .B(n187), .Y(n184) );
  INVXL U104 ( .A(n187), .Y(n190) );
  INVXL U105 ( .A(n191), .Y(n196) );
  NOR2BX1 U106 ( .AN(n35), .B(n39), .Y(n38) );
  OAI2BB1X1 U107 ( .A0N(n58), .A1N(n59), .B0(n60), .Y(n46) );
  INVX1 U108 ( .A(n159), .Y(n179) );
  NAND2X4 U109 ( .A(B[0]), .B(A[0]), .Y(n140) );
  NAND2X1 U110 ( .A(B[6]), .B(A[6]), .Y(n28) );
  OR2X2 U111 ( .A(A[12]), .B(B[12]), .Y(n195) );
  NAND2XL U112 ( .A(B[14]), .B(A[14]), .Y(n164) );
  NAND2X1 U113 ( .A(B[16]), .B(A[16]), .Y(n136) );
  OR2X2 U114 ( .A(A[18]), .B(B[18]), .Y(n124) );
  OAI2BB1X2 U115 ( .A0N(n216), .A1N(n36), .B0(n217), .Y(n20) );
  CLKINVX3 U116 ( .A(n165), .Y(n216) );
  INVX2 U117 ( .A(n174), .Y(n217) );
  NAND3BX4 U118 ( .AN(n172), .B(n42), .C(n171), .Y(n36) );
  NOR2BXL U119 ( .AN(n28), .B(n30), .Y(n29) );
  AOI21X2 U120 ( .A0(n60), .A1(n140), .B0(n139), .Y(n222) );
  INVX2 U121 ( .A(n37), .Y(n39) );
  OAI21X4 U122 ( .A0(n12), .A1(n215), .B0(n22), .Y(n17) );
  OAI21X2 U123 ( .A0(n119), .A1(n14), .B0(n109), .Y(n117) );
  AOI21XL U124 ( .A0(n192), .A1(n195), .B0(n196), .Y(n194) );
  INVXL U125 ( .A(n125), .Y(n143) );
  NOR2BXL U126 ( .AN(n104), .B(n100), .Y(n112) );
  NOR2BXL U127 ( .AN(n164), .B(n180), .Y(n189) );
  OAI2BB1X2 U128 ( .A0N(n81), .A1N(n87), .B0(n78), .Y(n85) );
  OAI2BB1X2 U129 ( .A0N(n116), .A1N(n117), .B0(n110), .Y(n114) );
  NAND2X2 U130 ( .A(n89), .B(n90), .Y(n68) );
  NOR2BX1 U131 ( .AN(n164), .B(n160), .Y(n155) );
  NOR2BXL U132 ( .AN(n42), .B(n172), .Y(n170) );
  NOR2BX1 U133 ( .AN(n79), .B(n71), .Y(n70) );
  NOR2BXL U134 ( .AN(n78), .B(n76), .Y(n88) );
  NOR2BXL U135 ( .AN(n191), .B(n181), .Y(n197) );
  NAND2XL U136 ( .A(n127), .B(n128), .Y(n123) );
  INVXL U137 ( .A(n90), .Y(n92) );
  NAND2X2 U138 ( .A(B[2]), .B(A[2]), .Y(n45) );
  OR2X4 U139 ( .A(A[1]), .B(B[1]), .Y(n58) );
  NOR2X2 U140 ( .A(A[11]), .B(B[11]), .Y(n10) );
  NAND2XL U141 ( .A(B[3]), .B(A[3]), .Y(n42) );
  NAND2XL U142 ( .A(B[11]), .B(A[11]), .Y(n206) );
  OR2X4 U143 ( .A(A[13]), .B(B[13]), .Y(n186) );
  OR2X4 U144 ( .A(A[14]), .B(B[14]), .Y(n158) );
  NAND2XL U145 ( .A(B[12]), .B(A[12]), .Y(n191) );
  NAND2XL U146 ( .A(B[17]), .B(A[17]), .Y(n137) );
  NAND2XL U147 ( .A(B[15]), .B(A[15]), .Y(n157) );
  NOR2XL U148 ( .A(A[20]), .B(B[20]), .Y(n14) );
  NOR2BX1 U149 ( .AN(n140), .B(n6), .Y(SUM[0]) );
  NOR2XL U150 ( .A(A[0]), .B(B[0]), .Y(n6) );
  NAND2XL U151 ( .A(B[24]), .B(A[24]), .Y(n77) );
  NAND2XL U152 ( .A(B[22]), .B(A[22]), .Y(n106) );
  NAND2XL U153 ( .A(B[25]), .B(A[25]), .Y(n78) );
  NAND2XL U154 ( .A(B[23]), .B(A[23]), .Y(n104) );
  INVX1 U155 ( .A(n154), .Y(n153) );
  NOR2X1 U156 ( .A(n99), .B(n100), .Y(n95) );
  NOR2X1 U157 ( .A(n8), .B(n10), .Y(n207) );
  NAND2X1 U158 ( .A(n205), .B(n206), .Y(n204) );
  XOR2X1 U159 ( .A(n85), .B(n86), .Y(SUM[26]) );
  NOR2BX1 U160 ( .AN(n73), .B(n74), .Y(n86) );
  INVX1 U161 ( .A(n97), .Y(n119) );
  AOI21X1 U162 ( .A0(n200), .A1(n174), .B0(n201), .Y(n199) );
  NOR2X1 U163 ( .A(n167), .B(n165), .Y(n198) );
  INVX1 U164 ( .A(n158), .Y(n180) );
  AOI21X1 U165 ( .A0(n129), .A1(n125), .B0(n130), .Y(n121) );
  INVX1 U166 ( .A(n131), .Y(n130) );
  NOR2BX1 U167 ( .AN(n205), .B(n8), .Y(n213) );
  XOR2X1 U168 ( .A(n17), .B(n18), .Y(SUM[9]) );
  XOR2X1 U169 ( .A(n145), .B(n146), .Y(SUM[18]) );
  NOR2BX1 U170 ( .AN(n133), .B(n144), .Y(n146) );
  XOR2X1 U171 ( .A(n117), .B(n118), .Y(SUM[21]) );
  NOR2BX1 U172 ( .AN(n110), .B(n98), .Y(n118) );
  NOR2BX1 U173 ( .AN(n206), .B(n10), .Y(n210) );
  INVX1 U174 ( .A(n114), .Y(n113) );
  NOR2BX1 U175 ( .AN(n79), .B(n15), .Y(n83) );
  NOR2BX1 U176 ( .AN(n131), .B(n143), .Y(n142) );
  NOR2BX1 U177 ( .AN(n157), .B(n179), .Y(n183) );
  OAI21XL U178 ( .A0(n184), .A1(n185), .B0(n164), .Y(n182) );
  NAND2X1 U179 ( .A(n186), .B(n158), .Y(n185) );
  XOR2X1 U180 ( .A(n193), .B(n194), .Y(SUM[13]) );
  NAND2X1 U181 ( .A(n186), .B(n162), .Y(n193) );
  NOR2BX1 U182 ( .AN(n25), .B(n11), .Y(n24) );
  XOR2X1 U183 ( .A(n32), .B(n33), .Y(n228) );
  XOR2X1 U184 ( .A(n147), .B(n148), .Y(SUM[17]) );
  NOR2BX1 U185 ( .AN(n137), .B(n135), .Y(n148) );
  XOR2X1 U186 ( .A(n114), .B(n115), .Y(SUM[22]) );
  NOR2BX1 U187 ( .AN(n106), .B(n99), .Y(n115) );
  AOI21X1 U188 ( .A0(n101), .A1(n102), .B0(n103), .Y(n93) );
  INVX1 U189 ( .A(n104), .Y(n103) );
  INVX1 U190 ( .A(n225), .Y(n172) );
  NAND2BX1 U191 ( .AN(n45), .B(n224), .Y(n225) );
  NAND2X1 U192 ( .A(n68), .B(n77), .Y(n87) );
  INVX1 U193 ( .A(n25), .Y(n221) );
  NAND2X1 U194 ( .A(n170), .B(n171), .Y(n168) );
  NOR2BX1 U195 ( .AN(n48), .B(n53), .Y(n52) );
  INVX1 U196 ( .A(n51), .Y(n53) );
  INVX1 U197 ( .A(n56), .Y(n54) );
  OAI21XL U198 ( .A0(n68), .A1(n69), .B0(n70), .Y(n64) );
  NAND3BX1 U199 ( .AN(n15), .B(n80), .C(n81), .Y(n69) );
  XOR2X1 U200 ( .A(n87), .B(n88), .Y(SUM[25]) );
  XOR2X1 U201 ( .A(n89), .B(n91), .Y(SUM[24]) );
  NOR2BX1 U202 ( .AN(n77), .B(n92), .Y(n91) );
  XOR2X1 U203 ( .A(n56), .B(n61), .Y(SUM[29]) );
  NOR2BX1 U204 ( .AN(n55), .B(n16), .Y(n61) );
  XOR2X1 U205 ( .A(n36), .B(n38), .Y(SUM[4]) );
  XOR2X1 U206 ( .A(n126), .B(n149), .Y(SUM[16]) );
  NOR2BX1 U207 ( .AN(n136), .B(n150), .Y(n149) );
  INVX1 U208 ( .A(n127), .Y(n150) );
  XOR2X1 U209 ( .A(n64), .B(n66), .Y(SUM[28]) );
  NOR2BX1 U210 ( .AN(n63), .B(n67), .Y(n66) );
  INVX1 U211 ( .A(n65), .Y(n67) );
  XOR2X1 U212 ( .A(n192), .B(n197), .Y(SUM[12]) );
  XOR2X1 U213 ( .A(n97), .B(n120), .Y(SUM[20]) );
  NOR2BX1 U214 ( .AN(n109), .B(n14), .Y(n120) );
  XOR2X1 U215 ( .A(n40), .B(n41), .Y(SUM[3]) );
  OAI21XL U216 ( .A0(n44), .A1(n13), .B0(n45), .Y(n40) );
  INVX1 U217 ( .A(n46), .Y(n44) );
  XOR2X1 U218 ( .A(n59), .B(n138), .Y(SUM[1]) );
  XOR2X1 U219 ( .A(n46), .B(n57), .Y(SUM[2]) );
  NOR2BX1 U220 ( .AN(n45), .B(n13), .Y(n57) );
  XOR2X1 U221 ( .A(n20), .B(n21), .Y(SUM[8]) );
  NOR2BX1 U222 ( .AN(n22), .B(n12), .Y(n21) );
  NOR2X1 U223 ( .A(n98), .B(n14), .Y(n96) );
  INVX1 U224 ( .A(n140), .Y(n59) );
  NAND2X1 U225 ( .A(n105), .B(n106), .Y(n101) );
  NAND2X1 U226 ( .A(n107), .B(n108), .Y(n105) );
  NAND2X1 U227 ( .A(n132), .B(n133), .Y(n129) );
  NAND2X1 U228 ( .A(n124), .B(n134), .Y(n132) );
  NAND2X1 U229 ( .A(n64), .B(n65), .Y(n62) );
  INVX1 U230 ( .A(n80), .Y(n74) );
  INVX1 U231 ( .A(n124), .Y(n144) );
  INVX1 U232 ( .A(n81), .Y(n76) );
  INVX1 U233 ( .A(n102), .Y(n100) );
  AOI21X1 U234 ( .A0(n72), .A1(n73), .B0(n15), .Y(n71) );
  NAND2BX1 U235 ( .AN(n74), .B(n75), .Y(n72) );
  OAI21XL U236 ( .A0(n76), .A1(n77), .B0(n78), .Y(n75) );
  NAND2X1 U237 ( .A(B[4]), .B(A[4]), .Y(n35) );
  NAND2X1 U238 ( .A(B[12]), .B(A[12]), .Y(n161) );
  OR2X2 U239 ( .A(A[15]), .B(B[15]), .Y(n159) );
  OR2X2 U240 ( .A(A[4]), .B(B[4]), .Y(n37) );
  OR2X2 U241 ( .A(A[19]), .B(B[19]), .Y(n125) );
  OR2X2 U242 ( .A(A[22]), .B(B[22]), .Y(n107) );
  OR2X2 U243 ( .A(A[17]), .B(B[17]), .Y(n128) );
  OR2X2 U244 ( .A(A[21]), .B(B[21]), .Y(n116) );
  NAND2X1 U245 ( .A(B[20]), .B(A[20]), .Y(n109) );
  OR2X2 U246 ( .A(A[25]), .B(B[25]), .Y(n81) );
  OR2X2 U247 ( .A(A[23]), .B(B[23]), .Y(n102) );
  OR2X2 U248 ( .A(A[24]), .B(B[24]), .Y(n90) );
  OR2X2 U249 ( .A(A[26]), .B(B[26]), .Y(n80) );
  NAND2X1 U250 ( .A(B[26]), .B(A[26]), .Y(n73) );
  NAND2X1 U251 ( .A(B[28]), .B(A[28]), .Y(n63) );
  NAND2X1 U252 ( .A(B[27]), .B(A[27]), .Y(n79) );
  OR2X2 U253 ( .A(A[28]), .B(B[28]), .Y(n65) );
  NOR2X1 U254 ( .A(A[27]), .B(B[27]), .Y(n15) );
  NAND2X1 U255 ( .A(B[30]), .B(A[30]), .Y(n48) );
  NAND2X1 U256 ( .A(B[29]), .B(A[29]), .Y(n55) );
  OR2X2 U257 ( .A(A[30]), .B(B[30]), .Y(n51) );
  NOR2X1 U258 ( .A(A[29]), .B(B[29]), .Y(n16) );
  XOR3X2 U259 ( .A(B[31]), .B(A[31]), .C(n47), .Y(SUM[31]) );
  NAND2X1 U260 ( .A(n48), .B(n49), .Y(n47) );
endmodule


module message_schedule_DW01_add_23 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207;

  NOR2X2 U2 ( .A(A[12]), .B(B[12]), .Y(n16) );
  NAND2X1 U3 ( .A(n94), .B(n103), .Y(n114) );
  NOR2X2 U4 ( .A(A[8]), .B(B[8]), .Y(n15) );
  AOI21X2 U5 ( .A0(n123), .A1(n142), .B0(n143), .Y(n141) );
  OR2X4 U6 ( .A(A[6]), .B(B[6]), .Y(n29) );
  AOI21X2 U7 ( .A0(n200), .A1(n201), .B0(n202), .Y(n199) );
  OAI21XL U8 ( .A0(n7), .A1(n31), .B0(n28), .Y(n202) );
  NAND2X1 U9 ( .A(B[10]), .B(A[10]), .Y(n188) );
  AOI21X2 U10 ( .A0(n64), .A1(n65), .B0(n66), .Y(n56) );
  NAND2X1 U11 ( .A(B[5]), .B(A[5]), .Y(n35) );
  AOI21X2 U12 ( .A0(n22), .A1(n25), .B0(n13), .Y(n186) );
  NOR2X2 U13 ( .A(n13), .B(n14), .Y(n190) );
  NOR2BXL U14 ( .AN(n188), .B(n13), .Y(n196) );
  OAI21X2 U15 ( .A0(n194), .A1(n13), .B0(n188), .Y(n192) );
  NOR2X2 U16 ( .A(A[10]), .B(B[10]), .Y(n13) );
  NOR2X1 U17 ( .A(n12), .B(n14), .Y(n185) );
  OAI21X1 U18 ( .A0(n188), .A1(n14), .B0(n189), .Y(n187) );
  NAND2X1 U19 ( .A(B[13]), .B(A[13]), .Y(n164) );
  OAI21XL U20 ( .A0(n102), .A1(n103), .B0(n104), .Y(n101) );
  OAI21XL U21 ( .A0(n134), .A1(n135), .B0(n136), .Y(n133) );
  NAND2X1 U22 ( .A(n190), .B(n191), .Y(n156) );
  INVX1 U23 ( .A(n29), .Y(n33) );
  OR2X2 U24 ( .A(A[18]), .B(B[18]), .Y(n123) );
  INVX1 U25 ( .A(n154), .Y(n198) );
  INVX1 U26 ( .A(n20), .Y(n197) );
  INVX1 U27 ( .A(n127), .Y(n134) );
  XOR2X1 U28 ( .A(n178), .B(n179), .Y(SUM[13]) );
  XOR2X1 U29 ( .A(n182), .B(n183), .Y(SUM[12]) );
  XOR2X1 U30 ( .A(n20), .B(n21), .Y(SUM[9]) );
  INVX2 U31 ( .A(n111), .Y(n110) );
  XOR2X1 U32 ( .A(n111), .B(n112), .Y(SUM[22]) );
  XOR2X1 U33 ( .A(n175), .B(n176), .Y(SUM[14]) );
  INVX1 U34 ( .A(n199), .Y(n167) );
  OR2X2 U35 ( .A(n16), .B(n180), .Y(n2) );
  NOR2BXL U36 ( .AN(n48), .B(n10), .Y(n59) );
  OAI21XL U37 ( .A0(n47), .A1(n10), .B0(n48), .Y(n44) );
  NOR2X2 U38 ( .A(n9), .B(n10), .Y(n204) );
  NOR2BXL U39 ( .AN(n28), .B(n7), .Y(n27) );
  NOR2X2 U40 ( .A(n7), .B(n33), .Y(n201) );
  NOR2X2 U41 ( .A(n7), .B(n33), .Y(n207) );
  OAI2BB1X1 U42 ( .A0N(n146), .A1N(n127), .B0(n136), .Y(n142) );
  NAND2X2 U43 ( .A(B[0]), .B(A[0]), .Y(n139) );
  XOR2X2 U44 ( .A(n85), .B(n86), .Y(SUM[26]) );
  NAND2X1 U45 ( .A(B[3]), .B(A[3]), .Y(n46) );
  OAI21X1 U46 ( .A0(n68), .A1(n69), .B0(n70), .Y(n64) );
  NAND2X4 U47 ( .A(n1), .B(n91), .Y(n68) );
  OAI21X4 U48 ( .A0(n9), .A1(n48), .B0(n46), .Y(n205) );
  NOR2X2 U49 ( .A(A[3]), .B(B[3]), .Y(n9) );
  XOR2X4 U50 ( .A(n82), .B(n83), .Y(SUM[27]) );
  OAI21X4 U51 ( .A0(n84), .A1(n74), .B0(n73), .Y(n82) );
  INVX4 U52 ( .A(n114), .Y(n113) );
  OAI21X4 U53 ( .A0(n113), .A1(n102), .B0(n104), .Y(n111) );
  XOR2X2 U54 ( .A(n108), .B(n109), .Y(SUM[23]) );
  XOR2X4 U55 ( .A(n172), .B(n173), .Y(SUM[15]) );
  NOR4X1 U56 ( .A(n169), .B(n154), .C(n155), .D(n156), .Y(n151) );
  NOR2BXL U57 ( .AN(n189), .B(n14), .Y(n193) );
  NOR2X2 U58 ( .A(A[11]), .B(B[11]), .Y(n14) );
  NAND3BX4 U59 ( .AN(n151), .B(n153), .C(n152), .Y(n125) );
  NAND2X2 U60 ( .A(n170), .B(n171), .Y(n155) );
  BUFX4 U61 ( .A(n90), .Y(n1) );
  OAI21X1 U62 ( .A0(n94), .A1(n95), .B0(n96), .Y(n90) );
  OAI21X2 U63 ( .A0(n15), .A1(n184), .B0(n25), .Y(n20) );
  OAI21X4 U64 ( .A0(n177), .A1(n11), .B0(n164), .Y(n175) );
  OAI21X2 U65 ( .A0(n34), .A1(n8), .B0(n35), .Y(n30) );
  NOR2X4 U66 ( .A(n8), .B(n43), .Y(n206) );
  AOI21X2 U67 ( .A0(n35), .A1(n39), .B0(n8), .Y(n200) );
  NOR2X2 U68 ( .A(A[5]), .B(B[5]), .Y(n8) );
  CLKINVX4 U69 ( .A(n169), .Y(n40) );
  AOI21X2 U70 ( .A0(n203), .A1(n204), .B0(n205), .Y(n169) );
  NOR2X2 U71 ( .A(A[2]), .B(B[2]), .Y(n10) );
  NAND2X4 U72 ( .A(n2), .B(n181), .Y(n178) );
  INVX1 U73 ( .A(n182), .Y(n180) );
  INVX4 U74 ( .A(n178), .Y(n177) );
  NAND2X1 U75 ( .A(B[1]), .B(A[1]), .Y(n62) );
  OR2XL U76 ( .A(n184), .B(n156), .Y(n3) );
  NAND2X2 U77 ( .A(n3), .B(n168), .Y(n182) );
  INVX4 U78 ( .A(n23), .Y(n184) );
  AOI21X2 U79 ( .A0(n185), .A1(n186), .B0(n187), .Y(n168) );
  NAND2X2 U80 ( .A(B[2]), .B(A[2]), .Y(n48) );
  NOR2X2 U81 ( .A(A[9]), .B(B[9]), .Y(n12) );
  NAND2XL U82 ( .A(B[9]), .B(A[9]), .Y(n22) );
  NAND2X1 U83 ( .A(n38), .B(n39), .Y(n36) );
  NOR2X2 U84 ( .A(A[13]), .B(B[13]), .Y(n11) );
  NAND2XL U85 ( .A(B[8]), .B(A[8]), .Y(n25) );
  INVX1 U86 ( .A(n195), .Y(n194) );
  OAI21X1 U87 ( .A0(n12), .A1(n197), .B0(n22), .Y(n195) );
  INVX1 U88 ( .A(n60), .Y(n138) );
  NAND3BXL U89 ( .AN(n18), .B(n106), .C(n107), .Y(n95) );
  NOR2BX1 U90 ( .AN(n73), .B(n74), .Y(n86) );
  NOR2X1 U91 ( .A(n15), .B(n12), .Y(n191) );
  INVX1 U92 ( .A(n41), .Y(n43) );
  OR2X1 U93 ( .A(A[16]), .B(B[16]), .Y(n126) );
  OAI2BB1X2 U94 ( .A0N(n198), .A1N(n40), .B0(n199), .Y(n23) );
  NOR2BXL U95 ( .AN(n165), .B(n17), .Y(n173) );
  NAND2XL U96 ( .A(n40), .B(n41), .Y(n38) );
  NOR2BX1 U97 ( .AN(n105), .B(n97), .Y(n96) );
  NOR2BXL U98 ( .AN(n99), .B(n100), .Y(n112) );
  NOR2BXL U99 ( .AN(n181), .B(n16), .Y(n183) );
  NOR2BXL U100 ( .AN(n35), .B(n8), .Y(n37) );
  NOR2BXL U101 ( .AN(n25), .B(n15), .Y(n24) );
  NOR2BXL U102 ( .AN(n105), .B(n18), .Y(n109) );
  OAI21X1 U103 ( .A0(n110), .A1(n100), .B0(n99), .Y(n108) );
  INVX2 U104 ( .A(n174), .Y(n161) );
  NAND2XL U105 ( .A(n125), .B(n126), .Y(n148) );
  NAND2X2 U106 ( .A(n116), .B(n117), .Y(n94) );
  NAND2X2 U107 ( .A(n87), .B(n78), .Y(n85) );
  XOR2X2 U108 ( .A(n53), .B(n6), .Y(SUM[30]) );
  NOR2BX1 U109 ( .AN(n79), .B(n71), .Y(n70) );
  OAI21X1 U110 ( .A0(n55), .A1(n56), .B0(n57), .Y(n53) );
  NOR2BXL U111 ( .AN(n104), .B(n102), .Y(n115) );
  NOR2BXL U112 ( .AN(n62), .B(n138), .Y(n137) );
  NAND2XL U113 ( .A(n53), .B(n54), .Y(n52) );
  NAND2XL U114 ( .A(n126), .B(n127), .Y(n122) );
  XOR2XL U115 ( .A(n63), .B(n56), .Y(SUM[29]) );
  XNOR2X1 U116 ( .A(n64), .B(n4), .Y(SUM[28]) );
  NAND2X1 U117 ( .A(n67), .B(n65), .Y(n4) );
  NOR2X2 U118 ( .A(A[7]), .B(B[7]), .Y(n7) );
  NAND2XL U119 ( .A(B[7]), .B(A[7]), .Y(n28) );
  NAND2XL U120 ( .A(B[14]), .B(A[14]), .Y(n160) );
  NAND2XL U121 ( .A(B[11]), .B(A[11]), .Y(n189) );
  NAND2BXL U122 ( .AN(n161), .B(n162), .Y(n159) );
  NAND2XL U123 ( .A(A[12]), .B(B[12]), .Y(n163) );
  NAND2XL U124 ( .A(B[17]), .B(A[17]), .Y(n136) );
  NAND2XL U125 ( .A(B[19]), .B(A[19]), .Y(n130) );
  NAND2XL U126 ( .A(B[12]), .B(A[12]), .Y(n181) );
  NAND2XL U127 ( .A(B[15]), .B(A[15]), .Y(n165) );
  NOR2BX1 U128 ( .AN(n139), .B(n5), .Y(SUM[0]) );
  NOR2XL U129 ( .A(A[0]), .B(B[0]), .Y(n5) );
  NAND2XL U130 ( .A(B[22]), .B(A[22]), .Y(n99) );
  NAND2XL U131 ( .A(B[21]), .B(A[21]), .Y(n104) );
  NAND2XL U132 ( .A(B[23]), .B(A[23]), .Y(n105) );
  OR2XL U133 ( .A(A[20]), .B(B[20]), .Y(n117) );
  NOR2X1 U134 ( .A(n156), .B(n155), .Y(n166) );
  AOI21X1 U135 ( .A0(n62), .A1(n139), .B0(n138), .Y(n203) );
  XOR2X1 U136 ( .A(n195), .B(n196), .Y(SUM[10]) );
  NOR2BX1 U137 ( .AN(n164), .B(n11), .Y(n179) );
  NOR2BX1 U138 ( .AN(n160), .B(n161), .Y(n176) );
  XOR2X1 U139 ( .A(n192), .B(n193), .Y(SUM[11]) );
  OAI2BB1X1 U140 ( .A0N(n174), .A1N(n175), .B0(n160), .Y(n172) );
  NAND2X1 U141 ( .A(n206), .B(n207), .Y(n154) );
  NOR2X1 U142 ( .A(n157), .B(n158), .Y(n153) );
  AOI2BB2X1 U143 ( .B0(n166), .B1(n167), .A0N(n168), .A1N(n155), .Y(n152) );
  INVX1 U144 ( .A(n36), .Y(n34) );
  XOR2X1 U145 ( .A(n88), .B(n89), .Y(SUM[25]) );
  NOR2BX1 U146 ( .AN(n78), .B(n76), .Y(n89) );
  NOR2X1 U147 ( .A(n17), .B(n161), .Y(n171) );
  NOR2X1 U148 ( .A(n11), .B(n16), .Y(n170) );
  XOR2X1 U149 ( .A(n142), .B(n144), .Y(SUM[18]) );
  NOR2BX1 U150 ( .AN(n132), .B(n145), .Y(n144) );
  INVX1 U151 ( .A(n123), .Y(n145) );
  NOR2BX1 U152 ( .AN(n22), .B(n12), .Y(n21) );
  XOR2X1 U153 ( .A(n30), .B(n32), .Y(SUM[6]) );
  NOR2BX1 U154 ( .AN(n31), .B(n33), .Y(n32) );
  XOR2X1 U155 ( .A(n40), .B(n42), .Y(SUM[4]) );
  NOR2BX1 U156 ( .AN(n39), .B(n43), .Y(n42) );
  NOR2BX1 U157 ( .AN(n79), .B(n19), .Y(n83) );
  INVX1 U158 ( .A(n85), .Y(n84) );
  XOR2X1 U159 ( .A(n140), .B(n141), .Y(SUM[19]) );
  NAND2X1 U160 ( .A(n130), .B(n124), .Y(n140) );
  INVX1 U161 ( .A(n132), .Y(n143) );
  XOR2X1 U162 ( .A(n26), .B(n27), .Y(SUM[7]) );
  OAI2BB1X1 U163 ( .A0N(n29), .A1N(n30), .B0(n31), .Y(n26) );
  XOR2X1 U164 ( .A(n36), .B(n37), .Y(SUM[5]) );
  XOR2X1 U165 ( .A(n146), .B(n147), .Y(SUM[17]) );
  NOR2BX1 U166 ( .AN(n136), .B(n134), .Y(n147) );
  XOR2X1 U167 ( .A(n23), .B(n24), .Y(SUM[8]) );
  XOR2X1 U168 ( .A(n114), .B(n115), .Y(SUM[21]) );
  NAND2X1 U169 ( .A(n120), .B(n121), .Y(n116) );
  AOI21X1 U170 ( .A0(n124), .A1(n128), .B0(n129), .Y(n120) );
  NAND4BXL U171 ( .AN(n122), .B(n123), .C(n124), .D(n125), .Y(n121) );
  INVX1 U172 ( .A(n130), .Y(n129) );
  NAND2X1 U173 ( .A(n68), .B(n77), .Y(n88) );
  NAND2X1 U174 ( .A(n148), .B(n135), .Y(n146) );
  NAND2X1 U175 ( .A(n81), .B(n88), .Y(n87) );
  NAND2X1 U176 ( .A(n131), .B(n132), .Y(n128) );
  NAND2X1 U177 ( .A(n123), .B(n133), .Y(n131) );
  AND2X2 U178 ( .A(n51), .B(n54), .Y(n6) );
  INVX1 U179 ( .A(n67), .Y(n66) );
  INVX1 U180 ( .A(n107), .Y(n102) );
  NAND3BX1 U181 ( .AN(n19), .B(n80), .C(n81), .Y(n69) );
  INVX1 U182 ( .A(n58), .Y(n55) );
  INVX1 U183 ( .A(n106), .Y(n100) );
  XOR2X1 U184 ( .A(n1), .B(n92), .Y(SUM[24]) );
  NOR2BX1 U185 ( .AN(n77), .B(n93), .Y(n92) );
  INVX1 U186 ( .A(n91), .Y(n93) );
  NAND2X1 U187 ( .A(n57), .B(n58), .Y(n63) );
  XOR2X1 U188 ( .A(n125), .B(n149), .Y(SUM[16]) );
  NOR2BX1 U189 ( .AN(n135), .B(n150), .Y(n149) );
  INVX1 U190 ( .A(n126), .Y(n150) );
  XOR2X1 U191 ( .A(n44), .B(n45), .Y(SUM[3]) );
  NOR2BX1 U192 ( .AN(n46), .B(n9), .Y(n45) );
  INVX1 U193 ( .A(n49), .Y(n47) );
  XOR2X1 U194 ( .A(n116), .B(n118), .Y(SUM[20]) );
  NOR2BX1 U195 ( .AN(n103), .B(n119), .Y(n118) );
  INVX1 U196 ( .A(n117), .Y(n119) );
  XOR2X1 U197 ( .A(n61), .B(n137), .Y(SUM[1]) );
  XOR2X1 U198 ( .A(n49), .B(n59), .Y(SUM[2]) );
  AOI21X1 U199 ( .A0(n98), .A1(n99), .B0(n18), .Y(n97) );
  NAND2BX1 U200 ( .AN(n100), .B(n101), .Y(n98) );
  OAI2BB1X1 U201 ( .A0N(n60), .A1N(n61), .B0(n62), .Y(n49) );
  INVX1 U202 ( .A(n139), .Y(n61) );
  INVX1 U203 ( .A(n165), .Y(n157) );
  NAND2X1 U204 ( .A(n51), .B(n52), .Y(n50) );
  INVX1 U205 ( .A(n80), .Y(n74) );
  INVX1 U206 ( .A(n81), .Y(n76) );
  AOI21X1 U207 ( .A0(n72), .A1(n73), .B0(n19), .Y(n71) );
  NAND2BX1 U208 ( .AN(n74), .B(n75), .Y(n72) );
  OAI21XL U209 ( .A0(n76), .A1(n77), .B0(n78), .Y(n75) );
  NAND2X1 U210 ( .A(B[4]), .B(A[4]), .Y(n39) );
  NAND2X1 U211 ( .A(B[6]), .B(A[6]), .Y(n31) );
  OR2X2 U212 ( .A(A[4]), .B(B[4]), .Y(n41) );
  XOR3X2 U213 ( .A(B[31]), .B(A[31]), .C(n50), .Y(SUM[31]) );
  OR2X2 U214 ( .A(A[1]), .B(B[1]), .Y(n60) );
  NOR2X1 U215 ( .A(A[15]), .B(B[15]), .Y(n17) );
  AOI21X1 U216 ( .A0(n159), .A1(n160), .B0(n17), .Y(n158) );
  OAI21XL U217 ( .A0(n11), .A1(n163), .B0(n164), .Y(n162) );
  OR2X2 U218 ( .A(A[17]), .B(B[17]), .Y(n127) );
  OR2X2 U219 ( .A(A[14]), .B(B[14]), .Y(n174) );
  NOR2X1 U220 ( .A(A[23]), .B(B[23]), .Y(n18) );
  NAND2X1 U221 ( .A(B[16]), .B(A[16]), .Y(n135) );
  NAND2X1 U222 ( .A(B[20]), .B(A[20]), .Y(n103) );
  OR2X2 U223 ( .A(A[19]), .B(B[19]), .Y(n124) );
  NAND2X1 U224 ( .A(B[18]), .B(A[18]), .Y(n132) );
  OR2X2 U225 ( .A(A[21]), .B(B[21]), .Y(n107) );
  OR2X2 U226 ( .A(A[22]), .B(B[22]), .Y(n106) );
  NOR2X1 U227 ( .A(A[27]), .B(B[27]), .Y(n19) );
  NAND2X1 U228 ( .A(B[24]), .B(A[24]), .Y(n77) );
  NAND2X1 U229 ( .A(B[26]), .B(A[26]), .Y(n73) );
  NAND2X1 U230 ( .A(B[25]), .B(A[25]), .Y(n78) );
  OR2X2 U231 ( .A(A[25]), .B(B[25]), .Y(n81) );
  OR2X2 U232 ( .A(A[24]), .B(B[24]), .Y(n91) );
  OR2X2 U233 ( .A(A[26]), .B(B[26]), .Y(n80) );
  NAND2X1 U234 ( .A(B[30]), .B(A[30]), .Y(n51) );
  NAND2X1 U235 ( .A(B[29]), .B(A[29]), .Y(n57) );
  NAND2X1 U236 ( .A(B[28]), .B(A[28]), .Y(n67) );
  OR2X2 U237 ( .A(A[28]), .B(B[28]), .Y(n65) );
  OR2X2 U238 ( .A(A[30]), .B(B[30]), .Y(n54) );
  NAND2X1 U239 ( .A(B[27]), .B(A[27]), .Y(n79) );
  OR2X2 U240 ( .A(A[29]), .B(B[29]), .Y(n58) );
endmodule


module message_schedule ( clk, reset, data, write_enable, inner_busy, Wt );
  input [7:0] data;
  output [31:0] Wt;
  input clk, reset, write_enable, inner_busy;
  wire   n2216, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451,
         N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462,
         N463, N464, N465, N474, N475, N476, N477, N478, N479, N480, N481,
         N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492,
         N493, N494, N495, N496, N497, N506, N507, N508, N509, N510, N511,
         N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522,
         N523, N524, N525, N526, N527, N528, N529, N538, N539, N540, N541,
         N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552,
         N553, N554, N555, N556, N557, N558, N559, N560, N561, N570, N571,
         N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582,
         N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593,
         N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612,
         N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623,
         N624, N625, N634, N635, N636, N637, N638, N639, N640, N641, N642,
         N643, N644, N645, N646, N647, N648, N649, N650, N651, N652, N653,
         N654, N655, N656, N657, N666, N667, N668, N669, N670, N671, N672,
         N673, N674, N675, N676, N677, N678, N679, N680, N681, N682, N683,
         N684, N685, N686, N687, N688, N689, N698, N699, N700, N701, N702,
         N703, N704, N705, N706, N707, N708, N709, N710, N711, N712, N713,
         N714, N715, N716, N717, N718, N719, N720, N721, N730, N731, N732,
         N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743,
         N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N762,
         N763, N764, N765, N766, N767, N768, N769, N770, N771, N772, N773,
         N774, N775, N776, N777, N778, N779, N780, N781, N782, N783, N784,
         N785, N794, N795, N796, N797, N798, N799, N800, N801, N802, N803,
         N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814,
         N815, N816, N817, N826, N827, N828, N829, N830, N831, N832, N833,
         N834, N835, N836, N837, N838, N839, N840, N841, N842, N843, N844,
         N845, N846, N847, N848, N849, N858, N859, N860, N861, N862, N863,
         N864, N865, N866, N867, N868, N869, N870, N871, N872, N873, N874,
         N875, N876, N877, N878, N879, N880, N881, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N911, N912, N913, N922, N923,
         N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934,
         N935, N936, N937, N938, N939, N940, N941, N942, N943, N944, N945,
         N1462, N1463, N1464, N1465, N1466, N1467, N1468, N2131, N2132, N2133,
         N2134, N2135, N2136, N2137, N2138, N2139, N2140, N2141, N2142, N2143,
         N2144, N2145, N2146, N2147, N2148, N2149, N2150, N2151, N2152, N2153,
         N2154, N2155, N2156, N2157, N2158, N2159, N2160, N2161, N2162, N2169,
         N2170, N2171, N2172, N2173, N2174, N2175, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1433,
         n1434, n1435, n1436, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1475, n1476, n1477, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1657, n1658, n1659, n1662, n1664, n1665, n1666, n1667, n1668,
         n1670, n1671, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1683,
         n1684, n1685, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1733, n1735, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2067, n2068, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76,
         N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62,
         N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48,
         N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34,
         N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, n49, n50, n51,
         n52, n53, n54, n55, n56, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n70, n71, n72, n74, n75, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n116, n117, n118, n119, n120, n121, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n135,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n169, n170, n172, n174, n175, n190, n545,
         n546, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1150, n1159, n1192, n1228,
         n1432, n1437, n1438, n1439, n1473, n1474, n1478, n1541, n1625, n1626,
         n1627, n1639, n1656, n1660, n1661, n1663, n1669, n1672, n1673, n1681,
         n1682, n1686, n1707, n1708, n1709, n1710, n1711, n1712, n1722, n1732,
         n1734, n1736, n1737, n1738, n1747, n1748, n1749, n1758, n1759, n1760,
         n1769, n1770, n1771, n1780, n1781, n1782, n1791, n1792, n1793, n1802,
         n1803, n1804, n1813, n1814, n1815, n1824, n1825, n1826, n1835, n1836,
         n1837, n1846, n1847, n1848, n1857, n1868, n1879, n1890, n1901, n1912,
         n1923, n1934, n1945, n1956, n1967, n1978, n1989, n2000, n2011, n2022,
         n2033, n2044, n2055, n2066, n2069, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212;
  wire   [31:0] R14;
  wire   [31:0] sigma0;
  wire   [31:0] R1;
  wire   [31:0] sigma1;
  wire   [31:0] R15;
  wire   [31:0] R6;
  wire   [31:0] logic_result;
  wire   [127:0] buffer;
  wire   [6:0] counter1;
  wire   [6:0] counter2;
  wire   [31:0] R2;
  wire   [31:0] R3;
  wire   [31:0] R4;
  wire   [31:0] R5;
  wire   [31:0] R7;
  wire   [31:0] R8;
  wire   [31:0] R9;
  wire   [31:0] R10;
  wire   [31:0] R11;
  wire   [31:0] R12;
  wire   [31:0] R13;

  AOI2BB1X4 U373 ( .A0N(n1369), .A1N(n62), .B0(reset), .Y(n1336) );
  AOI2BB1X4 U407 ( .A0N(n1405), .A1N(n62), .B0(reset), .Y(n1372) );
  NOR2X4 U441 ( .A(n701), .B(reset), .Y(n1409) );
  NOR2X4 U578 ( .A(n1550), .B(reset), .Y(n1551) );
  NOR2X4 U612 ( .A(n1586), .B(reset), .Y(n1587) );
  AOI2BB1X4 U647 ( .A0N(n1654), .A1N(n1655), .B0(reset), .Y(n1621) );
  NOR2X4 U680 ( .A(n1657), .B(reset), .Y(n1658) );
  AOI2BB1X4 U681 ( .A0N(n1690), .A1N(n1655), .B0(reset), .Y(n1657) );
  NAND3BX4 U682 ( .AN(counter1[6]), .B(n1584), .C(n1548), .Y(n1655) );
  AND3X4 U683 ( .A(n1441), .B(n1691), .C(n1334), .Y(n1584) );
  AND2X2 U689 ( .A(n1695), .B(n1262), .Y(n1152) );
  AND2X2 U690 ( .A(n1696), .B(n1263), .Y(n1153) );
  AND2X2 U698 ( .A(n1156), .B(n1155), .Y(n1334) );
  AND2X2 U709 ( .A(n1704), .B(n1701), .Y(n1654) );
  AND2X2 U710 ( .A(n1583), .B(n1619), .Y(n1548) );
  AND2X2 U714 ( .A(counter1[4]), .B(counter1[5]), .Y(n1704) );
  AND2X2 U716 ( .A(n1703), .B(n1702), .Y(n1546) );
  AND2X2 U719 ( .A(counter1[3]), .B(counter1[2]), .Y(n1701) );
  AND2X2 U722 ( .A(counter1[3]), .B(n1055), .Y(n1703) );
  AND2X2 U1105 ( .A(n2075), .B(n2076), .Y(n1718) );
  AND2X2 U1106 ( .A(n2077), .B(n2075), .Y(n1717) );
  AND2X2 U1108 ( .A(n2078), .B(n2076), .Y(n1720) );
  AND2X2 U1109 ( .A(n2077), .B(n2078), .Y(n1719) );
  AND2X2 U1112 ( .A(n2077), .B(n2079), .Y(n1721) );
  AND2X2 U1114 ( .A(n2080), .B(n2076), .Y(n1723) );
  AND2X2 U1120 ( .A(n2085), .B(n2075), .Y(n1729) );
  AND2X2 U1121 ( .A(n2075), .B(n2086), .Y(n1728) );
  AND2X2 U1122 ( .A(counter2[2]), .B(counter2[1]), .Y(n2075) );
  AND2X2 U1124 ( .A(n2078), .B(n2085), .Y(n1731) );
  AND2X2 U1125 ( .A(n2078), .B(n2086), .Y(n1730) );
  AND2X2 U1126 ( .A(counter2[2]), .B(n1060), .Y(n2078) );
  AND2X2 U1128 ( .A(n2085), .B(n2079), .Y(n1733) );
  AND2X2 U1132 ( .A(n2080), .B(n2085), .Y(n1735) );
  AND2X2 U1142 ( .A(write_enable), .B(n1062), .Y(n2089) );
  CLKINVX4 U1655 ( .A(reset), .Y(n1062) );
  message_schedule_DW01_inc_0 add_564 ( .A(counter2), .SUM({N2175, N2174, 
        N2173, N2172, N2171, N2170, N2169}) );
  message_schedule_DW01_inc_1 add_461 ( .A(counter1), .SUM({N1468, N1467, 
        N1466, N1465, N1464, N1463, N1462}) );
  message_schedule_DW01_add_19 add_0_root_add_0_root_add_35_3 ( .A({N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55}), .B({N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23}), .SUM(logic_result) );
  message_schedule_DW01_add_22 add_1_root_add_0_root_add_35_3 ( .A(sigma1), 
        .B(sigma0), .SUM({N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, 
        N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, 
        N30, N29, N28, N27, N26, N25, N24, N23}) );
  message_schedule_DW01_add_23 add_2_root_add_0_root_add_35_3 ( .A(R15), .B(R6), .SUM({N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, 
        N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, 
        N58, N57, N56, N55}) );
  DFFTRX1 counter1_reg_1_ ( .D(N1463), .RN(n2089), .CK(clk), .Q(counter1[1])
         );
  DFFTRX1 counter1_reg_0_ ( .D(N1462), .RN(n2089), .CK(clk), .Q(counter1[0])
         );
  DFFTRX1 R6_reg_31_ ( .D(R5[31]), .RN(n653), .CK(clk), .Q(R6[31]) );
  DFFTRX1 R15_reg_31_ ( .D(R14[31]), .RN(n652), .CK(clk), .Q(R15[31]) );
  DFFHQXL buffer_reg_14__24_ ( .D(n2159), .CK(clk), .Q(buffer[8]) );
  DFFHQXL buffer_reg_14__25_ ( .D(n2158), .CK(clk), .Q(buffer[9]) );
  DFFHQXL buffer_reg_14__26_ ( .D(n120), .CK(clk), .Q(buffer[10]) );
  DFFHQXL buffer_reg_14__27_ ( .D(n127), .CK(clk), .Q(buffer[11]) );
  DFFHQXL buffer_reg_14__28_ ( .D(n116), .CK(clk), .Q(buffer[12]) );
  DFFHQXL buffer_reg_14__29_ ( .D(n2157), .CK(clk), .Q(buffer[13]) );
  DFFHQXL buffer_reg_14__30_ ( .D(n2156), .CK(clk), .Q(buffer[14]) );
  DFFHQXL buffer_reg_14__31_ ( .D(n2155), .CK(clk), .Q(buffer[15]) );
  DFFHQXL buffer_reg_10__24_ ( .D(n1747), .CK(clk), .Q(buffer[40]) );
  DFFHQXL buffer_reg_10__25_ ( .D(n1738), .CK(clk), .Q(buffer[41]) );
  DFFHQXL buffer_reg_10__26_ ( .D(n1737), .CK(clk), .Q(buffer[42]) );
  DFFHQXL buffer_reg_10__27_ ( .D(n1736), .CK(clk), .Q(buffer[43]) );
  DFFHQXL buffer_reg_10__28_ ( .D(n1734), .CK(clk), .Q(buffer[44]) );
  DFFHQXL buffer_reg_10__29_ ( .D(n1732), .CK(clk), .Q(buffer[45]) );
  DFFHQXL buffer_reg_10__30_ ( .D(n1722), .CK(clk), .Q(buffer[46]) );
  DFFHQXL buffer_reg_10__31_ ( .D(n1712), .CK(clk), .Q(buffer[47]) );
  DFFHQXL buffer_reg_12__24_ ( .D(n2100), .CK(clk), .Q(buffer[24]) );
  DFFHQXL buffer_reg_12__25_ ( .D(n2099), .CK(clk), .Q(buffer[25]) );
  DFFHQXL buffer_reg_12__26_ ( .D(n2098), .CK(clk), .Q(buffer[26]) );
  DFFHQXL buffer_reg_12__27_ ( .D(n2097), .CK(clk), .Q(buffer[27]) );
  DFFHQXL buffer_reg_12__28_ ( .D(n2096), .CK(clk), .Q(buffer[28]) );
  DFFHQXL buffer_reg_12__29_ ( .D(n2095), .CK(clk), .Q(buffer[29]) );
  DFFHQXL buffer_reg_12__30_ ( .D(n2094), .CK(clk), .Q(buffer[30]) );
  DFFHQXL buffer_reg_12__31_ ( .D(n2093), .CK(clk), .Q(buffer[31]) );
  DFFHQX1 buffer_reg_4__24_ ( .D(n963), .CK(clk), .Q(buffer[88]) );
  DFFHQX1 buffer_reg_4__25_ ( .D(n962), .CK(clk), .Q(buffer[89]) );
  DFFHQX1 buffer_reg_4__26_ ( .D(n961), .CK(clk), .Q(buffer[90]) );
  DFFHQX1 buffer_reg_4__27_ ( .D(n960), .CK(clk), .Q(buffer[91]) );
  DFFHQX1 buffer_reg_4__28_ ( .D(n959), .CK(clk), .Q(buffer[92]) );
  DFFHQX1 buffer_reg_4__29_ ( .D(n958), .CK(clk), .Q(buffer[93]) );
  DFFHQX1 buffer_reg_4__30_ ( .D(n957), .CK(clk), .Q(buffer[94]) );
  DFFHQX1 buffer_reg_4__31_ ( .D(n956), .CK(clk), .Q(buffer[95]) );
  DFFHQXL buffer_reg_6__24_ ( .D(n1025), .CK(clk), .Q(buffer[72]) );
  DFFHQXL buffer_reg_6__25_ ( .D(n1024), .CK(clk), .Q(buffer[73]) );
  DFFHQXL buffer_reg_6__26_ ( .D(n1023), .CK(clk), .Q(buffer[74]) );
  DFFHQXL buffer_reg_6__27_ ( .D(n1022), .CK(clk), .Q(buffer[75]) );
  DFFHQXL buffer_reg_6__28_ ( .D(n1021), .CK(clk), .Q(buffer[76]) );
  DFFHQXL buffer_reg_6__29_ ( .D(n1020), .CK(clk), .Q(buffer[77]) );
  DFFHQXL buffer_reg_6__30_ ( .D(n1019), .CK(clk), .Q(buffer[78]) );
  DFFHQXL buffer_reg_6__31_ ( .D(n1018), .CK(clk), .Q(buffer[79]) );
  DFFHQXL buffer_reg_8__24_ ( .D(n1093), .CK(clk), .Q(buffer[56]) );
  DFFHQXL buffer_reg_8__25_ ( .D(n1092), .CK(clk), .Q(buffer[57]) );
  DFFHQXL buffer_reg_8__26_ ( .D(n1091), .CK(clk), .Q(buffer[58]) );
  DFFHQXL buffer_reg_8__27_ ( .D(n1090), .CK(clk), .Q(buffer[59]) );
  DFFHQXL buffer_reg_8__28_ ( .D(n1089), .CK(clk), .Q(buffer[60]) );
  DFFHQXL buffer_reg_8__29_ ( .D(n1088), .CK(clk), .Q(buffer[61]) );
  DFFHQXL buffer_reg_8__30_ ( .D(n1087), .CK(clk), .Q(buffer[62]) );
  DFFHQXL buffer_reg_8__31_ ( .D(n1086), .CK(clk), .Q(buffer[63]) );
  DFFHQXL buffer_reg_15__24_ ( .D(n2183), .CK(clk), .Q(buffer[0]) );
  DFFHQXL buffer_reg_15__25_ ( .D(n2182), .CK(clk), .Q(buffer[1]) );
  DFFHQXL buffer_reg_15__26_ ( .D(n92), .CK(clk), .Q(buffer[2]) );
  DFFHQXL buffer_reg_15__27_ ( .D(n2181), .CK(clk), .Q(buffer[3]) );
  DFFHQXL buffer_reg_15__28_ ( .D(n88), .CK(clk), .Q(buffer[4]) );
  DFFHQXL buffer_reg_15__29_ ( .D(n86), .CK(clk), .Q(buffer[5]) );
  DFFHQXL buffer_reg_15__30_ ( .D(n2180), .CK(clk), .Q(buffer[6]) );
  DFFHQXL buffer_reg_15__31_ ( .D(n102), .CK(clk), .Q(buffer[7]) );
  DFFHQXL buffer_reg_11__24_ ( .D(n1857), .CK(clk), .Q(buffer[32]) );
  DFFHQXL buffer_reg_11__25_ ( .D(n1848), .CK(clk), .Q(buffer[33]) );
  DFFHQXL buffer_reg_11__26_ ( .D(n1847), .CK(clk), .Q(buffer[34]) );
  DFFHQXL buffer_reg_11__27_ ( .D(n1846), .CK(clk), .Q(buffer[35]) );
  DFFHQXL buffer_reg_11__28_ ( .D(n1837), .CK(clk), .Q(buffer[36]) );
  DFFHQXL buffer_reg_11__29_ ( .D(n1836), .CK(clk), .Q(buffer[37]) );
  DFFHQXL buffer_reg_11__30_ ( .D(n1835), .CK(clk), .Q(buffer[38]) );
  DFFHQXL buffer_reg_11__31_ ( .D(n1826), .CK(clk), .Q(buffer[39]) );
  DFFHQXL buffer_reg_13__24_ ( .D(n2131), .CK(clk), .Q(buffer[16]) );
  DFFHQXL buffer_reg_13__25_ ( .D(n2130), .CK(clk), .Q(buffer[17]) );
  DFFHQXL buffer_reg_13__26_ ( .D(n2129), .CK(clk), .Q(buffer[18]) );
  DFFHQXL buffer_reg_13__27_ ( .D(n2128), .CK(clk), .Q(buffer[19]) );
  DFFHQXL buffer_reg_13__28_ ( .D(n2127), .CK(clk), .Q(buffer[20]) );
  DFFHQXL buffer_reg_13__29_ ( .D(n2126), .CK(clk), .Q(buffer[21]) );
  DFFHQXL buffer_reg_13__30_ ( .D(n2125), .CK(clk), .Q(buffer[22]) );
  DFFHQXL buffer_reg_13__31_ ( .D(n2124), .CK(clk), .Q(buffer[23]) );
  DFFHQX1 buffer_reg_5__24_ ( .D(n994), .CK(clk), .Q(buffer[80]) );
  DFFHQX1 buffer_reg_5__25_ ( .D(n993), .CK(clk), .Q(buffer[81]) );
  DFFHQX1 buffer_reg_5__26_ ( .D(n992), .CK(clk), .Q(buffer[82]) );
  DFFHQX1 buffer_reg_5__27_ ( .D(n991), .CK(clk), .Q(buffer[83]) );
  DFFHQX1 buffer_reg_5__29_ ( .D(n989), .CK(clk), .Q(buffer[85]) );
  DFFHQX1 buffer_reg_5__30_ ( .D(n988), .CK(clk), .Q(buffer[86]) );
  DFFHQX1 buffer_reg_5__31_ ( .D(n987), .CK(clk), .Q(buffer[87]) );
  DFFHQXL buffer_reg_7__24_ ( .D(n1065), .CK(clk), .Q(buffer[64]) );
  DFFHQXL buffer_reg_7__25_ ( .D(n1064), .CK(clk), .Q(buffer[65]) );
  DFFHQXL buffer_reg_7__26_ ( .D(n1063), .CK(clk), .Q(buffer[66]) );
  DFFHQXL buffer_reg_7__27_ ( .D(n1053), .CK(clk), .Q(buffer[67]) );
  DFFHQXL buffer_reg_7__28_ ( .D(n1052), .CK(clk), .Q(buffer[68]) );
  DFFHQXL buffer_reg_7__29_ ( .D(n1051), .CK(clk), .Q(buffer[69]) );
  DFFHQXL buffer_reg_7__30_ ( .D(n1050), .CK(clk), .Q(buffer[70]) );
  DFFHQXL buffer_reg_7__31_ ( .D(n1049), .CK(clk), .Q(buffer[71]) );
  DFFHQXL buffer_reg_9__24_ ( .D(n1439), .CK(clk), .Q(buffer[48]) );
  DFFHQXL buffer_reg_9__25_ ( .D(n1438), .CK(clk), .Q(buffer[49]) );
  DFFHQXL buffer_reg_9__26_ ( .D(n1437), .CK(clk), .Q(buffer[50]) );
  DFFHQXL buffer_reg_9__27_ ( .D(n1432), .CK(clk), .Q(buffer[51]) );
  DFFHQXL buffer_reg_9__28_ ( .D(n1228), .CK(clk), .Q(buffer[52]) );
  DFFHQXL buffer_reg_9__29_ ( .D(n1192), .CK(clk), .Q(buffer[53]) );
  DFFHQXL buffer_reg_9__30_ ( .D(n1159), .CK(clk), .Q(buffer[54]) );
  DFFHQXL buffer_reg_9__31_ ( .D(n1150), .CK(clk), .Q(buffer[55]) );
  DFFHQXL buffer_reg_14__0_ ( .D(n2199), .CK(clk), .Q(N890) );
  DFFHQXL buffer_reg_14__1_ ( .D(n2154), .CK(clk), .Q(N891) );
  DFFHQXL buffer_reg_14__2_ ( .D(n2153), .CK(clk), .Q(N892) );
  DFFHQXL buffer_reg_14__3_ ( .D(n2152), .CK(clk), .Q(N893) );
  DFFHQXL buffer_reg_14__4_ ( .D(n2151), .CK(clk), .Q(N894) );
  DFFHQXL buffer_reg_14__5_ ( .D(n2150), .CK(clk), .Q(N895) );
  DFFHQXL buffer_reg_14__6_ ( .D(n2149), .CK(clk), .Q(N896) );
  DFFHQXL buffer_reg_14__7_ ( .D(n2148), .CK(clk), .Q(N897) );
  DFFHQXL buffer_reg_14__8_ ( .D(n2174), .CK(clk), .Q(N898) );
  DFFHQXL buffer_reg_14__9_ ( .D(n2173), .CK(clk), .Q(N899) );
  DFFHQXL buffer_reg_14__10_ ( .D(n2172), .CK(clk), .Q(N900) );
  DFFHQXL buffer_reg_14__11_ ( .D(n2171), .CK(clk), .Q(N901) );
  DFFHQXL buffer_reg_14__12_ ( .D(n2170), .CK(clk), .Q(N902) );
  DFFHQXL buffer_reg_14__13_ ( .D(n2169), .CK(clk), .Q(N903) );
  DFFHQXL buffer_reg_14__14_ ( .D(n131), .CK(clk), .Q(N904) );
  DFFHQXL buffer_reg_14__15_ ( .D(n2168), .CK(clk), .Q(N905) );
  DFFHQXL buffer_reg_14__16_ ( .D(n2167), .CK(clk), .Q(N906) );
  DFFHQXL buffer_reg_14__17_ ( .D(n2166), .CK(clk), .Q(N907) );
  DFFHQXL buffer_reg_14__18_ ( .D(n2165), .CK(clk), .Q(N908) );
  DFFHQXL buffer_reg_14__19_ ( .D(n2164), .CK(clk), .Q(N909) );
  DFFHQXL buffer_reg_14__20_ ( .D(n2163), .CK(clk), .Q(N910) );
  DFFHQXL buffer_reg_14__21_ ( .D(n2162), .CK(clk), .Q(N911) );
  DFFHQXL buffer_reg_14__22_ ( .D(n2161), .CK(clk), .Q(N912) );
  DFFHQXL buffer_reg_14__23_ ( .D(n2160), .CK(clk), .Q(N913) );
  DFFHQXL buffer_reg_10__0_ ( .D(n2203), .CK(clk), .Q(N762) );
  DFFHQXL buffer_reg_10__1_ ( .D(n1711), .CK(clk), .Q(N763) );
  DFFHQXL buffer_reg_10__2_ ( .D(n1710), .CK(clk), .Q(N764) );
  DFFHQXL buffer_reg_10__3_ ( .D(n1709), .CK(clk), .Q(N765) );
  DFFHQXL buffer_reg_10__4_ ( .D(n1708), .CK(clk), .Q(N766) );
  DFFHQXL buffer_reg_10__5_ ( .D(n1707), .CK(clk), .Q(N767) );
  DFFHQXL buffer_reg_10__6_ ( .D(n1686), .CK(clk), .Q(N768) );
  DFFHQXL buffer_reg_10__7_ ( .D(n1682), .CK(clk), .Q(N769) );
  DFFHQXL buffer_reg_10__8_ ( .D(n1803), .CK(clk), .Q(N770) );
  DFFHQXL buffer_reg_10__9_ ( .D(n1802), .CK(clk), .Q(N771) );
  DFFHQXL buffer_reg_10__10_ ( .D(n1793), .CK(clk), .Q(N772) );
  DFFHQXL buffer_reg_10__11_ ( .D(n1792), .CK(clk), .Q(N773) );
  DFFHQXL buffer_reg_10__12_ ( .D(n1791), .CK(clk), .Q(N774) );
  DFFHQXL buffer_reg_10__13_ ( .D(n1782), .CK(clk), .Q(N775) );
  DFFHQXL buffer_reg_10__14_ ( .D(n1781), .CK(clk), .Q(N776) );
  DFFHQXL buffer_reg_10__15_ ( .D(n1780), .CK(clk), .Q(N777) );
  DFFHQXL buffer_reg_10__16_ ( .D(n1771), .CK(clk), .Q(N778) );
  DFFHQXL buffer_reg_10__17_ ( .D(n1770), .CK(clk), .Q(N779) );
  DFFHQXL buffer_reg_10__18_ ( .D(n1769), .CK(clk), .Q(N780) );
  DFFHQXL buffer_reg_10__19_ ( .D(n1760), .CK(clk), .Q(N781) );
  DFFHQXL buffer_reg_10__20_ ( .D(n1759), .CK(clk), .Q(N782) );
  DFFHQXL buffer_reg_10__21_ ( .D(n1758), .CK(clk), .Q(N783) );
  DFFHQXL buffer_reg_10__22_ ( .D(n1749), .CK(clk), .Q(N784) );
  DFFHQXL buffer_reg_10__23_ ( .D(n1748), .CK(clk), .Q(N785) );
  DFFHQXL buffer_reg_12__0_ ( .D(n2201), .CK(clk), .Q(N826) );
  DFFHQXL buffer_reg_12__1_ ( .D(n2092), .CK(clk), .Q(N827) );
  DFFHQXL buffer_reg_12__2_ ( .D(n2091), .CK(clk), .Q(N828) );
  DFFHQXL buffer_reg_12__3_ ( .D(n2090), .CK(clk), .Q(N829) );
  DFFHQXL buffer_reg_12__4_ ( .D(n2069), .CK(clk), .Q(N830) );
  DFFHQXL buffer_reg_12__5_ ( .D(n2066), .CK(clk), .Q(N831) );
  DFFHQXL buffer_reg_12__6_ ( .D(n2055), .CK(clk), .Q(N832) );
  DFFHQXL buffer_reg_12__7_ ( .D(n2044), .CK(clk), .Q(N833) );
  DFFHQXL buffer_reg_12__8_ ( .D(n2116), .CK(clk), .Q(N834) );
  DFFHQXL buffer_reg_12__9_ ( .D(n2115), .CK(clk), .Q(N835) );
  DFFHQXL buffer_reg_12__10_ ( .D(n2114), .CK(clk), .Q(N836) );
  DFFHQXL buffer_reg_12__11_ ( .D(n2113), .CK(clk), .Q(N837) );
  DFFHQXL buffer_reg_12__12_ ( .D(n2112), .CK(clk), .Q(N838) );
  DFFHQXL buffer_reg_12__13_ ( .D(n2111), .CK(clk), .Q(N839) );
  DFFHQXL buffer_reg_12__14_ ( .D(n2110), .CK(clk), .Q(N840) );
  DFFHQXL buffer_reg_12__15_ ( .D(n2109), .CK(clk), .Q(N841) );
  DFFHQXL buffer_reg_12__16_ ( .D(n2108), .CK(clk), .Q(N842) );
  DFFHQXL buffer_reg_12__17_ ( .D(n2107), .CK(clk), .Q(N843) );
  DFFHQXL buffer_reg_12__18_ ( .D(n2106), .CK(clk), .Q(N844) );
  DFFHQXL buffer_reg_12__19_ ( .D(n2105), .CK(clk), .Q(N845) );
  DFFHQXL buffer_reg_12__20_ ( .D(n2104), .CK(clk), .Q(N846) );
  DFFHQXL buffer_reg_12__21_ ( .D(n2103), .CK(clk), .Q(N847) );
  DFFHQXL buffer_reg_12__22_ ( .D(n2102), .CK(clk), .Q(N848) );
  DFFHQXL buffer_reg_12__23_ ( .D(n2101), .CK(clk), .Q(N849) );
  DFFHQX1 buffer_reg_4__0_ ( .D(n2209), .CK(clk), .Q(N570) );
  DFFHQX1 buffer_reg_4__1_ ( .D(n955), .CK(clk), .Q(N571) );
  DFFHQX1 buffer_reg_4__2_ ( .D(n954), .CK(clk), .Q(N572) );
  DFFHQX1 buffer_reg_4__3_ ( .D(n953), .CK(clk), .Q(N573) );
  DFFHQX1 buffer_reg_4__4_ ( .D(n952), .CK(clk), .Q(N574) );
  DFFHQX1 buffer_reg_4__5_ ( .D(n951), .CK(clk), .Q(N575) );
  DFFHQX1 buffer_reg_4__6_ ( .D(n950), .CK(clk), .Q(N576) );
  DFFHQX1 buffer_reg_4__7_ ( .D(n949), .CK(clk), .Q(N577) );
  DFFHQX1 buffer_reg_4__8_ ( .D(n979), .CK(clk), .Q(N578) );
  DFFHQX1 buffer_reg_4__9_ ( .D(n978), .CK(clk), .Q(N579) );
  DFFHQX1 buffer_reg_4__10_ ( .D(n977), .CK(clk), .Q(N580) );
  DFFHQX1 buffer_reg_4__11_ ( .D(n976), .CK(clk), .Q(N581) );
  DFFHQX1 buffer_reg_4__12_ ( .D(n975), .CK(clk), .Q(N582) );
  DFFHQX1 buffer_reg_4__13_ ( .D(n974), .CK(clk), .Q(N583) );
  DFFHQX1 buffer_reg_4__14_ ( .D(n973), .CK(clk), .Q(N584) );
  DFFHQX1 buffer_reg_4__15_ ( .D(n972), .CK(clk), .Q(N585) );
  DFFHQX1 buffer_reg_4__16_ ( .D(n971), .CK(clk), .Q(N586) );
  DFFHQX1 buffer_reg_4__17_ ( .D(n970), .CK(clk), .Q(N587) );
  DFFHQX1 buffer_reg_4__18_ ( .D(n969), .CK(clk), .Q(N588) );
  DFFHQX1 buffer_reg_4__19_ ( .D(n968), .CK(clk), .Q(N589) );
  DFFHQX1 buffer_reg_4__20_ ( .D(n967), .CK(clk), .Q(N590) );
  DFFHQX1 buffer_reg_4__21_ ( .D(n966), .CK(clk), .Q(N591) );
  DFFHQX1 buffer_reg_4__22_ ( .D(n965), .CK(clk), .Q(N592) );
  DFFHQX1 buffer_reg_4__23_ ( .D(n964), .CK(clk), .Q(N593) );
  DFFHQXL buffer_reg_6__0_ ( .D(n2207), .CK(clk), .Q(N634) );
  DFFHQXL buffer_reg_6__1_ ( .D(n1017), .CK(clk), .Q(N635) );
  DFFHQXL buffer_reg_6__2_ ( .D(n1016), .CK(clk), .Q(N636) );
  DFFHQXL buffer_reg_6__3_ ( .D(n1015), .CK(clk), .Q(N637) );
  DFFHQXL buffer_reg_6__4_ ( .D(n1014), .CK(clk), .Q(N638) );
  DFFHQXL buffer_reg_6__5_ ( .D(n1013), .CK(clk), .Q(N639) );
  DFFHQXL buffer_reg_6__6_ ( .D(n1012), .CK(clk), .Q(N640) );
  DFFHQXL buffer_reg_6__7_ ( .D(n1011), .CK(clk), .Q(N641) );
  DFFHQXL buffer_reg_6__8_ ( .D(n1041), .CK(clk), .Q(N642) );
  DFFHQXL buffer_reg_6__9_ ( .D(n1040), .CK(clk), .Q(N643) );
  DFFHQXL buffer_reg_6__10_ ( .D(n1039), .CK(clk), .Q(N644) );
  DFFHQXL buffer_reg_6__11_ ( .D(n1038), .CK(clk), .Q(N645) );
  DFFHQXL buffer_reg_6__12_ ( .D(n1037), .CK(clk), .Q(N646) );
  DFFHQXL buffer_reg_6__13_ ( .D(n1036), .CK(clk), .Q(N647) );
  DFFHQXL buffer_reg_6__14_ ( .D(n1035), .CK(clk), .Q(N648) );
  DFFHQXL buffer_reg_6__15_ ( .D(n1034), .CK(clk), .Q(N649) );
  DFFHQXL buffer_reg_6__16_ ( .D(n1033), .CK(clk), .Q(N650) );
  DFFHQXL buffer_reg_6__17_ ( .D(n1032), .CK(clk), .Q(N651) );
  DFFHQXL buffer_reg_6__18_ ( .D(n1031), .CK(clk), .Q(N652) );
  DFFHQXL buffer_reg_6__19_ ( .D(n1030), .CK(clk), .Q(N653) );
  DFFHQXL buffer_reg_6__20_ ( .D(n1029), .CK(clk), .Q(N654) );
  DFFHQXL buffer_reg_6__21_ ( .D(n1028), .CK(clk), .Q(N655) );
  DFFHQXL buffer_reg_6__22_ ( .D(n1027), .CK(clk), .Q(N656) );
  DFFHQXL buffer_reg_6__23_ ( .D(n1026), .CK(clk), .Q(N657) );
  DFFHQXL buffer_reg_8__0_ ( .D(n2205), .CK(clk), .Q(N698) );
  DFFHQXL buffer_reg_8__1_ ( .D(n106), .CK(clk), .Q(N699) );
  DFFHQXL buffer_reg_8__2_ ( .D(n98), .CK(clk), .Q(N700) );
  DFFHQXL buffer_reg_8__3_ ( .D(n78), .CK(clk), .Q(N701) );
  DFFHQXL buffer_reg_8__4_ ( .D(n1085), .CK(clk), .Q(N702) );
  DFFHQXL buffer_reg_8__5_ ( .D(n1084), .CK(clk), .Q(N703) );
  DFFHQXL buffer_reg_8__6_ ( .D(n1083), .CK(clk), .Q(N704) );
  DFFHQXL buffer_reg_8__7_ ( .D(n1082), .CK(clk), .Q(N705) );
  DFFHQXL buffer_reg_8__8_ ( .D(n83), .CK(clk), .Q(N706) );
  DFFHQXL buffer_reg_8__9_ ( .D(n1108), .CK(clk), .Q(N707) );
  DFFHQXL buffer_reg_8__10_ ( .D(n1107), .CK(clk), .Q(N708) );
  DFFHQXL buffer_reg_8__11_ ( .D(n1106), .CK(clk), .Q(N709) );
  DFFHQXL buffer_reg_8__12_ ( .D(n1105), .CK(clk), .Q(N710) );
  DFFHQXL buffer_reg_8__13_ ( .D(n1104), .CK(clk), .Q(N711) );
  DFFHQXL buffer_reg_8__14_ ( .D(n1103), .CK(clk), .Q(N712) );
  DFFHQXL buffer_reg_8__15_ ( .D(n1102), .CK(clk), .Q(N713) );
  DFFHQXL buffer_reg_8__16_ ( .D(n1101), .CK(clk), .Q(N714) );
  DFFHQXL buffer_reg_8__17_ ( .D(n1100), .CK(clk), .Q(N715) );
  DFFHQXL buffer_reg_8__18_ ( .D(n1099), .CK(clk), .Q(N716) );
  DFFHQXL buffer_reg_8__19_ ( .D(n1098), .CK(clk), .Q(N717) );
  DFFHQXL buffer_reg_8__20_ ( .D(n1097), .CK(clk), .Q(N718) );
  DFFHQXL buffer_reg_8__21_ ( .D(n1096), .CK(clk), .Q(N719) );
  DFFHQXL buffer_reg_8__22_ ( .D(n1095), .CK(clk), .Q(N720) );
  DFFHQXL buffer_reg_8__23_ ( .D(n1094), .CK(clk), .Q(N721) );
  DFFHQXL buffer_reg_15__0_ ( .D(n2198), .CK(clk), .Q(N922) );
  DFFHQXL buffer_reg_15__1_ ( .D(n2179), .CK(clk), .Q(N923) );
  DFFHQXL buffer_reg_15__2_ ( .D(n2178), .CK(clk), .Q(N924) );
  DFFHQXL buffer_reg_15__3_ ( .D(n118), .CK(clk), .Q(N925) );
  DFFHQXL buffer_reg_15__4_ ( .D(n2177), .CK(clk), .Q(N926) );
  DFFHQXL buffer_reg_15__5_ ( .D(n2176), .CK(clk), .Q(N927) );
  DFFHQXL buffer_reg_15__6_ ( .D(n2175), .CK(clk), .Q(N928) );
  DFFHQXL buffer_reg_15__7_ ( .D(n123), .CK(clk), .Q(N929) );
  DFFHQXL buffer_reg_15__8_ ( .D(n90), .CK(clk), .Q(N930) );
  DFFHQXL buffer_reg_15__9_ ( .D(n2195), .CK(clk), .Q(N931) );
  DFFHQXL buffer_reg_15__10_ ( .D(n2194), .CK(clk), .Q(N932) );
  DFFHQXL buffer_reg_15__11_ ( .D(n2193), .CK(clk), .Q(N933) );
  DFFHQXL buffer_reg_15__12_ ( .D(n2192), .CK(clk), .Q(N934) );
  DFFHQXL buffer_reg_15__13_ ( .D(n2191), .CK(clk), .Q(N935) );
  DFFHQXL buffer_reg_15__14_ ( .D(n2190), .CK(clk), .Q(N936) );
  DFFHQXL buffer_reg_15__15_ ( .D(n2189), .CK(clk), .Q(N937) );
  DFFHQXL buffer_reg_15__16_ ( .D(n81), .CK(clk), .Q(N938) );
  DFFHQXL buffer_reg_15__17_ ( .D(n96), .CK(clk), .Q(N939) );
  DFFHQXL buffer_reg_15__18_ ( .D(n2188), .CK(clk), .Q(N940) );
  DFFHQXL buffer_reg_15__19_ ( .D(n2187), .CK(clk), .Q(N941) );
  DFFHQXL buffer_reg_15__20_ ( .D(n94), .CK(clk), .Q(N942) );
  DFFHQXL buffer_reg_15__21_ ( .D(n2186), .CK(clk), .Q(N943) );
  DFFHQXL buffer_reg_15__22_ ( .D(n2185), .CK(clk), .Q(N944) );
  DFFHQXL buffer_reg_15__23_ ( .D(n2184), .CK(clk), .Q(N945) );
  DFFHQXL buffer_reg_11__0_ ( .D(n2202), .CK(clk), .Q(N794) );
  DFFHQXL buffer_reg_11__1_ ( .D(n1825), .CK(clk), .Q(N795) );
  DFFHQXL buffer_reg_11__2_ ( .D(n1824), .CK(clk), .Q(N796) );
  DFFHQXL buffer_reg_11__3_ ( .D(n1815), .CK(clk), .Q(N797) );
  DFFHQXL buffer_reg_11__4_ ( .D(n65), .CK(clk), .Q(N798) );
  DFFHQXL buffer_reg_11__5_ ( .D(n1814), .CK(clk), .Q(N799) );
  DFFHQXL buffer_reg_11__6_ ( .D(n1813), .CK(clk), .Q(N800) );
  DFFHQXL buffer_reg_11__7_ ( .D(n1804), .CK(clk), .Q(N801) );
  DFFHQXL buffer_reg_11__8_ ( .D(n2033), .CK(clk), .Q(N802) );
  DFFHQXL buffer_reg_11__9_ ( .D(n2022), .CK(clk), .Q(N803) );
  DFFHQXL buffer_reg_11__10_ ( .D(n2011), .CK(clk), .Q(N804) );
  DFFHQXL buffer_reg_11__11_ ( .D(n2000), .CK(clk), .Q(N805) );
  DFFHQXL buffer_reg_11__12_ ( .D(n1989), .CK(clk), .Q(N806) );
  DFFHQXL buffer_reg_11__13_ ( .D(n1978), .CK(clk), .Q(N807) );
  DFFHQXL buffer_reg_11__14_ ( .D(n1967), .CK(clk), .Q(N808) );
  DFFHQXL buffer_reg_11__15_ ( .D(n1956), .CK(clk), .Q(N809) );
  DFFHQXL buffer_reg_11__16_ ( .D(n1945), .CK(clk), .Q(N810) );
  DFFHQXL buffer_reg_11__17_ ( .D(n1934), .CK(clk), .Q(N811) );
  DFFHQXL buffer_reg_11__18_ ( .D(n1923), .CK(clk), .Q(N812) );
  DFFHQXL buffer_reg_11__20_ ( .D(n1901), .CK(clk), .Q(N814) );
  DFFHQXL buffer_reg_11__21_ ( .D(n1890), .CK(clk), .Q(N815) );
  DFFHQXL buffer_reg_11__22_ ( .D(n1879), .CK(clk), .Q(N816) );
  DFFHQXL buffer_reg_11__23_ ( .D(n1868), .CK(clk), .Q(N817) );
  DFFHQXL buffer_reg_13__0_ ( .D(n2200), .CK(clk), .Q(N858) );
  DFFHQXL buffer_reg_13__1_ ( .D(n2123), .CK(clk), .Q(N859) );
  DFFHQXL buffer_reg_13__2_ ( .D(n2122), .CK(clk), .Q(N860) );
  DFFHQXL buffer_reg_13__3_ ( .D(n2121), .CK(clk), .Q(N861) );
  DFFHQXL buffer_reg_13__4_ ( .D(n2120), .CK(clk), .Q(N862) );
  DFFHQXL buffer_reg_13__5_ ( .D(n2119), .CK(clk), .Q(N863) );
  DFFHQXL buffer_reg_13__6_ ( .D(n2118), .CK(clk), .Q(N864) );
  DFFHQXL buffer_reg_13__7_ ( .D(n2117), .CK(clk), .Q(N865) );
  DFFHQXL buffer_reg_13__8_ ( .D(n2147), .CK(clk), .Q(N866) );
  DFFHQXL buffer_reg_13__9_ ( .D(n2146), .CK(clk), .Q(N867) );
  DFFHQXL buffer_reg_13__10_ ( .D(n2145), .CK(clk), .Q(N868) );
  DFFHQXL buffer_reg_13__11_ ( .D(n2144), .CK(clk), .Q(N869) );
  DFFHQXL buffer_reg_13__12_ ( .D(n2143), .CK(clk), .Q(N870) );
  DFFHQXL buffer_reg_13__13_ ( .D(n2142), .CK(clk), .Q(N871) );
  DFFHQXL buffer_reg_13__14_ ( .D(n2141), .CK(clk), .Q(N872) );
  DFFHQXL buffer_reg_13__15_ ( .D(n2140), .CK(clk), .Q(N873) );
  DFFHQXL buffer_reg_13__16_ ( .D(n2139), .CK(clk), .Q(N874) );
  DFFHQXL buffer_reg_13__17_ ( .D(n2138), .CK(clk), .Q(N875) );
  DFFHQXL buffer_reg_13__18_ ( .D(n2137), .CK(clk), .Q(N876) );
  DFFHQXL buffer_reg_13__19_ ( .D(n2136), .CK(clk), .Q(N877) );
  DFFHQXL buffer_reg_13__20_ ( .D(n2135), .CK(clk), .Q(N878) );
  DFFHQXL buffer_reg_13__21_ ( .D(n2134), .CK(clk), .Q(N879) );
  DFFHQXL buffer_reg_13__22_ ( .D(n2133), .CK(clk), .Q(N880) );
  DFFHQXL buffer_reg_13__23_ ( .D(n2132), .CK(clk), .Q(N881) );
  DFFHQXL buffer_reg_5__0_ ( .D(n2208), .CK(clk), .Q(N602) );
  DFFHQXL buffer_reg_5__1_ ( .D(n986), .CK(clk), .Q(N603) );
  DFFHQXL buffer_reg_5__2_ ( .D(n985), .CK(clk), .Q(N604) );
  DFFHQXL buffer_reg_5__3_ ( .D(n984), .CK(clk), .Q(N605) );
  DFFHQXL buffer_reg_5__4_ ( .D(n983), .CK(clk), .Q(N606) );
  DFFHQXL buffer_reg_5__5_ ( .D(n982), .CK(clk), .Q(N607) );
  DFFHQXL buffer_reg_5__6_ ( .D(n981), .CK(clk), .Q(N608) );
  DFFHQXL buffer_reg_5__7_ ( .D(n980), .CK(clk), .Q(N609) );
  DFFHQXL buffer_reg_5__8_ ( .D(n1010), .CK(clk), .Q(N610) );
  DFFHQXL buffer_reg_5__9_ ( .D(n1009), .CK(clk), .Q(N611) );
  DFFHQXL buffer_reg_5__10_ ( .D(n1008), .CK(clk), .Q(N612) );
  DFFHQXL buffer_reg_5__11_ ( .D(n1007), .CK(clk), .Q(N613) );
  DFFHQXL buffer_reg_5__12_ ( .D(n1006), .CK(clk), .Q(N614) );
  DFFHQXL buffer_reg_5__13_ ( .D(n1005), .CK(clk), .Q(N615) );
  DFFHQXL buffer_reg_5__14_ ( .D(n1004), .CK(clk), .Q(N616) );
  DFFHQXL buffer_reg_5__15_ ( .D(n1003), .CK(clk), .Q(N617) );
  DFFHQXL buffer_reg_5__16_ ( .D(n1002), .CK(clk), .Q(N618) );
  DFFHQXL buffer_reg_5__17_ ( .D(n1001), .CK(clk), .Q(N619) );
  DFFHQXL buffer_reg_5__18_ ( .D(n1000), .CK(clk), .Q(N620) );
  DFFHQXL buffer_reg_5__19_ ( .D(n999), .CK(clk), .Q(N621) );
  DFFHQXL buffer_reg_5__20_ ( .D(n998), .CK(clk), .Q(N622) );
  DFFHQXL buffer_reg_5__21_ ( .D(n997), .CK(clk), .Q(N623) );
  DFFHQXL buffer_reg_5__22_ ( .D(n996), .CK(clk), .Q(N624) );
  DFFHQXL buffer_reg_5__23_ ( .D(n995), .CK(clk), .Q(N625) );
  DFFHQXL buffer_reg_7__0_ ( .D(n2206), .CK(clk), .Q(N666) );
  DFFHQXL buffer_reg_7__1_ ( .D(n1048), .CK(clk), .Q(N667) );
  DFFHQXL buffer_reg_7__2_ ( .D(n1047), .CK(clk), .Q(N668) );
  DFFHQXL buffer_reg_7__3_ ( .D(n1046), .CK(clk), .Q(N669) );
  DFFHQXL buffer_reg_7__4_ ( .D(n1045), .CK(clk), .Q(N670) );
  DFFHQXL buffer_reg_7__5_ ( .D(n1044), .CK(clk), .Q(N671) );
  DFFHQXL buffer_reg_7__6_ ( .D(n1043), .CK(clk), .Q(N672) );
  DFFHQXL buffer_reg_7__7_ ( .D(n1042), .CK(clk), .Q(N673) );
  DFFHQXL buffer_reg_7__8_ ( .D(n1081), .CK(clk), .Q(N674) );
  DFFHQXL buffer_reg_7__9_ ( .D(n1080), .CK(clk), .Q(N675) );
  DFFHQXL buffer_reg_7__10_ ( .D(n1079), .CK(clk), .Q(N676) );
  DFFHQXL buffer_reg_7__11_ ( .D(n1078), .CK(clk), .Q(N677) );
  DFFHQXL buffer_reg_7__12_ ( .D(n1077), .CK(clk), .Q(N678) );
  DFFHQXL buffer_reg_7__13_ ( .D(n1076), .CK(clk), .Q(N679) );
  DFFHQXL buffer_reg_7__14_ ( .D(n1075), .CK(clk), .Q(N680) );
  DFFHQXL buffer_reg_7__15_ ( .D(n1074), .CK(clk), .Q(N681) );
  DFFHQXL buffer_reg_7__16_ ( .D(n1073), .CK(clk), .Q(N682) );
  DFFHQXL buffer_reg_7__17_ ( .D(n1072), .CK(clk), .Q(N683) );
  DFFHQXL buffer_reg_7__18_ ( .D(n1071), .CK(clk), .Q(N684) );
  DFFHQXL buffer_reg_7__19_ ( .D(n1070), .CK(clk), .Q(N685) );
  DFFHQXL buffer_reg_7__20_ ( .D(n1069), .CK(clk), .Q(N686) );
  DFFHQXL buffer_reg_7__21_ ( .D(n1068), .CK(clk), .Q(N687) );
  DFFHQXL buffer_reg_7__22_ ( .D(n1067), .CK(clk), .Q(N688) );
  DFFHQXL buffer_reg_7__23_ ( .D(n1066), .CK(clk), .Q(N689) );
  DFFHQXL buffer_reg_9__0_ ( .D(n2204), .CK(clk), .Q(N730) );
  DFFHQXL buffer_reg_9__1_ ( .D(n108), .CK(clk), .Q(N731) );
  DFFHQXL buffer_reg_9__2_ ( .D(n100), .CK(clk), .Q(N732) );
  DFFHQXL buffer_reg_9__3_ ( .D(n1113), .CK(clk), .Q(N733) );
  DFFHQXL buffer_reg_9__4_ ( .D(n1112), .CK(clk), .Q(N734) );
  DFFHQXL buffer_reg_9__5_ ( .D(n1111), .CK(clk), .Q(N735) );
  DFFHQXL buffer_reg_9__6_ ( .D(n1110), .CK(clk), .Q(N736) );
  DFFHQXL buffer_reg_9__7_ ( .D(n1109), .CK(clk), .Q(N737) );
  DFFHQXL buffer_reg_9__8_ ( .D(n1681), .CK(clk), .Q(N738) );
  DFFHQXL buffer_reg_9__9_ ( .D(n1673), .CK(clk), .Q(N739) );
  DFFHQXL buffer_reg_9__10_ ( .D(n1672), .CK(clk), .Q(N740) );
  DFFHQXL buffer_reg_9__11_ ( .D(n1669), .CK(clk), .Q(N741) );
  DFFHQXL buffer_reg_9__12_ ( .D(n1663), .CK(clk), .Q(N742) );
  DFFHQXL buffer_reg_9__13_ ( .D(n1661), .CK(clk), .Q(N743) );
  DFFHQXL buffer_reg_9__14_ ( .D(n1660), .CK(clk), .Q(N744) );
  DFFHQXL buffer_reg_9__15_ ( .D(n1656), .CK(clk), .Q(N745) );
  DFFHQXL buffer_reg_9__16_ ( .D(n1639), .CK(clk), .Q(N746) );
  DFFHQXL buffer_reg_9__17_ ( .D(n1627), .CK(clk), .Q(N747) );
  DFFHQXL buffer_reg_9__18_ ( .D(n1626), .CK(clk), .Q(N748) );
  DFFHQXL buffer_reg_9__19_ ( .D(n1625), .CK(clk), .Q(N749) );
  DFFHQXL buffer_reg_9__20_ ( .D(n1541), .CK(clk), .Q(N750) );
  DFFHQXL buffer_reg_9__21_ ( .D(n1478), .CK(clk), .Q(N751) );
  DFFHQXL buffer_reg_9__22_ ( .D(n1474), .CK(clk), .Q(N752) );
  DFFHQXL buffer_reg_9__23_ ( .D(n1473), .CK(clk), .Q(N753) );
  DFFHQX1 Wt_reg_30_ ( .D(N2161), .CK(clk), .Q(Wt[30]) );
  DFFTRX1 counter2_reg_6_ ( .D(N2175), .RN(n1705), .CK(clk), .Q(counter2[6]), 
        .QN(n1056) );
  DFFTRX1 counter2_reg_4_ ( .D(N2173), .RN(n1705), .CK(clk), .Q(counter2[4]), 
        .QN(n1058) );
  DFFTRX1 counter2_reg_5_ ( .D(N2174), .RN(n1705), .CK(clk), .Q(counter2[5]), 
        .QN(n1057) );
  DFFTRX1 R15_reg_30_ ( .D(R14[30]), .RN(n651), .CK(clk), .Q(R15[30]) );
  DFFTRX1 R15_reg_29_ ( .D(R14[29]), .RN(n650), .CK(clk), .Q(R15[29]) );
  DFFTRX1 R15_reg_28_ ( .D(R14[28]), .RN(n649), .CK(clk), .Q(R15[28]) );
  DFFTRX1 R6_reg_30_ ( .D(R5[30]), .RN(n652), .CK(clk), .Q(R6[30]) );
  DFFTRX1 R6_reg_29_ ( .D(R5[29]), .RN(n651), .CK(clk), .Q(R6[29]) );
  DFFTRX1 R6_reg_28_ ( .D(R5[28]), .RN(n649), .CK(clk), .Q(R6[28]) );
  DFFTRX1 counter2_reg_3_ ( .D(N2172), .RN(n1705), .CK(clk), .Q(counter2[3]), 
        .QN(n1059) );
  DFFTRX1 counter2_reg_1_ ( .D(N2170), .RN(n1705), .CK(clk), .Q(counter2[1]), 
        .QN(n1060) );
  DFFTRX1 counter2_reg_0_ ( .D(N2169), .RN(n1705), .CK(clk), .Q(counter2[0]), 
        .QN(n1061) );
  DFFTRX1 counter2_reg_2_ ( .D(N2171), .RN(n1705), .CK(clk), .Q(counter2[2])
         );
  DFFTRX1 R15_reg_27_ ( .D(R14[27]), .RN(n647), .CK(clk), .Q(R15[27]) );
  DFFTRX1 R15_reg_26_ ( .D(R14[26]), .RN(n646), .CK(clk), .Q(R15[26]) );
  DFFTRX1 R15_reg_25_ ( .D(R14[25]), .RN(n645), .CK(clk), .Q(R15[25]) );
  DFFTRX1 R15_reg_24_ ( .D(R14[24]), .RN(n644), .CK(clk), .Q(R15[24]) );
  DFFTRX1 R6_reg_27_ ( .D(R5[27]), .RN(n648), .CK(clk), .Q(R6[27]) );
  DFFTRX1 R6_reg_26_ ( .D(R5[26]), .RN(n647), .CK(clk), .Q(R6[26]) );
  DFFTRX1 R6_reg_25_ ( .D(R5[25]), .RN(n646), .CK(clk), .Q(R6[25]) );
  DFFTRX1 R6_reg_24_ ( .D(R5[24]), .RN(n644), .CK(clk), .Q(R6[24]) );
  DFFTRX1 counter1_reg_6_ ( .D(N1468), .RN(n2089), .CK(clk), .Q(counter1[6])
         );
  DFFTRX1 counter1_reg_2_ ( .D(N1464), .RN(n2089), .CK(clk), .Q(counter1[2]), 
        .QN(n1055) );
  DFFTRX1 R15_reg_23_ ( .D(R14[23]), .RN(n642), .CK(clk), .Q(R15[23]) );
  DFFTRX1 R15_reg_22_ ( .D(R14[22]), .RN(n641), .CK(clk), .Q(R15[22]) );
  DFFTRX1 R15_reg_21_ ( .D(R14[21]), .RN(n640), .CK(clk), .Q(R15[21]) );
  DFFTRX1 R15_reg_20_ ( .D(R14[20]), .RN(n639), .CK(clk), .Q(R15[20]) );
  DFFTRX1 R15_reg_19_ ( .D(R14[19]), .RN(n637), .CK(clk), .Q(R15[19]) );
  DFFTRX1 R15_reg_18_ ( .D(R14[18]), .RN(n636), .CK(clk), .Q(R15[18]) );
  DFFTRX1 R6_reg_23_ ( .D(R5[23]), .RN(n643), .CK(clk), .Q(R6[23]) );
  DFFTRX1 R6_reg_22_ ( .D(R5[22]), .RN(n642), .CK(clk), .Q(R6[22]) );
  DFFTRX1 R6_reg_21_ ( .D(R5[21]), .RN(n641), .CK(clk), .Q(R6[21]) );
  DFFTRX1 R6_reg_20_ ( .D(R5[20]), .RN(n639), .CK(clk), .Q(R6[20]) );
  DFFTRX1 R6_reg_19_ ( .D(R5[19]), .RN(n638), .CK(clk), .Q(R6[19]) );
  DFFTRX1 R6_reg_18_ ( .D(R5[18]), .RN(n637), .CK(clk), .Q(R6[18]) );
  DFFTRX1 R6_reg_16_ ( .D(R5[16]), .RN(n634), .CK(clk), .Q(R6[16]) );
  DFFTRX1 R1_reg_9_ ( .D(Wt[9]), .RN(n626), .CK(clk), .Q(R1[9]) );
  DFFTRX1 R1_reg_7_ ( .D(Wt[7]), .RN(n623), .CK(clk), .Q(R1[7]) );
  DFFTRX1 counter1_reg_5_ ( .D(N1467), .RN(n2089), .CK(clk), .Q(counter1[5]), 
        .QN(n1054) );
  DFFHQX1 Wt_reg_17_ ( .D(N2148), .CK(clk), .Q(Wt[17]) );
  DFFTRX1 counter1_reg_3_ ( .D(N1465), .RN(n2089), .CK(clk), .Q(counter1[3])
         );
  DFFTRX1 counter1_reg_4_ ( .D(N1466), .RN(n2089), .CK(clk), .Q(counter1[4])
         );
  DFFTRX1 R15_reg_13_ ( .D(R14[13]), .RN(n630), .CK(clk), .Q(R15[13]) );
  DFFTRX1 R15_reg_11_ ( .D(R14[11]), .RN(n627), .CK(clk), .Q(R15[11]) );
  DFFTRX1 R6_reg_17_ ( .D(R5[17]), .RN(n636), .CK(clk), .Q(R6[17]) );
  DFFTRX1 R6_reg_15_ ( .D(R5[15]), .RN(n633), .CK(clk), .Q(R6[15]) );
  DFFTRX1 R6_reg_14_ ( .D(R5[14]), .RN(n632), .CK(clk), .Q(R6[14]) );
  DFFTRX1 R6_reg_11_ ( .D(R5[11]), .RN(n628), .CK(clk), .Q(R6[11]) );
  DFFTRX1 R6_reg_10_ ( .D(R5[10]), .RN(n627), .CK(clk), .Q(R6[10]) );
  DFFTRX1 R14_reg_2_ ( .D(R13[2]), .RN(n616), .CK(clk), .Q(R14[2]) );
  DFFTRX1 R15_reg_12_ ( .D(R14[12]), .RN(n629), .CK(clk), .Q(R15[12]) );
  DFFTRX1 R1_reg_6_ ( .D(Wt[6]), .RN(n622), .CK(clk), .Q(R1[6]) );
  DFFTRX1 R1_reg_5_ ( .D(Wt[5]), .RN(n621), .CK(clk), .Q(R1[5]) );
  DFFTRX1 R1_reg_4_ ( .D(Wt[4]), .RN(n620), .CK(clk), .Q(R1[4]) );
  DFFTRX1 R1_reg_3_ ( .D(Wt[3]), .RN(n618), .CK(clk), .Q(R1[3]) );
  DFFTRX1 R1_reg_8_ ( .D(Wt[8]), .RN(n625), .CK(clk), .Q(R1[8]) );
  DFFHQX1 Wt_reg_11_ ( .D(N2142), .CK(clk), .Q(Wt[11]) );
  DFFHQX1 Wt_reg_8_ ( .D(N2139), .CK(clk), .Q(Wt[8]) );
  DFFTRX1 R6_reg_12_ ( .D(R5[12]), .RN(n629), .CK(clk), .Q(R6[12]) );
  DFFTRX1 R15_reg_7_ ( .D(R14[7]), .RN(n622), .CK(clk), .Q(R15[7]) );
  DFFTRX1 R15_reg_3_ ( .D(R14[3]), .RN(n617), .CK(clk), .Q(R15[3]) );
  DFFTRX1 R15_reg_2_ ( .D(R14[2]), .RN(n616), .CK(clk), .Q(R15[2]) );
  DFFTRX1 R14_reg_0_ ( .D(R13[0]), .RN(n614), .CK(clk), .Q(R14[0]) );
  DFFTRX1 R1_reg_14_ ( .D(Wt[14]), .RN(n632), .CK(clk), .Q(R1[14]) );
  DFFTRX1 R2_reg_31_ ( .D(R1[31]), .RN(n653), .CK(clk), .Q(R2[31]) );
  DFFTRX1 R3_reg_31_ ( .D(R2[31]), .RN(n653), .CK(clk), .Q(R3[31]) );
  DFFTRX1 R4_reg_31_ ( .D(R3[31]), .RN(n653), .CK(clk), .Q(R4[31]) );
  DFFTRX1 R5_reg_31_ ( .D(R4[31]), .RN(n653), .CK(clk), .Q(R5[31]) );
  DFFTRX1 R7_reg_31_ ( .D(R6[31]), .RN(n653), .CK(clk), .Q(R7[31]) );
  DFFTRX1 R8_reg_31_ ( .D(R7[31]), .RN(n653), .CK(clk), .Q(R8[31]) );
  DFFTRX1 R9_reg_31_ ( .D(R8[31]), .RN(n653), .CK(clk), .Q(R9[31]) );
  DFFTRX1 R10_reg_31_ ( .D(R9[31]), .RN(n653), .CK(clk), .Q(R10[31]) );
  DFFTRX1 R11_reg_31_ ( .D(R10[31]), .RN(n653), .CK(clk), .Q(R11[31]) );
  DFFTRX1 R12_reg_31_ ( .D(R11[31]), .RN(n653), .CK(clk), .Q(R12[31]) );
  DFFTRX1 R13_reg_31_ ( .D(R12[31]), .RN(n652), .CK(clk), .Q(R13[31]) );
  DFFTRX1 R2_reg_30_ ( .D(R1[30]), .RN(n652), .CK(clk), .Q(R2[30]) );
  DFFTRX1 R3_reg_30_ ( .D(R2[30]), .RN(n652), .CK(clk), .Q(R3[30]) );
  DFFTRX1 R4_reg_30_ ( .D(R3[30]), .RN(n652), .CK(clk), .Q(R4[30]) );
  DFFTRX1 R5_reg_30_ ( .D(R4[30]), .RN(n652), .CK(clk), .Q(R5[30]) );
  DFFTRX1 R7_reg_30_ ( .D(R6[30]), .RN(n652), .CK(clk), .Q(R7[30]) );
  DFFTRX1 R8_reg_30_ ( .D(R7[30]), .RN(n652), .CK(clk), .Q(R8[30]) );
  DFFTRX1 R9_reg_30_ ( .D(R8[30]), .RN(n652), .CK(clk), .Q(R9[30]) );
  DFFTRX1 R10_reg_30_ ( .D(R9[30]), .RN(n651), .CK(clk), .Q(R10[30]) );
  DFFTRX1 R11_reg_30_ ( .D(R10[30]), .RN(n651), .CK(clk), .Q(R11[30]) );
  DFFTRX1 R12_reg_30_ ( .D(R11[30]), .RN(n651), .CK(clk), .Q(R12[30]) );
  DFFTRX1 R13_reg_30_ ( .D(R12[30]), .RN(n651), .CK(clk), .Q(R13[30]) );
  DFFTRX1 R2_reg_29_ ( .D(R1[29]), .RN(n651), .CK(clk), .Q(R2[29]) );
  DFFTRX1 R3_reg_29_ ( .D(R2[29]), .RN(n651), .CK(clk), .Q(R3[29]) );
  DFFTRX1 R4_reg_29_ ( .D(R3[29]), .RN(n651), .CK(clk), .Q(R4[29]) );
  DFFTRX1 R5_reg_29_ ( .D(R4[29]), .RN(n651), .CK(clk), .Q(R5[29]) );
  DFFTRX1 R7_reg_29_ ( .D(R6[29]), .RN(n650), .CK(clk), .Q(R7[29]) );
  DFFTRX1 R8_reg_29_ ( .D(R7[29]), .RN(n650), .CK(clk), .Q(R8[29]) );
  DFFTRX1 R9_reg_29_ ( .D(R8[29]), .RN(n650), .CK(clk), .Q(R9[29]) );
  DFFTRX1 R10_reg_29_ ( .D(R9[29]), .RN(n650), .CK(clk), .Q(R10[29]) );
  DFFTRX1 R11_reg_29_ ( .D(R10[29]), .RN(n650), .CK(clk), .Q(R11[29]) );
  DFFTRX1 R12_reg_29_ ( .D(R11[29]), .RN(n650), .CK(clk), .Q(R12[29]) );
  DFFTRX1 R13_reg_29_ ( .D(R12[29]), .RN(n650), .CK(clk), .Q(R13[29]) );
  DFFTRX1 R2_reg_28_ ( .D(R1[28]), .RN(n650), .CK(clk), .Q(R2[28]) );
  DFFTRX1 R3_reg_28_ ( .D(R2[28]), .RN(n650), .CK(clk), .Q(R3[28]) );
  DFFTRX1 R4_reg_28_ ( .D(R3[28]), .RN(n649), .CK(clk), .Q(R4[28]) );
  DFFTRX1 R5_reg_28_ ( .D(R4[28]), .RN(n649), .CK(clk), .Q(R5[28]) );
  DFFTRX1 R7_reg_28_ ( .D(R6[28]), .RN(n649), .CK(clk), .Q(R7[28]) );
  DFFTRX1 R8_reg_28_ ( .D(R7[28]), .RN(n649), .CK(clk), .Q(R8[28]) );
  DFFTRX1 R9_reg_28_ ( .D(R8[28]), .RN(n649), .CK(clk), .Q(R9[28]) );
  DFFTRX1 R10_reg_28_ ( .D(R9[28]), .RN(n649), .CK(clk), .Q(R10[28]) );
  DFFTRX1 R11_reg_28_ ( .D(R10[28]), .RN(n649), .CK(clk), .Q(R11[28]) );
  DFFTRX1 R12_reg_28_ ( .D(R11[28]), .RN(n649), .CK(clk), .Q(R12[28]) );
  DFFTRX1 R13_reg_28_ ( .D(R12[28]), .RN(n649), .CK(clk), .Q(R13[28]) );
  DFFTRX1 R2_reg_27_ ( .D(R1[27]), .RN(n648), .CK(clk), .Q(R2[27]) );
  DFFTRX1 R3_reg_27_ ( .D(R2[27]), .RN(n648), .CK(clk), .Q(R3[27]) );
  DFFTRX1 R4_reg_27_ ( .D(R3[27]), .RN(n648), .CK(clk), .Q(R4[27]) );
  DFFTRX1 R5_reg_27_ ( .D(R4[27]), .RN(n648), .CK(clk), .Q(R5[27]) );
  DFFTRX1 R7_reg_27_ ( .D(R6[27]), .RN(n648), .CK(clk), .Q(R7[27]) );
  DFFTRX1 R8_reg_27_ ( .D(R7[27]), .RN(n648), .CK(clk), .Q(R8[27]) );
  DFFTRX1 R9_reg_27_ ( .D(R8[27]), .RN(n648), .CK(clk), .Q(R9[27]) );
  DFFTRX1 R10_reg_27_ ( .D(R9[27]), .RN(n648), .CK(clk), .Q(R10[27]) );
  DFFTRX1 R11_reg_27_ ( .D(R10[27]), .RN(n648), .CK(clk), .Q(R11[27]) );
  DFFTRX1 R12_reg_27_ ( .D(R11[27]), .RN(n648), .CK(clk), .Q(R12[27]) );
  DFFTRX1 R13_reg_27_ ( .D(R12[27]), .RN(n647), .CK(clk), .Q(R13[27]) );
  DFFTRX1 R2_reg_26_ ( .D(R1[26]), .RN(n647), .CK(clk), .Q(R2[26]) );
  DFFTRX1 R3_reg_26_ ( .D(R2[26]), .RN(n647), .CK(clk), .Q(R3[26]) );
  DFFTRX1 R4_reg_26_ ( .D(R3[26]), .RN(n647), .CK(clk), .Q(R4[26]) );
  DFFTRX1 R5_reg_26_ ( .D(R4[26]), .RN(n647), .CK(clk), .Q(R5[26]) );
  DFFTRX1 R7_reg_26_ ( .D(R6[26]), .RN(n647), .CK(clk), .Q(R7[26]) );
  DFFTRX1 R8_reg_26_ ( .D(R7[26]), .RN(n647), .CK(clk), .Q(R8[26]) );
  DFFTRX1 R9_reg_26_ ( .D(R8[26]), .RN(n647), .CK(clk), .Q(R9[26]) );
  DFFTRX1 R10_reg_26_ ( .D(R9[26]), .RN(n646), .CK(clk), .Q(R10[26]) );
  DFFTRX1 R11_reg_26_ ( .D(R10[26]), .RN(n646), .CK(clk), .Q(R11[26]) );
  DFFTRX1 R12_reg_26_ ( .D(R11[26]), .RN(n646), .CK(clk), .Q(R12[26]) );
  DFFTRX1 R13_reg_26_ ( .D(R12[26]), .RN(n646), .CK(clk), .Q(R13[26]) );
  DFFTRX1 R2_reg_25_ ( .D(R1[25]), .RN(n646), .CK(clk), .Q(R2[25]) );
  DFFTRX1 R3_reg_25_ ( .D(R2[25]), .RN(n646), .CK(clk), .Q(R3[25]) );
  DFFTRX1 R4_reg_25_ ( .D(R3[25]), .RN(n646), .CK(clk), .Q(R4[25]) );
  DFFTRX1 R5_reg_25_ ( .D(R4[25]), .RN(n646), .CK(clk), .Q(R5[25]) );
  DFFTRX1 R7_reg_25_ ( .D(R6[25]), .RN(n645), .CK(clk), .Q(R7[25]) );
  DFFTRX1 R8_reg_25_ ( .D(R7[25]), .RN(n645), .CK(clk), .Q(R8[25]) );
  DFFTRX1 R9_reg_25_ ( .D(R8[25]), .RN(n645), .CK(clk), .Q(R9[25]) );
  DFFTRX1 R10_reg_25_ ( .D(R9[25]), .RN(n645), .CK(clk), .Q(R10[25]) );
  DFFTRX1 R11_reg_25_ ( .D(R10[25]), .RN(n645), .CK(clk), .Q(R11[25]) );
  DFFTRX1 R12_reg_25_ ( .D(R11[25]), .RN(n645), .CK(clk), .Q(R12[25]) );
  DFFTRX1 R13_reg_25_ ( .D(R12[25]), .RN(n645), .CK(clk), .Q(R13[25]) );
  DFFTRX1 R2_reg_24_ ( .D(R1[24]), .RN(n645), .CK(clk), .Q(R2[24]) );
  DFFTRX1 R3_reg_24_ ( .D(R2[24]), .RN(n645), .CK(clk), .Q(R3[24]) );
  DFFTRX1 R4_reg_24_ ( .D(R3[24]), .RN(n644), .CK(clk), .Q(R4[24]) );
  DFFTRX1 R5_reg_24_ ( .D(R4[24]), .RN(n644), .CK(clk), .Q(R5[24]) );
  DFFTRX1 R7_reg_24_ ( .D(R6[24]), .RN(n644), .CK(clk), .Q(R7[24]) );
  DFFTRX1 R8_reg_24_ ( .D(R7[24]), .RN(n644), .CK(clk), .Q(R8[24]) );
  DFFTRX1 R9_reg_24_ ( .D(R8[24]), .RN(n644), .CK(clk), .Q(R9[24]) );
  DFFTRX1 R10_reg_24_ ( .D(R9[24]), .RN(n644), .CK(clk), .Q(R10[24]) );
  DFFTRX1 R11_reg_24_ ( .D(R10[24]), .RN(n644), .CK(clk), .Q(R11[24]) );
  DFFTRX1 R12_reg_24_ ( .D(R11[24]), .RN(n644), .CK(clk), .Q(R12[24]) );
  DFFTRX1 R13_reg_24_ ( .D(R12[24]), .RN(n644), .CK(clk), .Q(R13[24]) );
  DFFTRX1 R2_reg_23_ ( .D(R1[23]), .RN(n643), .CK(clk), .Q(R2[23]) );
  DFFTRX1 R3_reg_23_ ( .D(R2[23]), .RN(n643), .CK(clk), .Q(R3[23]) );
  DFFTRX1 R4_reg_23_ ( .D(R3[23]), .RN(n643), .CK(clk), .Q(R4[23]) );
  DFFTRX1 R5_reg_23_ ( .D(R4[23]), .RN(n643), .CK(clk), .Q(R5[23]) );
  DFFTRX1 R7_reg_23_ ( .D(R6[23]), .RN(n643), .CK(clk), .Q(R7[23]) );
  DFFTRX1 R8_reg_23_ ( .D(R7[23]), .RN(n643), .CK(clk), .Q(R8[23]) );
  DFFTRX1 R9_reg_23_ ( .D(R8[23]), .RN(n643), .CK(clk), .Q(R9[23]) );
  DFFTRX1 R10_reg_23_ ( .D(R9[23]), .RN(n643), .CK(clk), .Q(R10[23]) );
  DFFTRX1 R11_reg_23_ ( .D(R10[23]), .RN(n643), .CK(clk), .Q(R11[23]) );
  DFFTRX1 R12_reg_23_ ( .D(R11[23]), .RN(n643), .CK(clk), .Q(R12[23]) );
  DFFTRX1 R13_reg_23_ ( .D(R12[23]), .RN(n642), .CK(clk), .Q(R13[23]) );
  DFFTRX1 R2_reg_22_ ( .D(R1[22]), .RN(n642), .CK(clk), .Q(R2[22]) );
  DFFTRX1 R3_reg_22_ ( .D(R2[22]), .RN(n642), .CK(clk), .Q(R3[22]) );
  DFFTRX1 R4_reg_22_ ( .D(R3[22]), .RN(n642), .CK(clk), .Q(R4[22]) );
  DFFTRX1 R5_reg_22_ ( .D(R4[22]), .RN(n642), .CK(clk), .Q(R5[22]) );
  DFFTRX1 R7_reg_22_ ( .D(R6[22]), .RN(n642), .CK(clk), .Q(R7[22]) );
  DFFTRX1 R8_reg_22_ ( .D(R7[22]), .RN(n642), .CK(clk), .Q(R8[22]) );
  DFFTRX1 R9_reg_22_ ( .D(R8[22]), .RN(n642), .CK(clk), .Q(R9[22]) );
  DFFTRX1 R10_reg_22_ ( .D(R9[22]), .RN(n641), .CK(clk), .Q(R10[22]) );
  DFFTRX1 R11_reg_22_ ( .D(R10[22]), .RN(n641), .CK(clk), .Q(R11[22]) );
  DFFTRX1 R12_reg_22_ ( .D(R11[22]), .RN(n641), .CK(clk), .Q(R12[22]) );
  DFFTRX1 R13_reg_22_ ( .D(R12[22]), .RN(n641), .CK(clk), .Q(R13[22]) );
  DFFTRX1 R2_reg_21_ ( .D(R1[21]), .RN(n641), .CK(clk), .Q(R2[21]) );
  DFFTRX1 R3_reg_21_ ( .D(R2[21]), .RN(n641), .CK(clk), .Q(R3[21]) );
  DFFTRX1 R4_reg_21_ ( .D(R3[21]), .RN(n641), .CK(clk), .Q(R4[21]) );
  DFFTRX1 R5_reg_21_ ( .D(R4[21]), .RN(n641), .CK(clk), .Q(R5[21]) );
  DFFTRX1 R7_reg_21_ ( .D(R6[21]), .RN(n640), .CK(clk), .Q(R7[21]) );
  DFFTRX1 R8_reg_21_ ( .D(R7[21]), .RN(n640), .CK(clk), .Q(R8[21]) );
  DFFTRX1 R9_reg_21_ ( .D(R8[21]), .RN(n640), .CK(clk), .Q(R9[21]) );
  DFFTRX1 R10_reg_21_ ( .D(R9[21]), .RN(n640), .CK(clk), .Q(R10[21]) );
  DFFTRX1 R11_reg_21_ ( .D(R10[21]), .RN(n640), .CK(clk), .Q(R11[21]) );
  DFFTRX1 R12_reg_21_ ( .D(R11[21]), .RN(n640), .CK(clk), .Q(R12[21]) );
  DFFTRX1 R13_reg_21_ ( .D(R12[21]), .RN(n640), .CK(clk), .Q(R13[21]) );
  DFFTRX1 R2_reg_20_ ( .D(R1[20]), .RN(n640), .CK(clk), .Q(R2[20]) );
  DFFTRX1 R3_reg_20_ ( .D(R2[20]), .RN(n640), .CK(clk), .Q(R3[20]) );
  DFFTRX1 R4_reg_20_ ( .D(R3[20]), .RN(n639), .CK(clk), .Q(R4[20]) );
  DFFTRX1 R5_reg_20_ ( .D(R4[20]), .RN(n639), .CK(clk), .Q(R5[20]) );
  DFFTRX1 R7_reg_20_ ( .D(R6[20]), .RN(n639), .CK(clk), .Q(R7[20]) );
  DFFTRX1 R8_reg_20_ ( .D(R7[20]), .RN(n639), .CK(clk), .Q(R8[20]) );
  DFFTRX1 R9_reg_20_ ( .D(R8[20]), .RN(n639), .CK(clk), .Q(R9[20]) );
  DFFTRX1 R10_reg_20_ ( .D(R9[20]), .RN(n639), .CK(clk), .Q(R10[20]) );
  DFFTRX1 R11_reg_20_ ( .D(R10[20]), .RN(n639), .CK(clk), .Q(R11[20]) );
  DFFTRX1 R12_reg_20_ ( .D(R11[20]), .RN(n639), .CK(clk), .Q(R12[20]) );
  DFFTRX1 R13_reg_20_ ( .D(R12[20]), .RN(n639), .CK(clk), .Q(R13[20]) );
  DFFTRX1 R2_reg_19_ ( .D(R1[19]), .RN(n638), .CK(clk), .Q(R2[19]) );
  DFFTRX1 R3_reg_19_ ( .D(R2[19]), .RN(n638), .CK(clk), .Q(R3[19]) );
  DFFTRX1 R4_reg_19_ ( .D(R3[19]), .RN(n638), .CK(clk), .Q(R4[19]) );
  DFFTRX1 R5_reg_19_ ( .D(R4[19]), .RN(n638), .CK(clk), .Q(R5[19]) );
  DFFTRX1 R7_reg_19_ ( .D(R6[19]), .RN(n638), .CK(clk), .Q(R7[19]) );
  DFFTRX1 R8_reg_19_ ( .D(R7[19]), .RN(n638), .CK(clk), .Q(R8[19]) );
  DFFTRX1 R9_reg_19_ ( .D(R8[19]), .RN(n638), .CK(clk), .Q(R9[19]) );
  DFFTRX1 R10_reg_19_ ( .D(R9[19]), .RN(n638), .CK(clk), .Q(R10[19]) );
  DFFTRX1 R11_reg_19_ ( .D(R10[19]), .RN(n638), .CK(clk), .Q(R11[19]) );
  DFFTRX1 R12_reg_19_ ( .D(R11[19]), .RN(n638), .CK(clk), .Q(R12[19]) );
  DFFTRX1 R13_reg_19_ ( .D(R12[19]), .RN(n637), .CK(clk), .Q(R13[19]) );
  DFFTRX1 R2_reg_18_ ( .D(R1[18]), .RN(n637), .CK(clk), .Q(R2[18]) );
  DFFTRX1 R3_reg_18_ ( .D(R2[18]), .RN(n637), .CK(clk), .Q(R3[18]) );
  DFFTRX1 R4_reg_18_ ( .D(R3[18]), .RN(n637), .CK(clk), .Q(R4[18]) );
  DFFTRX1 R5_reg_18_ ( .D(R4[18]), .RN(n637), .CK(clk), .Q(R5[18]) );
  DFFTRX1 R7_reg_18_ ( .D(R6[18]), .RN(n637), .CK(clk), .Q(R7[18]) );
  DFFTRX1 R8_reg_18_ ( .D(R7[18]), .RN(n637), .CK(clk), .Q(R8[18]) );
  DFFTRX1 R9_reg_18_ ( .D(R8[18]), .RN(n637), .CK(clk), .Q(R9[18]) );
  DFFTRX1 R10_reg_18_ ( .D(R9[18]), .RN(n636), .CK(clk), .Q(R10[18]) );
  DFFTRX1 R11_reg_18_ ( .D(R10[18]), .RN(n636), .CK(clk), .Q(R11[18]) );
  DFFTRX1 R12_reg_18_ ( .D(R11[18]), .RN(n636), .CK(clk), .Q(R12[18]) );
  DFFTRX1 R13_reg_18_ ( .D(R12[18]), .RN(n636), .CK(clk), .Q(R13[18]) );
  DFFTRX1 R2_reg_17_ ( .D(R1[17]), .RN(n636), .CK(clk), .Q(R2[17]) );
  DFFTRX1 R3_reg_17_ ( .D(R2[17]), .RN(n636), .CK(clk), .Q(R3[17]) );
  DFFTRX1 R4_reg_17_ ( .D(R3[17]), .RN(n636), .CK(clk), .Q(R4[17]) );
  DFFTRX1 R5_reg_17_ ( .D(R4[17]), .RN(n636), .CK(clk), .Q(R5[17]) );
  DFFTRX1 R7_reg_17_ ( .D(R6[17]), .RN(n635), .CK(clk), .Q(R7[17]) );
  DFFTRX1 R8_reg_17_ ( .D(R7[17]), .RN(n635), .CK(clk), .Q(R8[17]) );
  DFFTRX1 R9_reg_17_ ( .D(R8[17]), .RN(n635), .CK(clk), .Q(R9[17]) );
  DFFTRX1 R10_reg_17_ ( .D(R9[17]), .RN(n635), .CK(clk), .Q(R10[17]) );
  DFFTRX1 R11_reg_17_ ( .D(R10[17]), .RN(n635), .CK(clk), .Q(R11[17]) );
  DFFTRX1 R12_reg_17_ ( .D(R11[17]), .RN(n635), .CK(clk), .Q(R12[17]) );
  DFFTRX1 R13_reg_17_ ( .D(R12[17]), .RN(n635), .CK(clk), .Q(R13[17]) );
  DFFTRX1 R2_reg_16_ ( .D(R1[16]), .RN(n635), .CK(clk), .Q(R2[16]) );
  DFFTRX1 R3_reg_16_ ( .D(R2[16]), .RN(n635), .CK(clk), .Q(R3[16]) );
  DFFTRX1 R4_reg_16_ ( .D(R3[16]), .RN(n634), .CK(clk), .Q(R4[16]) );
  DFFTRX1 R5_reg_16_ ( .D(R4[16]), .RN(n634), .CK(clk), .Q(R5[16]) );
  DFFTRX1 R7_reg_16_ ( .D(R6[16]), .RN(n634), .CK(clk), .Q(R7[16]) );
  DFFTRX1 R8_reg_16_ ( .D(R7[16]), .RN(n634), .CK(clk), .Q(R8[16]) );
  DFFTRX1 R9_reg_16_ ( .D(R8[16]), .RN(n634), .CK(clk), .Q(R9[16]) );
  DFFTRX1 R10_reg_16_ ( .D(R9[16]), .RN(n634), .CK(clk), .Q(R10[16]) );
  DFFTRX1 R11_reg_16_ ( .D(R10[16]), .RN(n634), .CK(clk), .Q(R11[16]) );
  DFFTRX1 R12_reg_16_ ( .D(R11[16]), .RN(n634), .CK(clk), .Q(R12[16]) );
  DFFTRX1 R13_reg_16_ ( .D(R12[16]), .RN(n634), .CK(clk), .Q(R13[16]) );
  DFFTRX1 R2_reg_15_ ( .D(R1[15]), .RN(n633), .CK(clk), .Q(R2[15]) );
  DFFTRX1 R3_reg_15_ ( .D(R2[15]), .RN(n633), .CK(clk), .Q(R3[15]) );
  DFFTRX1 R4_reg_15_ ( .D(R3[15]), .RN(n633), .CK(clk), .Q(R4[15]) );
  DFFTRX1 R5_reg_15_ ( .D(R4[15]), .RN(n633), .CK(clk), .Q(R5[15]) );
  DFFTRX1 R7_reg_15_ ( .D(R6[15]), .RN(n633), .CK(clk), .Q(R7[15]) );
  DFFTRX1 R8_reg_15_ ( .D(R7[15]), .RN(n633), .CK(clk), .Q(R8[15]) );
  DFFTRX1 R9_reg_15_ ( .D(R8[15]), .RN(n633), .CK(clk), .Q(R9[15]) );
  DFFTRX1 R10_reg_15_ ( .D(R9[15]), .RN(n633), .CK(clk), .Q(R10[15]) );
  DFFTRX1 R11_reg_15_ ( .D(R10[15]), .RN(n633), .CK(clk), .Q(R11[15]) );
  DFFTRX1 R12_reg_15_ ( .D(R11[15]), .RN(n633), .CK(clk), .Q(R12[15]) );
  DFFTRX1 R13_reg_15_ ( .D(R12[15]), .RN(n632), .CK(clk), .Q(R13[15]) );
  DFFTRX1 R2_reg_14_ ( .D(R1[14]), .RN(n632), .CK(clk), .Q(R2[14]) );
  DFFTRX1 R3_reg_14_ ( .D(R2[14]), .RN(n632), .CK(clk), .Q(R3[14]) );
  DFFTRX1 R4_reg_14_ ( .D(R3[14]), .RN(n632), .CK(clk), .Q(R4[14]) );
  DFFTRX1 R5_reg_14_ ( .D(R4[14]), .RN(n632), .CK(clk), .Q(R5[14]) );
  DFFTRX1 R7_reg_14_ ( .D(R6[14]), .RN(n632), .CK(clk), .Q(R7[14]) );
  DFFTRX1 R8_reg_14_ ( .D(R7[14]), .RN(n632), .CK(clk), .Q(R8[14]) );
  DFFTRX1 R9_reg_14_ ( .D(R8[14]), .RN(n632), .CK(clk), .Q(R9[14]) );
  DFFTRX1 R10_reg_14_ ( .D(R9[14]), .RN(n631), .CK(clk), .Q(R10[14]) );
  DFFTRX1 R11_reg_14_ ( .D(R10[14]), .RN(n631), .CK(clk), .Q(R11[14]) );
  DFFTRX1 R12_reg_14_ ( .D(R11[14]), .RN(n631), .CK(clk), .Q(R12[14]) );
  DFFTRX1 R13_reg_14_ ( .D(R12[14]), .RN(n631), .CK(clk), .Q(R13[14]) );
  DFFTRX1 R2_reg_13_ ( .D(R1[13]), .RN(n631), .CK(clk), .Q(R2[13]) );
  DFFTRX1 R3_reg_13_ ( .D(R2[13]), .RN(n631), .CK(clk), .Q(R3[13]) );
  DFFTRX1 R4_reg_13_ ( .D(R3[13]), .RN(n631), .CK(clk), .Q(R4[13]) );
  DFFTRX1 R5_reg_13_ ( .D(R4[13]), .RN(n631), .CK(clk), .Q(R5[13]) );
  DFFTRX1 R7_reg_13_ ( .D(R6[13]), .RN(n630), .CK(clk), .Q(R7[13]) );
  DFFTRX1 R8_reg_13_ ( .D(R7[13]), .RN(n630), .CK(clk), .Q(R8[13]) );
  DFFTRX1 R9_reg_13_ ( .D(R8[13]), .RN(n630), .CK(clk), .Q(R9[13]) );
  DFFTRX1 R10_reg_13_ ( .D(R9[13]), .RN(n630), .CK(clk), .Q(R10[13]) );
  DFFTRX1 R11_reg_13_ ( .D(R10[13]), .RN(n630), .CK(clk), .Q(R11[13]) );
  DFFTRX1 R12_reg_13_ ( .D(R11[13]), .RN(n630), .CK(clk), .Q(R12[13]) );
  DFFTRX1 R13_reg_13_ ( .D(R12[13]), .RN(n630), .CK(clk), .Q(R13[13]) );
  DFFTRX1 R2_reg_12_ ( .D(R1[12]), .RN(n630), .CK(clk), .Q(R2[12]) );
  DFFTRX1 R3_reg_12_ ( .D(R2[12]), .RN(n630), .CK(clk), .Q(R3[12]) );
  DFFTRX1 R4_reg_12_ ( .D(R3[12]), .RN(n629), .CK(clk), .Q(R4[12]) );
  DFFTRX1 R5_reg_12_ ( .D(R4[12]), .RN(n629), .CK(clk), .Q(R5[12]) );
  DFFTRX1 R7_reg_12_ ( .D(R6[12]), .RN(n629), .CK(clk), .Q(R7[12]) );
  DFFTRX1 R8_reg_12_ ( .D(R7[12]), .RN(n629), .CK(clk), .Q(R8[12]) );
  DFFTRX1 R9_reg_12_ ( .D(R8[12]), .RN(n629), .CK(clk), .Q(R9[12]) );
  DFFTRX1 R10_reg_12_ ( .D(R9[12]), .RN(n629), .CK(clk), .Q(R10[12]) );
  DFFTRX1 R11_reg_12_ ( .D(R10[12]), .RN(n629), .CK(clk), .Q(R11[12]) );
  DFFTRX1 R12_reg_12_ ( .D(R11[12]), .RN(n629), .CK(clk), .Q(R12[12]) );
  DFFTRX1 R13_reg_12_ ( .D(R12[12]), .RN(n629), .CK(clk), .Q(R13[12]) );
  DFFTRX1 R2_reg_11_ ( .D(R1[11]), .RN(n628), .CK(clk), .Q(R2[11]) );
  DFFTRX1 R3_reg_11_ ( .D(R2[11]), .RN(n628), .CK(clk), .Q(R3[11]) );
  DFFTRX1 R4_reg_11_ ( .D(R3[11]), .RN(n628), .CK(clk), .Q(R4[11]) );
  DFFTRX1 R5_reg_11_ ( .D(R4[11]), .RN(n628), .CK(clk), .Q(R5[11]) );
  DFFTRX1 R7_reg_11_ ( .D(R6[11]), .RN(n628), .CK(clk), .Q(R7[11]) );
  DFFTRX1 R8_reg_11_ ( .D(R7[11]), .RN(n628), .CK(clk), .Q(R8[11]) );
  DFFTRX1 R9_reg_11_ ( .D(R8[11]), .RN(n628), .CK(clk), .Q(R9[11]) );
  DFFTRX1 R10_reg_11_ ( .D(R9[11]), .RN(n628), .CK(clk), .Q(R10[11]) );
  DFFTRX1 R11_reg_11_ ( .D(R10[11]), .RN(n628), .CK(clk), .Q(R11[11]) );
  DFFTRX1 R12_reg_11_ ( .D(R11[11]), .RN(n628), .CK(clk), .Q(R12[11]) );
  DFFTRX1 R13_reg_11_ ( .D(R12[11]), .RN(n627), .CK(clk), .Q(R13[11]) );
  DFFTRX1 R2_reg_10_ ( .D(R1[10]), .RN(n627), .CK(clk), .Q(R2[10]) );
  DFFTRX1 R3_reg_10_ ( .D(R2[10]), .RN(n627), .CK(clk), .Q(R3[10]) );
  DFFTRX1 R4_reg_10_ ( .D(R3[10]), .RN(n627), .CK(clk), .Q(R4[10]) );
  DFFTRX1 R5_reg_10_ ( .D(R4[10]), .RN(n627), .CK(clk), .Q(R5[10]) );
  DFFTRX1 R7_reg_10_ ( .D(R6[10]), .RN(n627), .CK(clk), .Q(R7[10]) );
  DFFTRX1 R8_reg_10_ ( .D(R7[10]), .RN(n627), .CK(clk), .Q(R8[10]) );
  DFFTRX1 R9_reg_10_ ( .D(R8[10]), .RN(n627), .CK(clk), .Q(R9[10]) );
  DFFTRX1 R10_reg_10_ ( .D(R9[10]), .RN(n626), .CK(clk), .Q(R10[10]) );
  DFFTRX1 R11_reg_10_ ( .D(R10[10]), .RN(n626), .CK(clk), .Q(R11[10]) );
  DFFTRX1 R12_reg_10_ ( .D(R11[10]), .RN(n626), .CK(clk), .Q(R12[10]) );
  DFFTRX1 R13_reg_10_ ( .D(R12[10]), .RN(n626), .CK(clk), .Q(R13[10]) );
  DFFTRX1 R2_reg_9_ ( .D(R1[9]), .RN(n626), .CK(clk), .Q(R2[9]) );
  DFFTRX1 R3_reg_9_ ( .D(R2[9]), .RN(n626), .CK(clk), .Q(R3[9]) );
  DFFTRX1 R4_reg_9_ ( .D(R3[9]), .RN(n626), .CK(clk), .Q(R4[9]) );
  DFFTRX1 R5_reg_9_ ( .D(R4[9]), .RN(n626), .CK(clk), .Q(R5[9]) );
  DFFTRX1 R7_reg_9_ ( .D(R6[9]), .RN(n625), .CK(clk), .Q(R7[9]) );
  DFFTRX1 R8_reg_9_ ( .D(R7[9]), .RN(n625), .CK(clk), .Q(R8[9]) );
  DFFTRX1 R9_reg_9_ ( .D(R8[9]), .RN(n625), .CK(clk), .Q(R9[9]) );
  DFFTRX1 R10_reg_9_ ( .D(R9[9]), .RN(n625), .CK(clk), .Q(R10[9]) );
  DFFTRX1 R11_reg_9_ ( .D(R10[9]), .RN(n625), .CK(clk), .Q(R11[9]) );
  DFFTRX1 R12_reg_9_ ( .D(R11[9]), .RN(n625), .CK(clk), .Q(R12[9]) );
  DFFTRX1 R13_reg_9_ ( .D(R12[9]), .RN(n625), .CK(clk), .Q(R13[9]) );
  DFFTRX1 R2_reg_8_ ( .D(R1[8]), .RN(n625), .CK(clk), .Q(R2[8]) );
  DFFTRX1 R3_reg_8_ ( .D(R2[8]), .RN(n625), .CK(clk), .Q(R3[8]) );
  DFFTRX1 R4_reg_8_ ( .D(R3[8]), .RN(n624), .CK(clk), .Q(R4[8]) );
  DFFTRX1 R5_reg_8_ ( .D(R4[8]), .RN(n624), .CK(clk), .Q(R5[8]) );
  DFFTRX1 R7_reg_8_ ( .D(R6[8]), .RN(n624), .CK(clk), .Q(R7[8]) );
  DFFTRX1 R8_reg_8_ ( .D(R7[8]), .RN(n624), .CK(clk), .Q(R8[8]) );
  DFFTRX1 R9_reg_8_ ( .D(R8[8]), .RN(n624), .CK(clk), .Q(R9[8]) );
  DFFTRX1 R10_reg_8_ ( .D(R9[8]), .RN(n624), .CK(clk), .Q(R10[8]) );
  DFFTRX1 R11_reg_8_ ( .D(R10[8]), .RN(n624), .CK(clk), .Q(R11[8]) );
  DFFTRX1 R12_reg_8_ ( .D(R11[8]), .RN(n624), .CK(clk), .Q(R12[8]) );
  DFFTRX1 R13_reg_8_ ( .D(R12[8]), .RN(n624), .CK(clk), .Q(R13[8]) );
  DFFTRX1 R2_reg_7_ ( .D(R1[7]), .RN(n623), .CK(clk), .Q(R2[7]) );
  DFFTRX1 R3_reg_7_ ( .D(R2[7]), .RN(n623), .CK(clk), .Q(R3[7]) );
  DFFTRX1 R4_reg_7_ ( .D(R3[7]), .RN(n623), .CK(clk), .Q(R4[7]) );
  DFFTRX1 R5_reg_7_ ( .D(R4[7]), .RN(n623), .CK(clk), .Q(R5[7]) );
  DFFTRX1 R7_reg_7_ ( .D(R6[7]), .RN(n623), .CK(clk), .Q(R7[7]) );
  DFFTRX1 R8_reg_7_ ( .D(R7[7]), .RN(n623), .CK(clk), .Q(R8[7]) );
  DFFTRX1 R9_reg_7_ ( .D(R8[7]), .RN(n623), .CK(clk), .Q(R9[7]) );
  DFFTRX1 R10_reg_7_ ( .D(R9[7]), .RN(n623), .CK(clk), .Q(R10[7]) );
  DFFTRX1 R11_reg_7_ ( .D(R10[7]), .RN(n623), .CK(clk), .Q(R11[7]) );
  DFFTRX1 R12_reg_7_ ( .D(R11[7]), .RN(n623), .CK(clk), .Q(R12[7]) );
  DFFTRX1 R13_reg_7_ ( .D(R12[7]), .RN(n622), .CK(clk), .Q(R13[7]) );
  DFFTRX1 R2_reg_6_ ( .D(R1[6]), .RN(n622), .CK(clk), .Q(R2[6]) );
  DFFTRX1 R3_reg_6_ ( .D(R2[6]), .RN(n622), .CK(clk), .Q(R3[6]) );
  DFFTRX1 R4_reg_6_ ( .D(R3[6]), .RN(n622), .CK(clk), .Q(R4[6]) );
  DFFTRX1 R5_reg_6_ ( .D(R4[6]), .RN(n622), .CK(clk), .Q(R5[6]) );
  DFFTRX1 R7_reg_6_ ( .D(R6[6]), .RN(n622), .CK(clk), .Q(R7[6]) );
  DFFTRX1 R8_reg_6_ ( .D(R7[6]), .RN(n622), .CK(clk), .Q(R8[6]) );
  DFFTRX1 R9_reg_6_ ( .D(R8[6]), .RN(n622), .CK(clk), .Q(R9[6]) );
  DFFTRX1 R10_reg_6_ ( .D(R9[6]), .RN(n621), .CK(clk), .Q(R10[6]) );
  DFFTRX1 R11_reg_6_ ( .D(R10[6]), .RN(n621), .CK(clk), .Q(R11[6]) );
  DFFTRX1 R12_reg_6_ ( .D(R11[6]), .RN(n621), .CK(clk), .Q(R12[6]) );
  DFFTRX1 R13_reg_6_ ( .D(R12[6]), .RN(n621), .CK(clk), .Q(R13[6]) );
  DFFTRX1 R2_reg_5_ ( .D(R1[5]), .RN(n621), .CK(clk), .Q(R2[5]) );
  DFFTRX1 R3_reg_5_ ( .D(R2[5]), .RN(n621), .CK(clk), .Q(R3[5]) );
  DFFTRX1 R4_reg_5_ ( .D(R3[5]), .RN(n621), .CK(clk), .Q(R4[5]) );
  DFFTRX1 R5_reg_5_ ( .D(R4[5]), .RN(n621), .CK(clk), .Q(R5[5]) );
  DFFTRX1 R7_reg_5_ ( .D(R6[5]), .RN(n620), .CK(clk), .Q(R7[5]) );
  DFFTRX1 R8_reg_5_ ( .D(R7[5]), .RN(n620), .CK(clk), .Q(R8[5]) );
  DFFTRX1 R9_reg_5_ ( .D(R8[5]), .RN(n620), .CK(clk), .Q(R9[5]) );
  DFFTRX1 R10_reg_5_ ( .D(R9[5]), .RN(n620), .CK(clk), .Q(R10[5]) );
  DFFTRX1 R11_reg_5_ ( .D(R10[5]), .RN(n620), .CK(clk), .Q(R11[5]) );
  DFFTRX1 R12_reg_5_ ( .D(R11[5]), .RN(n620), .CK(clk), .Q(R12[5]) );
  DFFTRX1 R13_reg_5_ ( .D(R12[5]), .RN(n620), .CK(clk), .Q(R13[5]) );
  DFFTRX1 R2_reg_4_ ( .D(R1[4]), .RN(n620), .CK(clk), .Q(R2[4]) );
  DFFTRX1 R3_reg_4_ ( .D(R2[4]), .RN(n620), .CK(clk), .Q(R3[4]) );
  DFFTRX1 R4_reg_4_ ( .D(R3[4]), .RN(n619), .CK(clk), .Q(R4[4]) );
  DFFTRX1 R5_reg_4_ ( .D(R4[4]), .RN(n619), .CK(clk), .Q(R5[4]) );
  DFFTRX1 R7_reg_4_ ( .D(R6[4]), .RN(n619), .CK(clk), .Q(R7[4]) );
  DFFTRX1 R8_reg_4_ ( .D(R7[4]), .RN(n619), .CK(clk), .Q(R8[4]) );
  DFFTRX1 R9_reg_4_ ( .D(R8[4]), .RN(n619), .CK(clk), .Q(R9[4]) );
  DFFTRX1 R10_reg_4_ ( .D(R9[4]), .RN(n619), .CK(clk), .Q(R10[4]) );
  DFFTRX1 R11_reg_4_ ( .D(R10[4]), .RN(n619), .CK(clk), .Q(R11[4]) );
  DFFTRX1 R12_reg_4_ ( .D(R11[4]), .RN(n619), .CK(clk), .Q(R12[4]) );
  DFFTRX1 R13_reg_4_ ( .D(R12[4]), .RN(n619), .CK(clk), .Q(R13[4]) );
  DFFTRX1 R2_reg_3_ ( .D(R1[3]), .RN(n618), .CK(clk), .Q(R2[3]) );
  DFFTRX1 R3_reg_3_ ( .D(R2[3]), .RN(n618), .CK(clk), .Q(R3[3]) );
  DFFTRX1 R4_reg_3_ ( .D(R3[3]), .RN(n618), .CK(clk), .Q(R4[3]) );
  DFFTRX1 R5_reg_3_ ( .D(R4[3]), .RN(n618), .CK(clk), .Q(R5[3]) );
  DFFTRX1 R7_reg_3_ ( .D(R6[3]), .RN(n618), .CK(clk), .Q(R7[3]) );
  DFFTRX1 R8_reg_3_ ( .D(R7[3]), .RN(n618), .CK(clk), .Q(R8[3]) );
  DFFTRX1 R9_reg_3_ ( .D(R8[3]), .RN(n618), .CK(clk), .Q(R9[3]) );
  DFFTRX1 R10_reg_3_ ( .D(R9[3]), .RN(n618), .CK(clk), .Q(R10[3]) );
  DFFTRX1 R11_reg_3_ ( .D(R10[3]), .RN(n618), .CK(clk), .Q(R11[3]) );
  DFFTRX1 R12_reg_3_ ( .D(R11[3]), .RN(n618), .CK(clk), .Q(R12[3]) );
  DFFTRX1 R13_reg_3_ ( .D(R12[3]), .RN(n617), .CK(clk), .Q(R13[3]) );
  DFFTRX1 R2_reg_2_ ( .D(R1[2]), .RN(n617), .CK(clk), .Q(R2[2]) );
  DFFTRX1 R3_reg_2_ ( .D(R2[2]), .RN(n617), .CK(clk), .Q(R3[2]) );
  DFFTRX1 R4_reg_2_ ( .D(R3[2]), .RN(n617), .CK(clk), .Q(R4[2]) );
  DFFTRX1 R5_reg_2_ ( .D(R4[2]), .RN(n617), .CK(clk), .Q(R5[2]) );
  DFFTRX1 R7_reg_2_ ( .D(R6[2]), .RN(n617), .CK(clk), .Q(R7[2]) );
  DFFTRX1 R8_reg_2_ ( .D(R7[2]), .RN(n617), .CK(clk), .Q(R8[2]) );
  DFFTRX1 R9_reg_2_ ( .D(R8[2]), .RN(n617), .CK(clk), .Q(R9[2]) );
  DFFTRX1 R10_reg_2_ ( .D(R9[2]), .RN(n616), .CK(clk), .Q(R10[2]) );
  DFFTRX1 R11_reg_2_ ( .D(R10[2]), .RN(n616), .CK(clk), .Q(R11[2]) );
  DFFTRX1 R12_reg_2_ ( .D(R11[2]), .RN(n616), .CK(clk), .Q(R12[2]) );
  DFFTRX1 R13_reg_2_ ( .D(R12[2]), .RN(n616), .CK(clk), .Q(R13[2]) );
  DFFTRX1 R2_reg_1_ ( .D(R1[1]), .RN(n616), .CK(clk), .Q(R2[1]) );
  DFFTRX1 R3_reg_1_ ( .D(R2[1]), .RN(n616), .CK(clk), .Q(R3[1]) );
  DFFTRX1 R4_reg_1_ ( .D(R3[1]), .RN(n616), .CK(clk), .Q(R4[1]) );
  DFFTRX1 R5_reg_1_ ( .D(R4[1]), .RN(n616), .CK(clk), .Q(R5[1]) );
  DFFTRX1 R7_reg_1_ ( .D(R6[1]), .RN(n615), .CK(clk), .Q(R7[1]) );
  DFFTRX1 R8_reg_1_ ( .D(R7[1]), .RN(n615), .CK(clk), .Q(R8[1]) );
  DFFTRX1 R9_reg_1_ ( .D(R8[1]), .RN(n615), .CK(clk), .Q(R9[1]) );
  DFFTRX1 R10_reg_1_ ( .D(R9[1]), .RN(n615), .CK(clk), .Q(R10[1]) );
  DFFTRX1 R11_reg_1_ ( .D(R10[1]), .RN(n615), .CK(clk), .Q(R11[1]) );
  DFFTRX1 R12_reg_1_ ( .D(R11[1]), .RN(n615), .CK(clk), .Q(R12[1]) );
  DFFTRX1 R13_reg_1_ ( .D(R12[1]), .RN(n615), .CK(clk), .Q(R13[1]) );
  DFFTRX1 R2_reg_0_ ( .D(R1[0]), .RN(n615), .CK(clk), .Q(R2[0]) );
  DFFTRX1 R3_reg_0_ ( .D(R2[0]), .RN(n615), .CK(clk), .Q(R3[0]) );
  DFFTRX1 R4_reg_0_ ( .D(R3[0]), .RN(n614), .CK(clk), .Q(R4[0]) );
  DFFTRX1 R5_reg_0_ ( .D(R4[0]), .RN(n614), .CK(clk), .Q(R5[0]) );
  DFFTRX1 R7_reg_0_ ( .D(R6[0]), .RN(n614), .CK(clk), .Q(R7[0]) );
  DFFTRX1 R8_reg_0_ ( .D(R7[0]), .RN(n614), .CK(clk), .Q(R8[0]) );
  DFFTRX1 R9_reg_0_ ( .D(R8[0]), .RN(n614), .CK(clk), .Q(R9[0]) );
  DFFTRX1 R10_reg_0_ ( .D(R9[0]), .RN(n614), .CK(clk), .Q(R10[0]) );
  DFFTRX1 R11_reg_0_ ( .D(R10[0]), .RN(n614), .CK(clk), .Q(R11[0]) );
  DFFTRX1 R12_reg_0_ ( .D(R11[0]), .RN(n614), .CK(clk), .Q(R12[0]) );
  DFFTRX1 R13_reg_0_ ( .D(R12[0]), .RN(n614), .CK(clk), .Q(R13[0]) );
  DFFHQXL Wt_reg_20_ ( .D(N2151), .CK(clk), .Q(Wt[20]) );
  DFFHQXL Wt_reg_18_ ( .D(N2149), .CK(clk), .Q(Wt[18]) );
  DFFHQXL Wt_reg_15_ ( .D(N2146), .CK(clk), .Q(n2216) );
  DFFTRX2 R1_reg_30_ ( .D(Wt[30]), .RN(n652), .CK(clk), .Q(R1[30]) );
  DFFTRX2 R1_reg_31_ ( .D(Wt[31]), .RN(n653), .CK(clk), .Q(R1[31]) );
  DFFHQXL buffer_reg_0__24_ ( .D(n839), .CK(clk), .Q(buffer[120]) );
  DFFHQXL buffer_reg_0__25_ ( .D(n838), .CK(clk), .Q(buffer[121]) );
  DFFHQXL buffer_reg_0__26_ ( .D(n837), .CK(clk), .Q(buffer[122]) );
  DFFHQXL buffer_reg_0__27_ ( .D(n836), .CK(clk), .Q(buffer[123]) );
  DFFHQXL buffer_reg_0__28_ ( .D(n835), .CK(clk), .Q(buffer[124]) );
  DFFHQXL buffer_reg_0__29_ ( .D(n834), .CK(clk), .Q(buffer[125]) );
  DFFHQXL buffer_reg_0__30_ ( .D(n833), .CK(clk), .Q(buffer[126]) );
  DFFHQXL buffer_reg_0__31_ ( .D(n832), .CK(clk), .Q(buffer[127]) );
  DFFHQXL buffer_reg_2__24_ ( .D(n901), .CK(clk), .Q(buffer[104]) );
  DFFHQXL buffer_reg_2__25_ ( .D(n900), .CK(clk), .Q(buffer[105]) );
  DFFHQXL buffer_reg_2__26_ ( .D(n899), .CK(clk), .Q(buffer[106]) );
  DFFHQXL buffer_reg_2__27_ ( .D(n898), .CK(clk), .Q(buffer[107]) );
  DFFHQXL buffer_reg_2__28_ ( .D(n897), .CK(clk), .Q(buffer[108]) );
  DFFHQXL buffer_reg_2__29_ ( .D(n896), .CK(clk), .Q(buffer[109]) );
  DFFHQXL buffer_reg_2__30_ ( .D(n895), .CK(clk), .Q(buffer[110]) );
  DFFHQXL buffer_reg_2__31_ ( .D(n894), .CK(clk), .Q(buffer[111]) );
  DFFHQXL buffer_reg_3__24_ ( .D(n932), .CK(clk), .Q(buffer[96]) );
  DFFHQXL buffer_reg_3__25_ ( .D(n931), .CK(clk), .Q(buffer[97]) );
  DFFHQXL buffer_reg_3__26_ ( .D(n930), .CK(clk), .Q(buffer[98]) );
  DFFHQXL buffer_reg_3__27_ ( .D(n929), .CK(clk), .Q(buffer[99]) );
  DFFHQXL buffer_reg_3__28_ ( .D(n928), .CK(clk), .Q(buffer[100]) );
  DFFHQXL buffer_reg_3__29_ ( .D(n927), .CK(clk), .Q(buffer[101]) );
  DFFHQXL buffer_reg_3__30_ ( .D(n926), .CK(clk), .Q(buffer[102]) );
  DFFHQXL buffer_reg_3__31_ ( .D(n925), .CK(clk), .Q(buffer[103]) );
  DFFHQXL buffer_reg_1__24_ ( .D(n870), .CK(clk), .Q(buffer[112]) );
  DFFHQXL buffer_reg_1__25_ ( .D(n869), .CK(clk), .Q(buffer[113]) );
  DFFHQXL buffer_reg_1__26_ ( .D(n868), .CK(clk), .Q(buffer[114]) );
  DFFHQXL buffer_reg_1__27_ ( .D(n867), .CK(clk), .Q(buffer[115]) );
  DFFHQXL buffer_reg_1__28_ ( .D(n866), .CK(clk), .Q(buffer[116]) );
  DFFHQXL buffer_reg_1__29_ ( .D(n865), .CK(clk), .Q(buffer[117]) );
  DFFHQXL buffer_reg_1__30_ ( .D(n864), .CK(clk), .Q(buffer[118]) );
  DFFHQXL buffer_reg_1__31_ ( .D(n863), .CK(clk), .Q(buffer[119]) );
  DFFHQXL buffer_reg_0__0_ ( .D(n2210), .CK(clk), .Q(N442) );
  DFFHQXL buffer_reg_0__1_ ( .D(n831), .CK(clk), .Q(N443) );
  DFFHQXL buffer_reg_0__2_ ( .D(n830), .CK(clk), .Q(N444) );
  DFFHQXL buffer_reg_0__3_ ( .D(n829), .CK(clk), .Q(N445) );
  DFFHQXL buffer_reg_0__4_ ( .D(n828), .CK(clk), .Q(N446) );
  DFFHQXL buffer_reg_0__5_ ( .D(n827), .CK(clk), .Q(N447) );
  DFFHQXL buffer_reg_0__6_ ( .D(n826), .CK(clk), .Q(N448) );
  DFFHQXL buffer_reg_0__7_ ( .D(n825), .CK(clk), .Q(N449) );
  DFFHQXL buffer_reg_2__0_ ( .D(n2212), .CK(clk), .Q(N506) );
  DFFHQXL buffer_reg_2__1_ ( .D(n893), .CK(clk), .Q(N507) );
  DFFHQXL buffer_reg_2__2_ ( .D(n892), .CK(clk), .Q(N508) );
  DFFHQXL buffer_reg_2__3_ ( .D(n891), .CK(clk), .Q(N509) );
  DFFHQXL buffer_reg_2__4_ ( .D(n890), .CK(clk), .Q(N510) );
  DFFHQXL buffer_reg_2__5_ ( .D(n889), .CK(clk), .Q(N511) );
  DFFHQXL buffer_reg_2__6_ ( .D(n888), .CK(clk), .Q(N512) );
  DFFHQXL buffer_reg_2__7_ ( .D(n887), .CK(clk), .Q(N513) );
  DFFHQXL buffer_reg_3__0_ ( .D(n2211), .CK(clk), .Q(N538) );
  DFFHQXL buffer_reg_3__1_ ( .D(n924), .CK(clk), .Q(N539) );
  DFFHQXL buffer_reg_3__2_ ( .D(n923), .CK(clk), .Q(N540) );
  DFFHQXL buffer_reg_3__3_ ( .D(n922), .CK(clk), .Q(N541) );
  DFFHQXL buffer_reg_3__4_ ( .D(n921), .CK(clk), .Q(N542) );
  DFFHQXL buffer_reg_3__5_ ( .D(n920), .CK(clk), .Q(N543) );
  DFFHQXL buffer_reg_3__6_ ( .D(n919), .CK(clk), .Q(N544) );
  DFFHQXL buffer_reg_3__7_ ( .D(n918), .CK(clk), .Q(N545) );
  DFFHQXL buffer_reg_1__0_ ( .D(n2197), .CK(clk), .Q(N474) );
  DFFHQXL buffer_reg_1__1_ ( .D(n862), .CK(clk), .Q(N475) );
  DFFHQXL buffer_reg_1__2_ ( .D(n861), .CK(clk), .Q(N476) );
  DFFHQXL buffer_reg_1__3_ ( .D(n860), .CK(clk), .Q(N477) );
  DFFHQXL buffer_reg_1__4_ ( .D(n859), .CK(clk), .Q(N478) );
  DFFHQXL buffer_reg_1__5_ ( .D(n858), .CK(clk), .Q(N479) );
  DFFHQXL buffer_reg_1__6_ ( .D(n857), .CK(clk), .Q(N480) );
  DFFHQXL buffer_reg_1__7_ ( .D(n856), .CK(clk), .Q(N481) );
  DFFHQXL buffer_reg_0__8_ ( .D(n855), .CK(clk), .Q(N450) );
  DFFHQXL buffer_reg_0__9_ ( .D(n854), .CK(clk), .Q(N451) );
  DFFHQXL buffer_reg_0__10_ ( .D(n853), .CK(clk), .Q(N452) );
  DFFHQXL buffer_reg_0__11_ ( .D(n852), .CK(clk), .Q(N453) );
  DFFHQXL buffer_reg_0__12_ ( .D(n851), .CK(clk), .Q(N454) );
  DFFHQXL buffer_reg_0__13_ ( .D(n850), .CK(clk), .Q(N455) );
  DFFHQXL buffer_reg_0__14_ ( .D(n849), .CK(clk), .Q(N456) );
  DFFHQXL buffer_reg_0__15_ ( .D(n848), .CK(clk), .Q(N457) );
  DFFHQXL buffer_reg_0__16_ ( .D(n847), .CK(clk), .Q(N458) );
  DFFHQXL buffer_reg_0__17_ ( .D(n846), .CK(clk), .Q(N459) );
  DFFHQXL buffer_reg_0__18_ ( .D(n845), .CK(clk), .Q(N460) );
  DFFHQXL buffer_reg_0__19_ ( .D(n844), .CK(clk), .Q(N461) );
  DFFHQXL buffer_reg_0__20_ ( .D(n843), .CK(clk), .Q(N462) );
  DFFHQXL buffer_reg_0__21_ ( .D(n842), .CK(clk), .Q(N463) );
  DFFHQXL buffer_reg_0__22_ ( .D(n841), .CK(clk), .Q(N464) );
  DFFHQXL buffer_reg_0__23_ ( .D(n840), .CK(clk), .Q(N465) );
  DFFHQXL buffer_reg_2__8_ ( .D(n917), .CK(clk), .Q(N514) );
  DFFHQXL buffer_reg_2__9_ ( .D(n916), .CK(clk), .Q(N515) );
  DFFHQXL buffer_reg_2__10_ ( .D(n915), .CK(clk), .Q(N516) );
  DFFHQXL buffer_reg_2__11_ ( .D(n914), .CK(clk), .Q(N517) );
  DFFHQXL buffer_reg_2__12_ ( .D(n913), .CK(clk), .Q(N518) );
  DFFHQXL buffer_reg_2__13_ ( .D(n912), .CK(clk), .Q(N519) );
  DFFHQXL buffer_reg_2__14_ ( .D(n911), .CK(clk), .Q(N520) );
  DFFHQXL buffer_reg_2__15_ ( .D(n910), .CK(clk), .Q(N521) );
  DFFHQXL buffer_reg_2__16_ ( .D(n909), .CK(clk), .Q(N522) );
  DFFHQXL buffer_reg_2__17_ ( .D(n908), .CK(clk), .Q(N523) );
  DFFHQXL buffer_reg_2__18_ ( .D(n907), .CK(clk), .Q(N524) );
  DFFHQXL buffer_reg_2__19_ ( .D(n906), .CK(clk), .Q(N525) );
  DFFHQXL buffer_reg_2__20_ ( .D(n905), .CK(clk), .Q(N526) );
  DFFHQXL buffer_reg_2__21_ ( .D(n904), .CK(clk), .Q(N527) );
  DFFHQXL buffer_reg_2__22_ ( .D(n903), .CK(clk), .Q(N528) );
  DFFHQXL buffer_reg_2__23_ ( .D(n902), .CK(clk), .Q(N529) );
  DFFHQXL buffer_reg_3__8_ ( .D(n948), .CK(clk), .Q(N546) );
  DFFHQXL buffer_reg_3__9_ ( .D(n947), .CK(clk), .Q(N547) );
  DFFHQXL buffer_reg_3__10_ ( .D(n946), .CK(clk), .Q(N548) );
  DFFHQXL buffer_reg_3__11_ ( .D(n945), .CK(clk), .Q(N549) );
  DFFHQXL buffer_reg_3__12_ ( .D(n944), .CK(clk), .Q(N550) );
  DFFHQXL buffer_reg_3__13_ ( .D(n943), .CK(clk), .Q(N551) );
  DFFHQXL buffer_reg_3__14_ ( .D(n942), .CK(clk), .Q(N552) );
  DFFHQXL buffer_reg_3__15_ ( .D(n941), .CK(clk), .Q(N553) );
  DFFHQXL buffer_reg_3__16_ ( .D(n940), .CK(clk), .Q(N554) );
  DFFHQXL buffer_reg_3__17_ ( .D(n939), .CK(clk), .Q(N555) );
  DFFHQXL buffer_reg_3__18_ ( .D(n938), .CK(clk), .Q(N556) );
  DFFHQXL buffer_reg_3__19_ ( .D(n937), .CK(clk), .Q(N557) );
  DFFHQXL buffer_reg_3__20_ ( .D(n936), .CK(clk), .Q(N558) );
  DFFHQXL buffer_reg_3__21_ ( .D(n935), .CK(clk), .Q(N559) );
  DFFHQXL buffer_reg_3__22_ ( .D(n934), .CK(clk), .Q(N560) );
  DFFHQXL buffer_reg_3__23_ ( .D(n933), .CK(clk), .Q(N561) );
  DFFHQXL buffer_reg_1__8_ ( .D(n886), .CK(clk), .Q(N482) );
  DFFHQXL buffer_reg_1__9_ ( .D(n885), .CK(clk), .Q(N483) );
  DFFHQXL buffer_reg_1__10_ ( .D(n884), .CK(clk), .Q(N484) );
  DFFHQXL buffer_reg_1__11_ ( .D(n883), .CK(clk), .Q(N485) );
  DFFHQXL buffer_reg_1__12_ ( .D(n882), .CK(clk), .Q(N486) );
  DFFHQXL buffer_reg_1__13_ ( .D(n881), .CK(clk), .Q(N487) );
  DFFHQXL buffer_reg_1__14_ ( .D(n880), .CK(clk), .Q(N488) );
  DFFHQXL buffer_reg_1__15_ ( .D(n879), .CK(clk), .Q(N489) );
  DFFHQXL buffer_reg_1__16_ ( .D(n878), .CK(clk), .Q(N490) );
  DFFHQXL buffer_reg_1__17_ ( .D(n877), .CK(clk), .Q(N491) );
  DFFHQXL buffer_reg_1__18_ ( .D(n876), .CK(clk), .Q(N492) );
  DFFHQXL buffer_reg_1__19_ ( .D(n875), .CK(clk), .Q(N493) );
  DFFHQXL buffer_reg_1__20_ ( .D(n874), .CK(clk), .Q(N494) );
  DFFHQXL buffer_reg_1__21_ ( .D(n873), .CK(clk), .Q(N495) );
  DFFHQXL buffer_reg_1__22_ ( .D(n872), .CK(clk), .Q(N496) );
  DFFHQXL buffer_reg_1__23_ ( .D(n871), .CK(clk), .Q(N497) );
  DFFHQXL Wt_reg_29_ ( .D(N2160), .CK(clk), .Q(Wt[29]) );
  DFFHQXL Wt_reg_28_ ( .D(N2159), .CK(clk), .Q(Wt[28]) );
  DFFHQXL Wt_reg_27_ ( .D(N2158), .CK(clk), .Q(Wt[27]) );
  DFFHQXL Wt_reg_24_ ( .D(N2155), .CK(clk), .Q(Wt[24]) );
  DFFHQXL Wt_reg_26_ ( .D(N2157), .CK(clk), .Q(Wt[26]) );
  DFFHQXL Wt_reg_25_ ( .D(N2156), .CK(clk), .Q(Wt[25]) );
  DFFHQXL Wt_reg_22_ ( .D(N2153), .CK(clk), .Q(Wt[22]) );
  DFFHQXL Wt_reg_23_ ( .D(N2154), .CK(clk), .Q(Wt[23]) );
  DFFHQXL Wt_reg_21_ ( .D(N2152), .CK(clk), .Q(Wt[21]) );
  DFFTRX2 R1_reg_23_ ( .D(Wt[23]), .RN(n643), .CK(clk), .Q(R1[23]) );
  DFFTRX4 R14_reg_18_ ( .D(R13[18]), .RN(n636), .CK(clk), .Q(R14[18]) );
  DFFTRX4 R1_reg_17_ ( .D(Wt[17]), .RN(n636), .CK(clk), .Q(R1[17]) );
  DFFTRX4 R14_reg_7_ ( .D(R13[7]), .RN(n622), .CK(clk), .Q(R14[7]) );
  DFFHQXL Wt_reg_31_ ( .D(N2162), .CK(clk), .Q(Wt[31]) );
  DFFTRX4 R1_reg_19_ ( .D(Wt[19]), .RN(n638), .CK(clk), .Q(R1[19]) );
  DFFHQX1 Wt_reg_9_ ( .D(N2140), .CK(clk), .Q(Wt[9]) );
  DFFHQX2 Wt_reg_2_ ( .D(N2133), .CK(clk), .Q(Wt[2]) );
  DFFTRX2 R14_reg_9_ ( .D(R13[9]), .RN(n625), .CK(clk), .Q(R14[9]) );
  DFFTRX4 R6_reg_1_ ( .D(R5[1]), .RN(n616), .CK(clk), .Q(R6[1]) );
  DFFTRX2 R1_reg_27_ ( .D(Wt[27]), .RN(n648), .CK(clk), .Q(R1[27]) );
  DFFTRX2 R1_reg_26_ ( .D(Wt[26]), .RN(n647), .CK(clk), .Q(R1[26]) );
  DFFTRX2 R14_reg_26_ ( .D(R13[26]), .RN(n646), .CK(clk), .Q(R14[26]) );
  DFFTRX2 R14_reg_27_ ( .D(R13[27]), .RN(n647), .CK(clk), .Q(R14[27]) );
  DFFTRX2 R14_reg_31_ ( .D(R13[31]), .RN(n652), .CK(clk), .Q(R14[31]) );
  DFFTRX2 R1_reg_28_ ( .D(Wt[28]), .RN(n650), .CK(clk), .Q(R1[28]) );
  DFFTRX2 R1_reg_29_ ( .D(Wt[29]), .RN(n651), .CK(clk), .Q(R1[29]) );
  DFFTRX2 R14_reg_16_ ( .D(R13[16]), .RN(n634), .CK(clk), .Q(R14[16]) );
  DFFTRX2 R14_reg_15_ ( .D(R13[15]), .RN(n632), .CK(clk), .Q(R14[15]) );
  DFFTRX2 R14_reg_23_ ( .D(R13[23]), .RN(n642), .CK(clk), .Q(R14[23]) );
  DFFTRX2 R6_reg_6_ ( .D(R5[6]), .RN(n622), .CK(clk), .Q(R6[6]) );
  DFFTRX2 R14_reg_10_ ( .D(R13[10]), .RN(n626), .CK(clk), .Q(R14[10]) );
  DFFTRX2 R1_reg_18_ ( .D(Wt[18]), .RN(n637), .CK(clk), .Q(R1[18]) );
  DFFTRX2 R14_reg_5_ ( .D(R13[5]), .RN(n620), .CK(clk), .Q(R14[5]) );
  DFFTRX2 R14_reg_4_ ( .D(R13[4]), .RN(n619), .CK(clk), .Q(R14[4]) );
  DFFTRX4 R14_reg_19_ ( .D(R13[19]), .RN(n637), .CK(clk), .Q(R14[19]) );
  DFFHQX2 Wt_reg_13_ ( .D(N2144), .CK(clk), .Q(Wt[13]) );
  DFFTRX4 R15_reg_1_ ( .D(R14[1]), .RN(n615), .CK(clk), .Q(R15[1]) );
  DFFTRX2 R6_reg_0_ ( .D(R5[0]), .RN(n614), .CK(clk), .Q(R6[0]) );
  DFFHQX2 Wt_reg_6_ ( .D(N2137), .CK(clk), .Q(Wt[6]) );
  DFFHQX2 Wt_reg_10_ ( .D(N2141), .CK(clk), .Q(Wt[10]) );
  DFFTRX2 R1_reg_10_ ( .D(Wt[10]), .RN(n627), .CK(clk), .Q(R1[10]) );
  DFFTRX2 R15_reg_0_ ( .D(R14[0]), .RN(n614), .CK(clk), .Q(R15[0]) );
  DFFTRX4 R1_reg_20_ ( .D(Wt[20]), .RN(n640), .CK(clk), .Q(R1[20]) );
  DFFXL buffer_reg_11__19_ ( .D(n1912), .CK(clk), .Q(N813) );
  DFFHQXL buffer_reg_5__28_ ( .D(n990), .CK(clk), .Q(buffer[84]) );
  DFFTRX2 R14_reg_30_ ( .D(R13[30]), .RN(n651), .CK(clk), .Q(R14[30]) );
  DFFTRX2 R14_reg_3_ ( .D(R13[3]), .RN(n617), .CK(clk), .Q(R14[3]) );
  DFFTRX2 R14_reg_12_ ( .D(R13[12]), .RN(n629), .CK(clk), .Q(R14[12]) );
  DFFTRX2 R14_reg_11_ ( .D(R13[11]), .RN(n627), .CK(clk), .Q(R14[11]) );
  DFFTRX2 R14_reg_13_ ( .D(R13[13]), .RN(n630), .CK(clk), .Q(R14[13]) );
  DFFTRX2 R14_reg_29_ ( .D(R13[29]), .RN(n650), .CK(clk), .Q(R14[29]) );
  DFFHQX1 Wt_reg_19_ ( .D(N2150), .CK(clk), .Q(Wt[19]) );
  DFFTRX1 R15_reg_9_ ( .D(R14[9]), .RN(n625), .CK(clk), .Q(R15[9]) );
  DFFTRX2 R1_reg_25_ ( .D(Wt[25]), .RN(n646), .CK(clk), .Q(R1[25]) );
  DFFTRX2 R1_reg_24_ ( .D(Wt[24]), .RN(n645), .CK(clk), .Q(R1[24]) );
  DFFTRX1 R15_reg_16_ ( .D(R14[16]), .RN(n634), .CK(clk), .Q(R15[16]) );
  DFFTRX2 R14_reg_17_ ( .D(R13[17]), .RN(n635), .CK(clk), .Q(R14[17]) );
  DFFTRX1 R15_reg_17_ ( .D(R14[17]), .RN(n635), .CK(clk), .Q(R15[17]) );
  DFFTRX2 R14_reg_22_ ( .D(R13[22]), .RN(n641), .CK(clk), .Q(R14[22]) );
  DFFTRX1 R15_reg_15_ ( .D(R14[15]), .RN(n632), .CK(clk), .Q(R15[15]) );
  DFFTRX2 R14_reg_14_ ( .D(R13[14]), .RN(n631), .CK(clk), .Q(R14[14]) );
  DFFTRX1 R15_reg_14_ ( .D(R14[14]), .RN(n631), .CK(clk), .Q(R15[14]) );
  DFFTRX1 R15_reg_8_ ( .D(R14[8]), .RN(n624), .CK(clk), .Q(R15[8]) );
  DFFTRX1 R15_reg_10_ ( .D(R14[10]), .RN(n626), .CK(clk), .Q(R15[10]) );
  DFFTRX1 R15_reg_5_ ( .D(R14[5]), .RN(n620), .CK(clk), .Q(R15[5]) );
  DFFTRX2 R14_reg_25_ ( .D(R13[25]), .RN(n645), .CK(clk), .Q(R14[25]) );
  DFFTRX2 R15_reg_4_ ( .D(R14[4]), .RN(n619), .CK(clk), .Q(R15[4]) );
  DFFHQX1 Wt_reg_16_ ( .D(N2147), .CK(clk), .Q(Wt[16]) );
  DFFHQX2 Wt_reg_12_ ( .D(N2143), .CK(clk), .Q(Wt[12]) );
  DFFTRX2 R1_reg_12_ ( .D(Wt[12]), .RN(n630), .CK(clk), .Q(R1[12]) );
  DFFTRX1 R6_reg_13_ ( .D(R5[13]), .RN(n631), .CK(clk), .Q(R6[13]) );
  DFFTRX1 R1_reg_15_ ( .D(Wt[15]), .RN(n633), .CK(clk), .Q(R1[15]) );
  DFFTRX1 R6_reg_8_ ( .D(R5[8]), .RN(n624), .CK(clk), .Q(R6[8]) );
  DFFTRX1 R6_reg_9_ ( .D(R5[9]), .RN(n626), .CK(clk), .Q(R6[9]) );
  DFFTRX1 R14_reg_1_ ( .D(R13[1]), .RN(n615), .CK(clk), .Q(R14[1]) );
  DFFX2 Wt_reg_14_ ( .D(N2145), .CK(clk), .Q(Wt[14]) );
  DFFTRX2 R6_reg_4_ ( .D(R5[4]), .RN(n619), .CK(clk), .Q(R6[4]) );
  DFFTRX1 R6_reg_7_ ( .D(R5[7]), .RN(n623), .CK(clk), .Q(R6[7]) );
  DFFTRX1 R6_reg_3_ ( .D(R5[3]), .RN(n618), .CK(clk), .Q(R6[3]) );
  DFFTRX1 R6_reg_2_ ( .D(R5[2]), .RN(n617), .CK(clk), .Q(R6[2]) );
  DFFTRX2 R1_reg_22_ ( .D(Wt[22]), .RN(n642), .CK(clk), .Q(R1[22]) );
  DFFTRX2 R14_reg_8_ ( .D(R13[8]), .RN(n624), .CK(clk), .Q(R14[8]) );
  DFFHQX2 Wt_reg_3_ ( .D(N2134), .CK(clk), .Q(Wt[3]) );
  DFFHQX2 Wt_reg_4_ ( .D(N2135), .CK(clk), .Q(Wt[4]) );
  DFFHQX2 Wt_reg_5_ ( .D(N2136), .CK(clk), .Q(Wt[5]) );
  DFFHQX2 Wt_reg_0_ ( .D(N2131), .CK(clk), .Q(Wt[0]) );
  DFFTRX2 R1_reg_0_ ( .D(Wt[0]), .RN(n615), .CK(clk), .Q(R1[0]) );
  DFFHQX4 Wt_reg_7_ ( .D(N2138), .CK(clk), .Q(Wt[7]) );
  DFFTRX2 R14_reg_6_ ( .D(R13[6]), .RN(n621), .CK(clk), .Q(R14[6]) );
  DFFTRX4 R15_reg_6_ ( .D(R14[6]), .RN(n621), .CK(clk), .Q(R15[6]) );
  DFFTRX2 R1_reg_13_ ( .D(Wt[13]), .RN(n631), .CK(clk), .Q(R1[13]) );
  DFFTRX4 R14_reg_28_ ( .D(R13[28]), .RN(n649), .CK(clk), .Q(R14[28]) );
  DFFTRX2 R1_reg_2_ ( .D(Wt[2]), .RN(n617), .CK(clk), .Q(R1[2]) );
  DFFTRX2 R1_reg_16_ ( .D(Wt[16]), .RN(n635), .CK(clk), .Q(R1[16]) );
  DFFTRX4 R14_reg_24_ ( .D(R13[24]), .RN(n644), .CK(clk), .Q(R14[24]) );
  DFFTRX2 R1_reg_11_ ( .D(Wt[11]), .RN(n628), .CK(clk), .Q(R1[11]) );
  DFFTRX4 R14_reg_20_ ( .D(R13[20]), .RN(n639), .CK(clk), .Q(R14[20]) );
  DFFHQX4 Wt_reg_1_ ( .D(N2132), .CK(clk), .Q(Wt[1]) );
  DFFTRX1 R1_reg_1_ ( .D(Wt[1]), .RN(n616), .CK(clk), .Q(R1[1]) );
  DFFTRX2 R6_reg_5_ ( .D(R5[5]), .RN(n621), .CK(clk), .Q(R6[5]) );
  DFFTRX4 R14_reg_21_ ( .D(R13[21]), .RN(n640), .CK(clk), .Q(R14[21]) );
  DFFTRX4 R1_reg_21_ ( .D(Wt[21]), .RN(n641), .CK(clk), .Q(R1[21]) );
  OR2X4 U3 ( .A(n1477), .B(reset), .Y(n56) );
  INVX16 U4 ( .A(n713), .Y(n711) );
  INVX4 U5 ( .A(n1621), .Y(n153) );
  INVX8 U6 ( .A(n59), .Y(n1225) );
  NOR2X4 U7 ( .A(n1657), .B(reset), .Y(n77) );
  INVX8 U8 ( .A(n737), .Y(n736) );
  INVX4 U9 ( .A(n738), .Y(n735) );
  NOR2X4 U10 ( .A(n741), .B(reset), .Y(n1116) );
  INVX8 U11 ( .A(n110), .Y(n113) );
  INVX4 U12 ( .A(n49), .Y(n727) );
  XOR2X1 U13 ( .A(R1[14]), .B(R1[16]), .Y(sigma1[29]) );
  XOR3X4 U14 ( .A(R1[23]), .B(R1[25]), .C(R1[16]), .Y(sigma1[6]) );
  INVX8 U15 ( .A(n706), .Y(n703) );
  INVX8 U16 ( .A(n705), .Y(n704) );
  NOR2X4 U17 ( .A(n708), .B(reset), .Y(n1373) );
  XOR3X4 U18 ( .A(R1[25]), .B(R1[2]), .C(R1[0]), .Y(sigma1[15]) );
  XOR3X2 U19 ( .A(R14[28]), .B(R14[17]), .C(R14[13]), .Y(sigma0[10]) );
  INVX12 U20 ( .A(n713), .Y(n712) );
  CLKINVX4 U21 ( .A(n1337), .Y(n713) );
  INVX4 U22 ( .A(n1658), .Y(n105) );
  XOR3X4 U23 ( .A(R1[20]), .B(R1[22]), .C(R1[13]), .Y(sigma1[3]) );
  XOR2XL U24 ( .A(R1[13]), .B(R1[15]), .Y(sigma1[28]) );
  XOR3X4 U25 ( .A(R14[21]), .B(R14[10]), .C(R14[6]), .Y(sigma0[3]) );
  NOR2X2 U26 ( .A(n146), .B(reset), .Y(n1514) );
  INVX8 U27 ( .A(n153), .Y(n154) );
  XOR3X2 U28 ( .A(R1[27]), .B(R1[29]), .C(R1[20]), .Y(sigma1[10]) );
  INVXL U29 ( .A(n1191), .Y(n730) );
  CLKINVX3 U30 ( .A(n1444), .Y(n692) );
  CLKINVX3 U31 ( .A(n1409), .Y(n698) );
  AOI2BB1X2 U32 ( .A0N(n1510), .A1N(n1511), .B0(reset), .Y(n1477) );
  INVX1 U33 ( .A(data[3]), .Y(n119) );
  INVX4 U34 ( .A(n110), .Y(n112) );
  BUFX4 U35 ( .A(n77), .Y(n175) );
  CLKINVX3 U36 ( .A(n702), .Y(n699) );
  CLKINVX3 U37 ( .A(n72), .Y(n681) );
  INVX1 U38 ( .A(N807), .Y(n114) );
  AOI22X1 U39 ( .A0(n142), .A1(N811), .B0(N803), .B1(n113), .Y(n1528) );
  INVX1 U40 ( .A(n1630), .Y(n2160) );
  INVX1 U41 ( .A(n1637), .Y(n2167) );
  XOR3X2 U42 ( .A(R14[19]), .B(R14[30]), .C(R14[15]), .Y(sigma0[12]) );
  XOR3X2 U43 ( .A(R14[27]), .B(R14[16]), .C(R14[12]), .Y(sigma0[9]) );
  NOR2X2 U44 ( .A(n716), .B(reset), .Y(n1337) );
  CLKINVX3 U45 ( .A(n1373), .Y(n705) );
  NOR2X2 U46 ( .A(n721), .B(reset), .Y(n1266) );
  INVX8 U47 ( .A(n734), .Y(n733) );
  INVX8 U48 ( .A(n56), .Y(n172) );
  CLKINVX3 U49 ( .A(n135), .Y(Wt[15]) );
  INVX1 U50 ( .A(n2216), .Y(n135) );
  NAND2X1 U51 ( .A(logic_result[23]), .B(n605), .Y(n790) );
  NAND2X1 U52 ( .A(n815), .B(n814), .Y(N2160) );
  NAND2X1 U53 ( .A(logic_result[29]), .B(n606), .Y(n814) );
  AOI22X1 U54 ( .A0(n733), .A1(N485), .B0(N477), .B1(n731), .Y(n1179) );
  AOI22X1 U55 ( .A0(n729), .A1(N517), .B0(N509), .B1(n727), .Y(n1212) );
  AOI22X1 U56 ( .A0(n740), .A1(N453), .B0(N445), .B1(n735), .Y(n1136) );
  AOI22X1 U57 ( .A0(n733), .A1(buffer[112]), .B0(N490), .B1(n732), .Y(n1166)
         );
  AOI22X1 U58 ( .A0(n728), .A1(buffer[104]), .B0(N522), .B1(n727), .Y(n1199)
         );
  AOI22X1 U59 ( .A0(n739), .A1(buffer[120]), .B0(N458), .B1(n736), .Y(n1123)
         );
  INVX1 U60 ( .A(N732), .Y(n101) );
  INVX1 U61 ( .A(N731), .Y(n109) );
  INVX1 U62 ( .A(n1475), .Y(n2204) );
  AOI22X1 U63 ( .A0(n142), .A1(N806), .B0(N798), .B1(n112), .Y(n1533) );
  INVX1 U64 ( .A(N803), .Y(n74) );
  INVX1 U65 ( .A(n1538), .Y(n1804) );
  INVX1 U66 ( .A(data[4]), .Y(n66) );
  INVX1 U67 ( .A(n112), .Y(n67) );
  INVX1 U68 ( .A(N797), .Y(n64) );
  AOI22X2 U69 ( .A0(n677), .A1(N943), .B0(N935), .B1(n174), .Y(n1668) );
  OAI2BB2X1 U70 ( .B0(n95), .B1(n105), .A0N(n677), .A1N(N942), .Y(n94) );
  INVX1 U71 ( .A(N934), .Y(n95) );
  OAI2BB2X1 U72 ( .B0(n97), .B1(n105), .A0N(n677), .A1N(N939), .Y(n96) );
  INVX1 U73 ( .A(N931), .Y(n97) );
  INVX1 U74 ( .A(N938), .Y(n82) );
  INVX1 U75 ( .A(n1675), .Y(n2190) );
  INVX1 U76 ( .A(n1676), .Y(n2191) );
  INVX1 U77 ( .A(n1677), .Y(n2192) );
  INVX1 U78 ( .A(n1678), .Y(n2193) );
  INVX1 U79 ( .A(n1679), .Y(n2194) );
  INVX1 U80 ( .A(n1680), .Y(n2195) );
  OAI2BB2X1 U81 ( .B0(n91), .B1(n105), .A0N(n678), .A1N(N930), .Y(n90) );
  INVX1 U82 ( .A(N922), .Y(n91) );
  INVX1 U83 ( .A(N929), .Y(n124) );
  INVX1 U84 ( .A(data[7]), .Y(n125) );
  INVX1 U85 ( .A(n1684), .Y(n2176) );
  INVX1 U86 ( .A(n1687), .Y(n2178) );
  INVX1 U87 ( .A(N706), .Y(n85) );
  INVX1 U88 ( .A(n1433), .Y(n1082) );
  INVX1 U89 ( .A(N704), .Y(n61) );
  INVX1 U90 ( .A(N703), .Y(n63) );
  INVX1 U91 ( .A(N702), .Y(n70) );
  INVX1 U92 ( .A(N701), .Y(n79) );
  INVX1 U93 ( .A(n697), .Y(n80) );
  INVX1 U94 ( .A(N700), .Y(n99) );
  INVX1 U95 ( .A(N699), .Y(n107) );
  INVX1 U96 ( .A(n1440), .Y(n2205) );
  INVX1 U97 ( .A(n1632), .Y(n2162) );
  INVX1 U98 ( .A(n1636), .Y(n2166) );
  INVX1 U99 ( .A(N896), .Y(n132) );
  AOI22X1 U100 ( .A0(n154), .A1(N903), .B0(N895), .B1(n72), .Y(n1640) );
  INVX1 U101 ( .A(N894), .Y(n130) );
  INVX1 U102 ( .A(N898), .Y(n133) );
  INVX1 U103 ( .A(n1646), .Y(n2148) );
  AOI22X1 U104 ( .A0(n154), .A1(N896), .B0(data[6]), .B1(n72), .Y(n1647) );
  AOI22X1 U105 ( .A0(n154), .A1(N895), .B0(data[5]), .B1(n72), .Y(n1648) );
  INVX1 U106 ( .A(n1650), .Y(n2152) );
  AOI22X1 U107 ( .A0(n693), .A1(buffer[48]), .B0(N746), .B1(n691), .Y(n1451)
         );
  AOI22X1 U108 ( .A0(n144), .A1(buffer[37]), .B0(N815), .B1(n111), .Y(n1516)
         );
  AOI22X1 U109 ( .A0(n144), .A1(buffer[33]), .B0(N811), .B1(n111), .Y(n1520)
         );
  OAI22X1 U110 ( .A0(n71), .A1(n103), .B0(n104), .B1(n105), .Y(n102) );
  INVX1 U111 ( .A(buffer[7]), .Y(n103) );
  INVX1 U112 ( .A(N945), .Y(n104) );
  OAI2BB2X1 U113 ( .B0(n87), .B1(n105), .A0N(n677), .A1N(buffer[5]), .Y(n86)
         );
  INVX1 U114 ( .A(N943), .Y(n87) );
  OAI2BB2X1 U115 ( .B0(n89), .B1(n105), .A0N(n678), .A1N(buffer[4]), .Y(n88)
         );
  INVX1 U116 ( .A(N942), .Y(n89) );
  INVX1 U117 ( .A(N941), .Y(n126) );
  OAI2BB2X1 U118 ( .B0(n93), .B1(n105), .A0N(n677), .A1N(buffer[2]), .Y(n92)
         );
  INVX1 U119 ( .A(N940), .Y(n93) );
  AOI22X1 U120 ( .A0(n699), .A1(buffer[56]), .B0(N714), .B1(n697), .Y(n1416)
         );
  INVX1 U121 ( .A(n1620), .Y(n2155) );
  INVX1 U122 ( .A(N910), .Y(n117) );
  INVX1 U123 ( .A(buffer[11]), .Y(n128) );
  INVX1 U124 ( .A(N909), .Y(n129) );
  INVX1 U125 ( .A(N908), .Y(n121) );
  INVX1 U126 ( .A(n1628), .Y(n2158) );
  AOI22X1 U127 ( .A0(n154), .A1(buffer[9]), .B0(N907), .B1(n75), .Y(n1628) );
  AOI22X1 U128 ( .A0(n154), .A1(buffer[8]), .B0(N906), .B1(n72), .Y(n1629) );
  AOI31X4 U129 ( .A0(n1224), .A1(n1225), .A2(n190), .B0(reset), .Y(n1191) );
  AOI22X1 U130 ( .A0(n677), .A1(buffer[1]), .B0(N939), .B1(n1658), .Y(n1664)
         );
  AOI22X1 U131 ( .A0(n678), .A1(N941), .B0(N933), .B1(n1658), .Y(n1670) );
  AOI22X1 U132 ( .A0(n677), .A1(N935), .B0(N927), .B1(n1658), .Y(n1676) );
  INVX2 U133 ( .A(n700), .Y(n84) );
  XOR3X2 U134 ( .A(R1[29]), .B(R1[31]), .C(R1[22]), .Y(sigma1[12]) );
  INVX8 U135 ( .A(n722), .Y(n721) );
  INVX4 U136 ( .A(n1265), .Y(n722) );
  AOI22X1 U137 ( .A0(n721), .A1(N577), .B0(data[7]), .B1(n138), .Y(n1290) );
  AOI22X1 U138 ( .A0(n721), .A1(N575), .B0(data[5]), .B1(n140), .Y(n1292) );
  AOI22X1 U139 ( .A0(n721), .A1(N574), .B0(data[4]), .B1(n140), .Y(n1293) );
  AOI22X1 U140 ( .A0(n721), .A1(N573), .B0(data[3]), .B1(n140), .Y(n1294) );
  AOI22X1 U141 ( .A0(n721), .A1(N572), .B0(data[2]), .B1(n138), .Y(n1295) );
  AOI22X1 U142 ( .A0(n721), .A1(N571), .B0(data[1]), .B1(n138), .Y(n1296) );
  AOI22X1 U143 ( .A0(n721), .A1(N570), .B0(data[0]), .B1(n139), .Y(n1297) );
  INVX1 U144 ( .A(n141), .Y(n148) );
  INVX1 U145 ( .A(n1658), .Y(n675) );
  CLKINVX3 U146 ( .A(n1266), .Y(n137) );
  INVX4 U147 ( .A(n1408), .Y(n702) );
  CLKINVX3 U148 ( .A(n730), .Y(n728) );
  OR2X2 U149 ( .A(n1191), .B(reset), .Y(n49) );
  CLKINVX3 U150 ( .A(n1301), .Y(n157) );
  OR2X2 U151 ( .A(n733), .B(reset), .Y(n50) );
  OR2X4 U152 ( .A(n725), .B(reset), .Y(n51) );
  CLKINVX3 U153 ( .A(n137), .Y(n139) );
  CLKINVX3 U154 ( .A(n137), .Y(n138) );
  INVX2 U155 ( .A(n676), .Y(n174) );
  NAND2X1 U156 ( .A(n2080), .B(n2086), .Y(n52) );
  NAND2X1 U157 ( .A(n2086), .B(n2079), .Y(n53) );
  NAND2X1 U158 ( .A(n2077), .B(n2080), .Y(n54) );
  NAND2X1 U159 ( .A(n2079), .B(n2076), .Y(n55) );
  INVX4 U160 ( .A(n709), .Y(n707) );
  INVX4 U161 ( .A(n717), .Y(n715) );
  BUFX8 U162 ( .A(n1622), .Y(n72) );
  CLKINVX3 U163 ( .A(n137), .Y(n140) );
  CLKINVX3 U164 ( .A(n1586), .Y(n684) );
  CLKINVX3 U165 ( .A(n684), .Y(n150) );
  CLKINVX3 U166 ( .A(n684), .Y(n149) );
  CLKINVX3 U167 ( .A(n1550), .Y(n687) );
  CLKINVX3 U168 ( .A(n687), .Y(n152) );
  CLKINVX3 U169 ( .A(n687), .Y(n151) );
  NOR2X2 U170 ( .A(n1443), .B(reset), .Y(n1444) );
  INVX4 U171 ( .A(n50), .Y(n732) );
  INVX4 U172 ( .A(n51), .Y(n724) );
  CLKINVX3 U173 ( .A(n158), .Y(n162) );
  CLKINVX3 U174 ( .A(n158), .Y(n161) );
  CLKINVX3 U175 ( .A(n157), .Y(n159) );
  CLKINVX3 U176 ( .A(n157), .Y(n160) );
  NAND3BX4 U177 ( .AN(n58), .B(n1692), .C(write_enable), .Y(n59) );
  INVX1 U178 ( .A(n1154), .Y(n58) );
  AOI2BB2X1 U179 ( .B0(N891), .B1(n75), .A0N(n60), .A1N(n153), .Y(n1644) );
  INVX1 U180 ( .A(N899), .Y(n60) );
  INVX1 U181 ( .A(n1116), .Y(n737) );
  CLKINVX8 U182 ( .A(n1551), .Y(n685) );
  CLKINVX8 U183 ( .A(n1587), .Y(n682) );
  AOI2BB2X2 U184 ( .B0(n154), .B1(N907), .A0N(n60), .A1N(n680), .Y(n1636) );
  AOI22X1 U185 ( .A0(n700), .A1(N707), .B0(N699), .B1(n696), .Y(n1431) );
  AOI22X1 U186 ( .A0(n154), .A1(N911), .B0(N903), .B1(n75), .Y(n1632) );
  AOI2BB2XL U187 ( .B0(data[6]), .B1(n697), .A0N(n84), .A1N(n61), .Y(n1434) );
  BUFX3 U188 ( .A(n1370), .Y(n62) );
  AOI2BB2XL U189 ( .B0(data[5]), .B1(n696), .A0N(n84), .A1N(n63), .Y(n1435) );
  AOI2BB2X1 U190 ( .B0(data[3]), .B1(n113), .A0N(n148), .A1N(n64), .Y(n1542)
         );
  OAI2BB2X1 U191 ( .B0(n66), .B1(n67), .A0N(n141), .A1N(N798), .Y(n65) );
  XOR3X2 U192 ( .A(R1[20]), .B(R1[18]), .C(R1[11]), .Y(sigma1[1]) );
  AOI2BB2XL U193 ( .B0(data[4]), .B1(n697), .A0N(n84), .A1N(n70), .Y(n1436) );
  INVXL U194 ( .A(n1657), .Y(n71) );
  INVX12 U195 ( .A(n1657), .Y(n679) );
  INVX4 U196 ( .A(n679), .Y(n677) );
  INVX20 U197 ( .A(n719), .Y(n718) );
  XOR3X2 U198 ( .A(R14[20]), .B(R14[31]), .C(R14[16]), .Y(sigma0[13]) );
  INVX1 U199 ( .A(n1477), .Y(n689) );
  INVX8 U200 ( .A(n689), .Y(n688) );
  NOR2X2 U201 ( .A(n1621), .B(reset), .Y(n1622) );
  AOI2BB2X1 U202 ( .B0(N795), .B1(n113), .A0N(n145), .A1N(n74), .Y(n1536) );
  INVX4 U203 ( .A(n1513), .Y(n145) );
  NOR2X4 U204 ( .A(n1621), .B(reset), .Y(n75) );
  INVX2 U205 ( .A(n72), .Y(n680) );
  AOI22X1 U206 ( .A0(n154), .A1(buffer[14]), .B0(N912), .B1(n72), .Y(n1623) );
  INVX12 U207 ( .A(n726), .Y(n725) );
  OAI22X1 U208 ( .A0(n84), .A1(n79), .B0(n119), .B1(n80), .Y(n78) );
  CLKINVX8 U209 ( .A(n702), .Y(n701) );
  OAI2BB2X1 U210 ( .B0(n71), .B1(n82), .A0N(N930), .A1N(n175), .Y(n81) );
  OAI2BB2X1 U211 ( .B0(n84), .B1(n85), .A0N(N698), .A1N(n1409), .Y(n83) );
  CLKINVX3 U212 ( .A(n695), .Y(n694) );
  CLKINVX3 U213 ( .A(n695), .Y(n693) );
  CLKINVX3 U214 ( .A(n1443), .Y(n695) );
  AOI22X1 U215 ( .A0(n700), .A1(N714), .B0(N706), .B1(n696), .Y(n1424) );
  INVX8 U216 ( .A(n698), .Y(n696) );
  AOI22X1 U217 ( .A0(n694), .A1(N746), .B0(N738), .B1(n690), .Y(n1459) );
  INVX8 U218 ( .A(n692), .Y(n690) );
  AOI22X1 U219 ( .A0(n678), .A1(buffer[6]), .B0(N944), .B1(n175), .Y(n1659) );
  AOI22X1 U220 ( .A0(n677), .A1(N936), .B0(N928), .B1(n1658), .Y(n1675) );
  OAI2BB2X1 U221 ( .B0(n84), .B1(n99), .A0N(data[2]), .A1N(n1409), .Y(n98) );
  OAI2BB2X1 U222 ( .B0(n695), .B1(n101), .A0N(data[2]), .A1N(n1444), .Y(n100)
         );
  OAI2BB2X1 U223 ( .B0(n84), .B1(n107), .A0N(data[1]), .A1N(n1409), .Y(n106)
         );
  OAI2BB2X1 U224 ( .B0(n695), .B1(n109), .A0N(data[1]), .A1N(n1444), .Y(n108)
         );
  CLKINVX8 U225 ( .A(n1514), .Y(n110) );
  INVX8 U226 ( .A(n110), .Y(n111) );
  AOI2BB2X1 U227 ( .B0(n142), .B1(N815), .A0N(n114), .A1N(n110), .Y(n1524) );
  OAI2BB2X1 U228 ( .B0(n117), .B1(n680), .A0N(n154), .A1N(buffer[12]), .Y(n116) );
  OAI2BB2X1 U229 ( .B0(n119), .B1(n675), .A0N(n678), .A1N(N925), .Y(n118) );
  OAI2BB2XL U230 ( .B0(n121), .B1(n680), .A0N(n154), .A1N(buffer[10]), .Y(n120) );
  INVX8 U231 ( .A(n682), .Y(n169) );
  INVX8 U232 ( .A(n685), .Y(n170) );
  OAI22XL U233 ( .A0(n679), .A1(n124), .B0(n125), .B1(n675), .Y(n123) );
  AOI2BB2X1 U234 ( .B0(n677), .B1(buffer[3]), .A0N(n126), .A1N(n676), .Y(n1662) );
  OAI22XL U235 ( .A0(n153), .A1(n128), .B0(n129), .B1(n681), .Y(n127) );
  AOI2BB2X1 U236 ( .B0(n154), .B1(N902), .A0N(n130), .A1N(n681), .Y(n1641) );
  OAI2BB2XL U237 ( .B0(n132), .B1(n681), .A0N(n154), .A1N(N904), .Y(n131) );
  AOI2BB2XL U238 ( .B0(N890), .B1(n72), .A0N(n153), .A1N(n133), .Y(n1645) );
  AOI31X2 U239 ( .A0(n1333), .A1(n190), .A2(n1334), .B0(reset), .Y(n1300) );
  AOI22X1 U240 ( .A0(n718), .A1(N624), .B0(N616), .B1(n161), .Y(n1310) );
  NAND2X4 U241 ( .A(n807), .B(n806), .Y(N2158) );
  AOI22X1 U242 ( .A0(n715), .A1(N653), .B0(N645), .B1(n711), .Y(n1349) );
  AOI22X1 U243 ( .A0(n715), .A1(N652), .B0(N644), .B1(n711), .Y(n1350) );
  AOI22X1 U244 ( .A0(n715), .A1(N651), .B0(N643), .B1(n711), .Y(n1351) );
  AOI22X1 U245 ( .A0(n715), .A1(N650), .B0(N642), .B1(n711), .Y(n1352) );
  AOI22X1 U246 ( .A0(n715), .A1(N649), .B0(N641), .B1(n711), .Y(n1353) );
  AOI22X1 U247 ( .A0(n715), .A1(N648), .B0(N640), .B1(n711), .Y(n1354) );
  AOI22X1 U248 ( .A0(n678), .A1(N922), .B0(data[0]), .B1(n175), .Y(n1689) );
  AOI22X1 U249 ( .A0(n707), .A1(N685), .B0(N677), .B1(n704), .Y(n1385) );
  AOI22X1 U250 ( .A0(n707), .A1(N684), .B0(N676), .B1(n704), .Y(n1386) );
  AOI22X1 U251 ( .A0(n707), .A1(N683), .B0(N675), .B1(n704), .Y(n1387) );
  AOI22X1 U252 ( .A0(n707), .A1(N682), .B0(N674), .B1(n704), .Y(n1388) );
  AOI22X1 U253 ( .A0(n707), .A1(N681), .B0(N673), .B1(n704), .Y(n1389) );
  AOI22X1 U254 ( .A0(n707), .A1(N680), .B0(N672), .B1(n704), .Y(n1390) );
  AOI22X2 U255 ( .A0(n678), .A1(N931), .B0(N923), .B1(n174), .Y(n1680) );
  AOI22X2 U256 ( .A0(n678), .A1(N933), .B0(N925), .B1(n174), .Y(n1678) );
  AOI22X2 U257 ( .A0(n677), .A1(N932), .B0(N924), .B1(n174), .Y(n1679) );
  AOI22X2 U258 ( .A0(n677), .A1(N940), .B0(N932), .B1(n174), .Y(n1671) );
  NAND4X2 U259 ( .A(n1334), .B(n1547), .C(n1548), .D(n1441), .Y(n1511) );
  AOI22X1 U260 ( .A0(n707), .A1(N688), .B0(N680), .B1(n704), .Y(n1382) );
  AOI22X1 U261 ( .A0(n707), .A1(N687), .B0(N679), .B1(n704), .Y(n1383) );
  AOI22X1 U262 ( .A0(n707), .A1(N686), .B0(N678), .B1(n704), .Y(n1384) );
  AOI22X1 U263 ( .A0(n678), .A1(N937), .B0(N929), .B1(n175), .Y(n1674) );
  AOI22X1 U264 ( .A0(n678), .A1(N934), .B0(N926), .B1(n175), .Y(n1677) );
  CLKINVX3 U265 ( .A(n742), .Y(n741) );
  NAND2X2 U266 ( .A(n767), .B(n766), .Y(N2146) );
  AND2X4 U267 ( .A(n1153), .B(n1298), .Y(n1406) );
  AND2X4 U268 ( .A(n1152), .B(n1225), .Y(n1298) );
  AOI31X4 U269 ( .A0(n1261), .A1(n1298), .A2(n190), .B0(reset), .Y(n1265) );
  XOR2XL U270 ( .A(R1[15]), .B(R1[17]), .Y(sigma1[30]) );
  AOI22X1 U271 ( .A0(n154), .A1(N909), .B0(N901), .B1(n72), .Y(n1634) );
  AOI22X1 U272 ( .A0(n154), .A1(N894), .B0(data[4]), .B1(n75), .Y(n1649) );
  AOI22X1 U273 ( .A0(n154), .A1(N892), .B0(data[2]), .B1(n75), .Y(n1651) );
  AOI31X4 U274 ( .A0(n190), .A1(n1156), .A2(n1441), .B0(reset), .Y(n1408) );
  AOI31X4 U275 ( .A0(n190), .A1(n1155), .A2(n1441), .B0(reset), .Y(n1443) );
  AOI22X1 U276 ( .A0(n678), .A1(buffer[0]), .B0(N938), .B1(n175), .Y(n1665) );
  NAND2X4 U277 ( .A(n819), .B(n818), .Y(N2161) );
  NAND2X2 U278 ( .A(logic_result[15]), .B(n605), .Y(n766) );
  AND2X4 U279 ( .A(n1151), .B(n1406), .Y(n1441) );
  AOI2BB1X4 U280 ( .A0N(n1546), .A1N(n1511), .B0(reset), .Y(n1513) );
  INVX4 U281 ( .A(n702), .Y(n700) );
  NAND2X4 U282 ( .A(logic_result[30]), .B(n606), .Y(n818) );
  XOR2XL U283 ( .A(R1[12]), .B(R1[14]), .Y(sigma1[27]) );
  XOR2X1 U284 ( .A(R1[10]), .B(R1[12]), .Y(sigma1[25]) );
  XOR3X2 U285 ( .A(R1[19]), .B(R1[21]), .C(R1[12]), .Y(sigma1[2]) );
  INVX8 U286 ( .A(n692), .Y(n691) );
  INVX8 U287 ( .A(n698), .Y(n697) );
  AOI22X1 U288 ( .A0(n721), .A1(N576), .B0(data[6]), .B1(n138), .Y(n1291) );
  INVX4 U289 ( .A(n1300), .Y(n719) );
  NAND2X4 U290 ( .A(logic_result[27]), .B(n606), .Y(n806) );
  AOI22XL U291 ( .A0(n725), .A1(buffer[96]), .B0(N554), .B1(n724), .Y(n1235)
         );
  INVX8 U292 ( .A(n709), .Y(n708) );
  INVX8 U293 ( .A(n717), .Y(n716) );
  INVX2 U294 ( .A(n145), .Y(n141) );
  BUFX3 U295 ( .A(n143), .Y(n142) );
  INVX1 U296 ( .A(n145), .Y(n143) );
  BUFX3 U297 ( .A(n143), .Y(n144) );
  INVX8 U298 ( .A(n145), .Y(n146) );
  INVXL U299 ( .A(n145), .Y(n147) );
  AOI31X4 U300 ( .A0(n1547), .A1(n1619), .A2(n1584), .B0(reset), .Y(n1586) );
  INVX4 U301 ( .A(n684), .Y(n683) );
  AOI31X4 U302 ( .A0(n1547), .A1(n1583), .A2(n1584), .B0(reset), .Y(n1550) );
  INVX4 U303 ( .A(n687), .Y(n686) );
  INVXL U304 ( .A(n153), .Y(n155) );
  INVX8 U305 ( .A(n679), .Y(n678) );
  XOR3X4 U306 ( .A(R14[20]), .B(R14[9]), .C(R14[5]), .Y(sigma0[2]) );
  INVX1 U307 ( .A(n157), .Y(n156) );
  CLKINVX2 U308 ( .A(n1301), .Y(n158) );
  XOR2XL U309 ( .A(R14[6]), .B(R14[17]), .Y(sigma0[31]) );
  XOR2XL U310 ( .A(R14[4]), .B(R14[15]), .Y(sigma0[29]) );
  XOR3X2 U311 ( .A(R14[25]), .B(R14[14]), .C(R14[10]), .Y(sigma0[7]) );
  XOR2XL U312 ( .A(R14[5]), .B(R14[16]), .Y(sigma0[30]) );
  XOR2X1 U313 ( .A(R1[16]), .B(R1[18]), .Y(sigma1[31]) );
  XOR3X4 U314 ( .A(R14[18]), .B(R14[29]), .C(R14[14]), .Y(sigma0[11]) );
  XOR3X2 U315 ( .A(R1[22]), .B(R1[24]), .C(R1[15]), .Y(sigma1[5]) );
  CLKINVX2 U316 ( .A(n77), .Y(n676) );
  INVX4 U317 ( .A(n51), .Y(n723) );
  INVX4 U318 ( .A(n50), .Y(n731) );
  CLKINVX3 U319 ( .A(n1373), .Y(n706) );
  INVX4 U320 ( .A(n714), .Y(n710) );
  CLKINVX3 U321 ( .A(n1337), .Y(n714) );
  INVX4 U322 ( .A(n1372), .Y(n709) );
  INVX4 U323 ( .A(n1336), .Y(n717) );
  NOR3X1 U324 ( .A(n1654), .B(counter1[6]), .C(n1690), .Y(n1547) );
  INVX2 U325 ( .A(n1115), .Y(n742) );
  INVXL U326 ( .A(n1227), .Y(n726) );
  INVXL U327 ( .A(n1158), .Y(n734) );
  INVXL U328 ( .A(n1115), .Y(n743) );
  NAND2XL U329 ( .A(n1700), .B(n1704), .Y(n1619) );
  NAND2XL U330 ( .A(n1704), .B(n1694), .Y(n1583) );
  NAND2XL U331 ( .A(n1693), .B(n1701), .Y(n1695) );
  AND3X2 U332 ( .A(n1691), .B(n1548), .C(n1547), .Y(n190) );
  AND2X1 U333 ( .A(n1701), .B(n1702), .Y(n1510) );
  AND2X1 U334 ( .A(n1699), .B(n1701), .Y(n1369) );
  AND2X1 U335 ( .A(n1703), .B(n1704), .Y(n1690) );
  AND2X1 U336 ( .A(n1699), .B(n1703), .Y(n1405) );
  NOR2X4 U337 ( .A(n718), .B(reset), .Y(n1301) );
  AOI22XL U338 ( .A0(n718), .A1(N625), .B0(N617), .B1(n156), .Y(n1309) );
  AOI22XL U339 ( .A0(n693), .A1(N753), .B0(N745), .B1(n690), .Y(n1452) );
  AOI22XL U340 ( .A0(n699), .A1(N721), .B0(N713), .B1(n696), .Y(n1417) );
  AOI22XL U341 ( .A0(n693), .A1(buffer[55]), .B0(N753), .B1(n691), .Y(n1442)
         );
  AOI22XL U342 ( .A0(n699), .A1(buffer[63]), .B0(N721), .B1(n697), .Y(n1407)
         );
  AOI22XL U343 ( .A0(n707), .A1(N689), .B0(N681), .B1(n704), .Y(n1381) );
  AOI22XL U344 ( .A0(n715), .A1(N657), .B0(N649), .B1(n711), .Y(n1345) );
  AOI22XL U345 ( .A0(n715), .A1(buffer[79]), .B0(N657), .B1(n712), .Y(n1335)
         );
  AOI22XL U346 ( .A0(n707), .A1(buffer[71]), .B0(N689), .B1(n703), .Y(n1371)
         );
  AOI22XL U347 ( .A0(n678), .A1(N945), .B0(N937), .B1(n175), .Y(n1666) );
  AOI22XL U348 ( .A0(n155), .A1(N913), .B0(N905), .B1(n75), .Y(n1630) );
  AOI22XL U349 ( .A0(n683), .A1(N881), .B0(N873), .B1(n169), .Y(n1595) );
  AOI22XL U350 ( .A0(n686), .A1(N849), .B0(N841), .B1(n170), .Y(n1559) );
  AOI22XL U351 ( .A0(n142), .A1(N817), .B0(N809), .B1(n112), .Y(n1522) );
  AOI22XL U352 ( .A0(n688), .A1(N785), .B0(N777), .B1(n172), .Y(n1486) );
  AOI22XL U353 ( .A0(n693), .A1(N741), .B0(N733), .B1(n691), .Y(n1464) );
  AOI22XL U354 ( .A0(n700), .A1(N709), .B0(N701), .B1(n697), .Y(n1429) );
  AOI22XL U355 ( .A0(n707), .A1(N677), .B0(N669), .B1(n703), .Y(n1393) );
  AOI22XL U356 ( .A0(n715), .A1(N645), .B0(N637), .B1(n710), .Y(n1357) );
  AOI22XL U357 ( .A0(n718), .A1(N613), .B0(N605), .B1(n160), .Y(n1321) );
  AOI22XL U358 ( .A0(n725), .A1(N545), .B0(data[7]), .B1(n723), .Y(n1252) );
  AOI22XL U359 ( .A0(n725), .A1(N544), .B0(data[6]), .B1(n723), .Y(n1253) );
  AOI22XL U360 ( .A0(n725), .A1(N543), .B0(data[5]), .B1(n724), .Y(n1254) );
  AOI22XL U361 ( .A0(n725), .A1(N542), .B0(data[4]), .B1(n723), .Y(n1255) );
  AOI22XL U362 ( .A0(n725), .A1(N541), .B0(data[3]), .B1(n724), .Y(n1256) );
  AOI22XL U363 ( .A0(n725), .A1(N540), .B0(data[2]), .B1(n724), .Y(n1257) );
  AOI22XL U364 ( .A0(n725), .A1(N539), .B0(data[1]), .B1(n723), .Y(n1258) );
  AOI22XL U365 ( .A0(n725), .A1(N538), .B0(data[0]), .B1(n724), .Y(n1259) );
  AOI22XL U366 ( .A0(n728), .A1(N513), .B0(data[7]), .B1(n727), .Y(n1216) );
  AOI22XL U367 ( .A0(n728), .A1(N512), .B0(data[6]), .B1(n727), .Y(n1217) );
  AOI22XL U368 ( .A0(n728), .A1(N511), .B0(data[5]), .B1(n727), .Y(n1218) );
  AOI22XL U369 ( .A0(n728), .A1(N510), .B0(data[4]), .B1(n727), .Y(n1219) );
  AOI22XL U370 ( .A0(n728), .A1(N509), .B0(data[3]), .B1(n727), .Y(n1220) );
  AOI22XL U371 ( .A0(n728), .A1(N508), .B0(data[2]), .B1(n727), .Y(n1221) );
  AOI22XL U372 ( .A0(n728), .A1(N507), .B0(data[1]), .B1(n727), .Y(n1222) );
  AOI22XL U374 ( .A0(n728), .A1(N506), .B0(data[0]), .B1(n727), .Y(n1223) );
  AOI22XL U375 ( .A0(n733), .A1(N481), .B0(data[7]), .B1(n732), .Y(n1183) );
  AOI22XL U376 ( .A0(n733), .A1(N480), .B0(data[6]), .B1(n732), .Y(n1184) );
  AOI22XL U377 ( .A0(n733), .A1(N479), .B0(data[5]), .B1(n731), .Y(n1185) );
  AOI22XL U378 ( .A0(n733), .A1(N478), .B0(data[4]), .B1(n732), .Y(n1186) );
  AOI22XL U379 ( .A0(n733), .A1(N477), .B0(data[3]), .B1(n731), .Y(n1187) );
  AOI22XL U380 ( .A0(n733), .A1(N476), .B0(data[2]), .B1(n732), .Y(n1188) );
  AOI22XL U381 ( .A0(n733), .A1(N475), .B0(data[1]), .B1(n732), .Y(n1189) );
  AOI22XL U382 ( .A0(n733), .A1(N474), .B0(data[0]), .B1(n731), .Y(n1697) );
  AOI22XL U383 ( .A0(n741), .A1(N449), .B0(data[7]), .B1(n735), .Y(n1140) );
  AOI22XL U384 ( .A0(n741), .A1(N448), .B0(data[6]), .B1(n735), .Y(n1141) );
  AOI22XL U385 ( .A0(n741), .A1(N447), .B0(data[5]), .B1(n735), .Y(n1142) );
  AOI22XL U386 ( .A0(n741), .A1(N446), .B0(data[4]), .B1(n735), .Y(n1143) );
  AOI22XL U387 ( .A0(n741), .A1(N445), .B0(data[3]), .B1(n735), .Y(n1144) );
  AOI22XL U388 ( .A0(n741), .A1(N444), .B0(data[2]), .B1(n735), .Y(n1145) );
  AOI22XL U389 ( .A0(n741), .A1(N443), .B0(data[1]), .B1(n735), .Y(n1146) );
  AOI22XL U390 ( .A0(n741), .A1(N442), .B0(data[0]), .B1(n735), .Y(n1147) );
  NOR2XL U391 ( .A(counter1[4]), .B(counter1[5]), .Y(n1693) );
  NOR2XL U392 ( .A(counter1[2]), .B(counter1[3]), .Y(n1700) );
  NOR2XL U393 ( .A(n1055), .B(counter1[3]), .Y(n1694) );
  NOR2XL U394 ( .A(n1054), .B(counter1[4]), .Y(n1702) );
  XOR2XL U395 ( .A(R1[8]), .B(R1[10]), .Y(sigma1[23]) );
  XOR2XL U396 ( .A(R1[9]), .B(R1[11]), .Y(sigma1[24]) );
  AND2X1 U397 ( .A(counter1[4]), .B(n1054), .Y(n1699) );
  NAND3XL U398 ( .A(n1062), .B(n2087), .C(inner_busy), .Y(n2070) );
  AND3X1 U399 ( .A(n1706), .B(n1062), .C(inner_busy), .Y(n1705) );
  INVX1 U400 ( .A(n666), .Y(n614) );
  INVX1 U401 ( .A(n666), .Y(n615) );
  INVX1 U402 ( .A(n666), .Y(n616) );
  INVX1 U403 ( .A(n666), .Y(n617) );
  INVX1 U404 ( .A(n665), .Y(n618) );
  INVX1 U405 ( .A(n665), .Y(n619) );
  INVX1 U406 ( .A(n664), .Y(n620) );
  INVX1 U408 ( .A(n664), .Y(n621) );
  INVX1 U409 ( .A(n664), .Y(n622) );
  INVX1 U410 ( .A(n665), .Y(n623) );
  INVX1 U411 ( .A(n663), .Y(n624) );
  INVX1 U412 ( .A(n663), .Y(n625) );
  INVX1 U413 ( .A(n663), .Y(n626) );
  INVX1 U414 ( .A(n662), .Y(n627) );
  INVX1 U415 ( .A(n662), .Y(n628) );
  INVX1 U416 ( .A(n662), .Y(n629) );
  INVX1 U417 ( .A(n661), .Y(n630) );
  INVX1 U418 ( .A(n661), .Y(n631) );
  INVX1 U419 ( .A(n660), .Y(n632) );
  INVX1 U420 ( .A(n660), .Y(n633) );
  INVX1 U421 ( .A(n660), .Y(n634) );
  INVX1 U422 ( .A(n661), .Y(n635) );
  INVX1 U423 ( .A(n659), .Y(n636) );
  INVX1 U424 ( .A(n659), .Y(n637) );
  INVX1 U425 ( .A(n658), .Y(n638) );
  INVX1 U426 ( .A(n658), .Y(n639) );
  INVX1 U427 ( .A(n658), .Y(n640) );
  INVX1 U428 ( .A(n659), .Y(n641) );
  INVX1 U429 ( .A(n657), .Y(n642) );
  INVX1 U430 ( .A(n657), .Y(n643) );
  INVX1 U431 ( .A(n656), .Y(n644) );
  INVX1 U432 ( .A(n656), .Y(n645) );
  INVX1 U433 ( .A(n657), .Y(n646) );
  INVX1 U434 ( .A(n656), .Y(n647) );
  INVX1 U435 ( .A(n655), .Y(n648) );
  INVX1 U436 ( .A(n655), .Y(n649) );
  INVX1 U437 ( .A(n654), .Y(n650) );
  INVX1 U438 ( .A(n654), .Y(n651) );
  INVX1 U439 ( .A(n654), .Y(n652) );
  INVX1 U440 ( .A(n655), .Y(n653) );
  INVX1 U442 ( .A(n612), .Y(n666) );
  INVX1 U443 ( .A(n612), .Y(n665) );
  INVX1 U444 ( .A(n612), .Y(n664) );
  INVX1 U445 ( .A(n611), .Y(n663) );
  INVX1 U446 ( .A(n611), .Y(n662) );
  INVX1 U447 ( .A(n610), .Y(n661) );
  INVX1 U448 ( .A(n610), .Y(n660) );
  INVX1 U449 ( .A(n609), .Y(n659) );
  INVX1 U450 ( .A(n609), .Y(n658) );
  INVX1 U451 ( .A(n608), .Y(n657) );
  INVX1 U452 ( .A(n608), .Y(n656) );
  INVX1 U453 ( .A(n607), .Y(n606) );
  INVX1 U454 ( .A(n613), .Y(n612) );
  INVX1 U455 ( .A(n613), .Y(n611) );
  INVX1 U456 ( .A(n613), .Y(n610) );
  INVX1 U457 ( .A(n613), .Y(n609) );
  INVX1 U458 ( .A(n613), .Y(n608) );
  INVX1 U459 ( .A(n611), .Y(n655) );
  INVX1 U460 ( .A(n610), .Y(n654) );
  INVX1 U461 ( .A(n53), .Y(n670) );
  INVX1 U462 ( .A(n52), .Y(n668) );
  INVX1 U463 ( .A(n54), .Y(n672) );
  INVX1 U464 ( .A(n55), .Y(n674) );
  NAND3XL U465 ( .A(n190), .B(n1406), .C(n1334), .Y(n1370) );
  INVX1 U466 ( .A(n722), .Y(n720) );
  INVX1 U467 ( .A(n730), .Y(n729) );
  INVX1 U468 ( .A(n742), .Y(n740) );
  NOR2X1 U469 ( .A(n1369), .B(n1405), .Y(n1151) );
  BUFX3 U470 ( .A(n820), .Y(n604) );
  INVX1 U471 ( .A(n760), .Y(n820) );
  INVX1 U472 ( .A(n607), .Y(n605) );
  INVX1 U473 ( .A(n545), .Y(n607) );
  INVX1 U474 ( .A(n2196), .Y(n613) );
  AND3X2 U475 ( .A(n1151), .B(n1696), .C(n1334), .Y(n1261) );
  NOR2X1 U476 ( .A(n1510), .B(n1546), .Y(n1691) );
  AND3X2 U477 ( .A(n1261), .B(n1695), .C(n1263), .Y(n1224) );
  INVX1 U478 ( .A(n53), .Y(n669) );
  INVX1 U479 ( .A(n52), .Y(n667) );
  INVX1 U480 ( .A(n54), .Y(n671) );
  INVX1 U481 ( .A(n55), .Y(n673) );
  INVX1 U482 ( .A(n1116), .Y(n738) );
  NAND2X1 U483 ( .A(n811), .B(n810), .Y(N2159) );
  OAI21XL U484 ( .A0(n809), .A1(n808), .B0(n604), .Y(n811) );
  NAND2X1 U485 ( .A(logic_result[28]), .B(n606), .Y(n810) );
  NAND4X1 U486 ( .A(n1763), .B(n1764), .C(n1761), .D(n1762), .Y(n809) );
  OAI21XL U487 ( .A0(n817), .A1(n816), .B0(n604), .Y(n819) );
  NAND4X1 U488 ( .A(n1741), .B(n1742), .C(n1739), .D(n1740), .Y(n817) );
  NAND2X1 U489 ( .A(n791), .B(n790), .Y(N2154) );
  OAI21XL U490 ( .A0(n789), .A1(n788), .B0(n604), .Y(n791) );
  NAND4X1 U491 ( .A(n1818), .B(n1819), .C(n1816), .D(n1817), .Y(n789) );
  NAND2X1 U492 ( .A(n799), .B(n798), .Y(N2156) );
  OAI21XL U493 ( .A0(n797), .A1(n796), .B0(n604), .Y(n799) );
  NAND2X1 U494 ( .A(logic_result[25]), .B(n606), .Y(n798) );
  NAND4X1 U495 ( .A(n1796), .B(n1797), .C(n1794), .D(n1795), .Y(n797) );
  NAND2X1 U496 ( .A(n803), .B(n802), .Y(N2157) );
  OAI21XL U497 ( .A0(n801), .A1(n800), .B0(n604), .Y(n803) );
  NAND2X1 U498 ( .A(logic_result[26]), .B(n606), .Y(n802) );
  NAND4X1 U499 ( .A(n1785), .B(n1786), .C(n1783), .D(n1784), .Y(n801) );
  OAI21XL U500 ( .A0(n805), .A1(n804), .B0(n604), .Y(n807) );
  NAND4X1 U501 ( .A(n1774), .B(n1775), .C(n1772), .D(n1773), .Y(n805) );
  OAI21XL U502 ( .A0(n813), .A1(n812), .B0(n604), .Y(n815) );
  NAND4X1 U503 ( .A(n1752), .B(n1753), .C(n1750), .D(n1751), .Y(n813) );
  NAND2X1 U504 ( .A(n824), .B(n823), .Y(N2162) );
  OAI21XL U505 ( .A0(n822), .A1(n821), .B0(n604), .Y(n824) );
  NAND2X1 U506 ( .A(logic_result[31]), .B(n605), .Y(n823) );
  NAND4X1 U507 ( .A(n1715), .B(n1716), .C(n1713), .D(n1714), .Y(n822) );
  OAI2BB2X1 U508 ( .B0(n757), .B1(n760), .A0N(logic_result[10]), .A1N(n606), 
        .Y(N2141) );
  NOR2X1 U509 ( .A(n1957), .B(n1958), .Y(n757) );
  NAND4X1 U510 ( .A(n1959), .B(n1960), .C(n1961), .D(n1962), .Y(n1958) );
  INVX1 U511 ( .A(n743), .Y(n739) );
  NAND2X1 U512 ( .A(n773), .B(n772), .Y(N2149) );
  OAI21XL U513 ( .A0(n1870), .A1(n1869), .B0(n604), .Y(n773) );
  NAND2X1 U514 ( .A(logic_result[18]), .B(n605), .Y(n772) );
  NAND4X1 U515 ( .A(n1871), .B(n1872), .C(n1873), .D(n1874), .Y(n1870) );
  NAND2X1 U516 ( .A(n795), .B(n794), .Y(N2155) );
  OAI21XL U517 ( .A0(n793), .A1(n792), .B0(n604), .Y(n795) );
  NAND2X1 U518 ( .A(logic_result[24]), .B(n606), .Y(n794) );
  NAND4X1 U519 ( .A(n1807), .B(n1808), .C(n1805), .D(n1806), .Y(n793) );
  NAND2X1 U520 ( .A(n763), .B(n762), .Y(N2144) );
  OAI21XL U521 ( .A0(n1925), .A1(n1924), .B0(n604), .Y(n763) );
  NAND2X1 U522 ( .A(logic_result[13]), .B(n605), .Y(n762) );
  NAND4X1 U523 ( .A(n1926), .B(n1927), .C(n1928), .D(n1929), .Y(n1925) );
  NAND2X1 U524 ( .A(n765), .B(n764), .Y(N2145) );
  OAI21XL U525 ( .A0(n1914), .A1(n1913), .B0(n604), .Y(n765) );
  NAND2X1 U526 ( .A(logic_result[14]), .B(n605), .Y(n764) );
  NAND4X1 U527 ( .A(n1915), .B(n1916), .C(n1917), .D(n1918), .Y(n1914) );
  NAND2X1 U528 ( .A(n769), .B(n768), .Y(N2147) );
  OAI21XL U529 ( .A0(n1892), .A1(n1891), .B0(n604), .Y(n769) );
  NAND2X1 U530 ( .A(logic_result[16]), .B(n605), .Y(n768) );
  NAND4X1 U531 ( .A(n1893), .B(n1894), .C(n1895), .D(n1896), .Y(n1892) );
  NAND2X1 U532 ( .A(n759), .B(n758), .Y(N2142) );
  OAI21XL U533 ( .A0(n1947), .A1(n1946), .B0(n604), .Y(n759) );
  NAND2X1 U534 ( .A(logic_result[11]), .B(n605), .Y(n758) );
  NAND4X1 U535 ( .A(n1948), .B(n1949), .C(n1950), .D(n1951), .Y(n1947) );
  OAI21XL U536 ( .A0(n1903), .A1(n1902), .B0(n604), .Y(n767) );
  NAND4X1 U537 ( .A(n1904), .B(n1905), .C(n1906), .D(n1907), .Y(n1903) );
  NAND2X1 U538 ( .A(n771), .B(n770), .Y(N2148) );
  OAI21XL U539 ( .A0(n1881), .A1(n1880), .B0(n604), .Y(n771) );
  NAND2X1 U540 ( .A(logic_result[17]), .B(n605), .Y(n770) );
  NAND4X1 U541 ( .A(n1882), .B(n1883), .C(n1884), .D(n1885), .Y(n1881) );
  NAND2X1 U542 ( .A(n775), .B(n774), .Y(N2150) );
  OAI21XL U543 ( .A0(n1859), .A1(n1858), .B0(n604), .Y(n775) );
  NAND2X1 U544 ( .A(logic_result[19]), .B(n605), .Y(n774) );
  NAND4X1 U545 ( .A(n1860), .B(n1861), .C(n1862), .D(n1863), .Y(n1859) );
  NAND2X1 U546 ( .A(n779), .B(n778), .Y(N2151) );
  OAI21XL U547 ( .A0(n777), .A1(n776), .B0(n604), .Y(n779) );
  NAND2X1 U548 ( .A(logic_result[20]), .B(n605), .Y(n778) );
  NAND4X1 U549 ( .A(n1851), .B(n1852), .C(n1849), .D(n1850), .Y(n777) );
  NAND2X1 U550 ( .A(n783), .B(n782), .Y(N2152) );
  OAI21XL U551 ( .A0(n781), .A1(n780), .B0(n604), .Y(n783) );
  NAND2X1 U552 ( .A(logic_result[21]), .B(n605), .Y(n782) );
  NAND4X1 U553 ( .A(n1840), .B(n1841), .C(n1838), .D(n1839), .Y(n781) );
  NAND2X1 U554 ( .A(n787), .B(n786), .Y(N2153) );
  OAI21XL U555 ( .A0(n785), .A1(n784), .B0(n604), .Y(n787) );
  NAND2X1 U556 ( .A(logic_result[22]), .B(n605), .Y(n786) );
  NAND4X1 U557 ( .A(n1829), .B(n1830), .C(n1827), .D(n1828), .Y(n785) );
  INVX1 U558 ( .A(n2070), .Y(n2196) );
  INVX1 U559 ( .A(n2070), .Y(n745) );
  NAND2X1 U560 ( .A(n1699), .B(n1700), .Y(n1263) );
  NAND2X1 U561 ( .A(n1693), .B(n1703), .Y(n1262) );
  NAND2X1 U562 ( .A(n744), .B(n745), .Y(n760) );
  INVX1 U563 ( .A(n746), .Y(n744) );
  AND2X2 U564 ( .A(n746), .B(n745), .Y(n545) );
  NAND2X1 U565 ( .A(n1693), .B(n1694), .Y(n1154) );
  OAI2BB2X1 U566 ( .B0(n747), .B1(n760), .A0N(logic_result[0]), .A1N(n605), 
        .Y(N2131) );
  NOR2X1 U567 ( .A(n2067), .B(n2068), .Y(n747) );
  OAI2BB2X1 U568 ( .B0(n748), .B1(n760), .A0N(logic_result[1]), .A1N(n605), 
        .Y(N2132) );
  NOR2X1 U569 ( .A(n2056), .B(n2057), .Y(n748) );
  NAND4X1 U570 ( .A(n2058), .B(n2059), .C(n2060), .D(n2061), .Y(n2057) );
  OAI2BB2X1 U571 ( .B0(n749), .B1(n760), .A0N(logic_result[2]), .A1N(n605), 
        .Y(N2133) );
  NOR2X1 U572 ( .A(n2045), .B(n2046), .Y(n749) );
  NAND4X1 U573 ( .A(n2047), .B(n2048), .C(n2049), .D(n2050), .Y(n2046) );
  OAI2BB2X1 U574 ( .B0(n750), .B1(n760), .A0N(logic_result[3]), .A1N(n545), 
        .Y(N2134) );
  NOR2X1 U575 ( .A(n2034), .B(n2035), .Y(n750) );
  NAND4X1 U576 ( .A(n2036), .B(n2037), .C(n2038), .D(n2039), .Y(n2035) );
  OAI2BB2X1 U577 ( .B0(n751), .B1(n760), .A0N(logic_result[4]), .A1N(n606), 
        .Y(N2135) );
  NOR2X1 U579 ( .A(n2023), .B(n2024), .Y(n751) );
  NAND4X1 U580 ( .A(n2025), .B(n2026), .C(n2027), .D(n2028), .Y(n2024) );
  OAI2BB2X1 U581 ( .B0(n752), .B1(n760), .A0N(logic_result[5]), .A1N(n606), 
        .Y(N2136) );
  NOR2X1 U582 ( .A(n2012), .B(n2013), .Y(n752) );
  NAND4X1 U583 ( .A(n2014), .B(n2015), .C(n2016), .D(n2017), .Y(n2013) );
  OAI2BB2X1 U584 ( .B0(n753), .B1(n760), .A0N(logic_result[6]), .A1N(n606), 
        .Y(N2137) );
  NOR2X1 U585 ( .A(n2001), .B(n2002), .Y(n753) );
  NAND4X1 U586 ( .A(n2003), .B(n2004), .C(n2005), .D(n2006), .Y(n2002) );
  OAI2BB2X1 U587 ( .B0(n754), .B1(n760), .A0N(logic_result[7]), .A1N(n606), 
        .Y(N2138) );
  NOR2X1 U588 ( .A(n1990), .B(n1991), .Y(n754) );
  NAND4X1 U589 ( .A(n1992), .B(n1993), .C(n1994), .D(n1995), .Y(n1991) );
  OAI2BB2X1 U590 ( .B0(n755), .B1(n760), .A0N(logic_result[8]), .A1N(n606), 
        .Y(N2139) );
  NOR2X1 U591 ( .A(n1979), .B(n1980), .Y(n755) );
  NAND4X1 U592 ( .A(n1981), .B(n1982), .C(n1983), .D(n1984), .Y(n1980) );
  OAI2BB2X1 U593 ( .B0(n756), .B1(n760), .A0N(logic_result[9]), .A1N(n606), 
        .Y(N2140) );
  NOR2X1 U594 ( .A(n1968), .B(n1969), .Y(n756) );
  NAND4X1 U595 ( .A(n1970), .B(n1971), .C(n1972), .D(n1973), .Y(n1969) );
  OAI2BB2X1 U596 ( .B0(n761), .B1(n760), .A0N(logic_result[12]), .A1N(n606), 
        .Y(N2143) );
  NOR2X1 U597 ( .A(n1935), .B(n1936), .Y(n761) );
  NAND4X1 U598 ( .A(n1937), .B(n1938), .C(n1939), .D(n1940), .Y(n1936) );
  NAND2X1 U599 ( .A(n1693), .B(n1700), .Y(n1692) );
  NAND2X1 U600 ( .A(n1699), .B(n1694), .Y(n1696) );
  NAND2X1 U601 ( .A(n1702), .B(n1694), .Y(n1156) );
  NAND2X1 U602 ( .A(n1700), .B(n1702), .Y(n1155) );
  AND3X1 U603 ( .A(n1298), .B(n1263), .C(n1151), .Y(n1333) );
  AOI31X1 U604 ( .A0(n1698), .A1(n190), .A2(n1224), .B0(reset), .Y(n1158) );
  AND3X1 U605 ( .A(n1692), .B(n1262), .C(write_enable), .Y(n1698) );
  AOI31X1 U606 ( .A0(n1260), .A1(n190), .A2(n1261), .B0(reset), .Y(n1227) );
  AND3X1 U607 ( .A(n1262), .B(n1263), .C(n1225), .Y(n1260) );
  AOI2BB1X1 U608 ( .A0N(n1148), .A1N(n1149), .B0(reset), .Y(n1115) );
  NAND4X1 U609 ( .A(n190), .B(n1151), .C(n1152), .D(n1153), .Y(n1149) );
  NAND4XL U610 ( .A(write_enable), .B(n1154), .C(n1155), .D(n1156), .Y(n1148)
         );
  XOR3X2 U611 ( .A(R14[21]), .B(R14[17]), .C(R14[0]), .Y(sigma0[14]) );
  XOR3X2 U613 ( .A(R14[26]), .B(R14[15]), .C(R14[11]), .Y(sigma0[8]) );
  XOR3X2 U614 ( .A(R14[19]), .B(R14[8]), .C(R14[4]), .Y(sigma0[1]) );
  XOR3X2 U615 ( .A(R14[18]), .B(R14[7]), .C(R14[3]), .Y(sigma0[0]) );
  XOR3X2 U616 ( .A(R14[23]), .B(R14[12]), .C(R14[8]), .Y(sigma0[5]) );
  XOR3X2 U617 ( .A(R14[22]), .B(R14[11]), .C(R14[7]), .Y(sigma0[4]) );
  XOR3X2 U618 ( .A(R14[24]), .B(R14[13]), .C(R14[9]), .Y(sigma0[6]) );
  XOR3X2 U619 ( .A(R14[18]), .B(R14[22]), .C(R14[1]), .Y(sigma0[15]) );
  XOR3X2 U620 ( .A(R1[19]), .B(R1[17]), .C(R1[10]), .Y(sigma1[0]) );
  XOR3X2 U621 ( .A(R1[28]), .B(R1[30]), .C(R1[21]), .Y(sigma1[11]) );
  XOR3X2 U622 ( .A(R1[23]), .B(R1[30]), .C(R1[0]), .Y(sigma1[13]) );
  XOR3X2 U623 ( .A(R1[24]), .B(R1[31]), .C(R1[1]), .Y(sigma1[14]) );
  XOR3X2 U624 ( .A(R1[21]), .B(R1[23]), .C(R1[14]), .Y(sigma1[4]) );
  XOR3X2 U625 ( .A(R1[25]), .B(R1[27]), .C(R1[18]), .Y(sigma1[8]) );
  XOR3X2 U626 ( .A(R1[24]), .B(R1[26]), .C(R1[17]), .Y(sigma1[7]) );
  XOR3X2 U627 ( .A(R1[26]), .B(R1[28]), .C(R1[19]), .Y(sigma1[9]) );
  INVX1 U628 ( .A(n1666), .Y(n2184) );
  INVX1 U629 ( .A(n1667), .Y(n2185) );
  AOI22XL U630 ( .A0(n678), .A1(N944), .B0(N936), .B1(n175), .Y(n1667) );
  INVX1 U631 ( .A(n1668), .Y(n2186) );
  INVX1 U632 ( .A(n1670), .Y(n2187) );
  INVX1 U633 ( .A(n1671), .Y(n2188) );
  INVX1 U634 ( .A(n1674), .Y(n2189) );
  INVX1 U635 ( .A(n1683), .Y(n2175) );
  AOI22XL U636 ( .A0(n678), .A1(N928), .B0(data[6]), .B1(n1658), .Y(n1683) );
  AOI22XL U637 ( .A0(n678), .A1(N927), .B0(data[5]), .B1(n1658), .Y(n1684) );
  INVX1 U638 ( .A(n1685), .Y(n2177) );
  AOI22XL U639 ( .A0(n678), .A1(N926), .B0(data[4]), .B1(n1658), .Y(n1685) );
  AOI22XL U640 ( .A0(n678), .A1(N924), .B0(data[2]), .B1(n1658), .Y(n1687) );
  INVX1 U641 ( .A(n1688), .Y(n2179) );
  AOI22XL U642 ( .A0(n678), .A1(N923), .B0(data[1]), .B1(n175), .Y(n1688) );
  INVX1 U643 ( .A(n1689), .Y(n2198) );
  INVX1 U644 ( .A(n1595), .Y(n2132) );
  INVX1 U645 ( .A(n1596), .Y(n2133) );
  AOI22XL U646 ( .A0(n683), .A1(N880), .B0(N872), .B1(n169), .Y(n1596) );
  INVX1 U648 ( .A(n1597), .Y(n2134) );
  AOI22XL U649 ( .A0(n683), .A1(N879), .B0(N871), .B1(n169), .Y(n1597) );
  INVX1 U650 ( .A(n1598), .Y(n2135) );
  AOI22XL U651 ( .A0(n149), .A1(N878), .B0(N870), .B1(n169), .Y(n1598) );
  INVX1 U652 ( .A(n1599), .Y(n2136) );
  AOI22XL U653 ( .A0(n149), .A1(N877), .B0(N869), .B1(n169), .Y(n1599) );
  INVX1 U654 ( .A(n1600), .Y(n2137) );
  AOI22XL U655 ( .A0(n150), .A1(N876), .B0(N868), .B1(n169), .Y(n1600) );
  INVX1 U656 ( .A(n1601), .Y(n2138) );
  AOI22XL U657 ( .A0(n683), .A1(N875), .B0(N867), .B1(n169), .Y(n1601) );
  INVX1 U658 ( .A(n1602), .Y(n2139) );
  AOI22XL U659 ( .A0(n150), .A1(N874), .B0(N866), .B1(n169), .Y(n1602) );
  INVX1 U660 ( .A(n1603), .Y(n2140) );
  AOI22XL U661 ( .A0(n683), .A1(N873), .B0(N865), .B1(n169), .Y(n1603) );
  INVX1 U662 ( .A(n1604), .Y(n2141) );
  AOI22XL U663 ( .A0(n149), .A1(N872), .B0(N864), .B1(n169), .Y(n1604) );
  INVX1 U664 ( .A(n1605), .Y(n2142) );
  AOI22XL U665 ( .A0(n150), .A1(N871), .B0(N863), .B1(n169), .Y(n1605) );
  INVX1 U666 ( .A(n1606), .Y(n2143) );
  AOI22XL U667 ( .A0(n683), .A1(N870), .B0(N862), .B1(n169), .Y(n1606) );
  INVX1 U668 ( .A(n1607), .Y(n2144) );
  AOI22XL U669 ( .A0(n683), .A1(N869), .B0(N861), .B1(n169), .Y(n1607) );
  INVX1 U670 ( .A(n1608), .Y(n2145) );
  AOI22XL U671 ( .A0(n683), .A1(N868), .B0(N860), .B1(n169), .Y(n1608) );
  INVX1 U672 ( .A(n1609), .Y(n2146) );
  AOI22XL U673 ( .A0(n149), .A1(N867), .B0(N859), .B1(n169), .Y(n1609) );
  INVX1 U674 ( .A(n1610), .Y(n2147) );
  AOI22XL U675 ( .A0(n150), .A1(N866), .B0(N858), .B1(n169), .Y(n1610) );
  INVX1 U676 ( .A(n1611), .Y(n2117) );
  AOI22XL U677 ( .A0(n683), .A1(N865), .B0(data[7]), .B1(n169), .Y(n1611) );
  INVX1 U678 ( .A(n1612), .Y(n2118) );
  AOI22XL U679 ( .A0(n149), .A1(N864), .B0(data[6]), .B1(n169), .Y(n1612) );
  INVX1 U684 ( .A(n1613), .Y(n2119) );
  AOI22XL U685 ( .A0(n150), .A1(N863), .B0(data[5]), .B1(n169), .Y(n1613) );
  INVX1 U686 ( .A(n1614), .Y(n2120) );
  AOI22XL U687 ( .A0(n683), .A1(N862), .B0(data[4]), .B1(n169), .Y(n1614) );
  INVX1 U688 ( .A(n1615), .Y(n2121) );
  AOI22XL U691 ( .A0(n150), .A1(N861), .B0(data[3]), .B1(n169), .Y(n1615) );
  INVX1 U692 ( .A(n1616), .Y(n2122) );
  AOI22XL U693 ( .A0(n683), .A1(N860), .B0(data[2]), .B1(n169), .Y(n1616) );
  INVX1 U694 ( .A(n1617), .Y(n2123) );
  AOI22XL U695 ( .A0(n683), .A1(N859), .B0(data[1]), .B1(n169), .Y(n1617) );
  INVX1 U696 ( .A(n1618), .Y(n2200) );
  AOI22XL U697 ( .A0(n149), .A1(N858), .B0(data[0]), .B1(n169), .Y(n1618) );
  INVX1 U699 ( .A(n1522), .Y(n1868) );
  INVX1 U700 ( .A(n1523), .Y(n1879) );
  AOI22XL U701 ( .A0(n147), .A1(N816), .B0(N808), .B1(n111), .Y(n1523) );
  INVX1 U702 ( .A(n1524), .Y(n1890) );
  INVX1 U703 ( .A(n1525), .Y(n1901) );
  AOI22XL U704 ( .A0(n144), .A1(N814), .B0(N806), .B1(n113), .Y(n1525) );
  INVX1 U705 ( .A(n1526), .Y(n1912) );
  AOI22XL U706 ( .A0(n146), .A1(N813), .B0(N805), .B1(n111), .Y(n1526) );
  INVX1 U707 ( .A(n1527), .Y(n1923) );
  AOI22XL U708 ( .A0(n141), .A1(N812), .B0(N804), .B1(n112), .Y(n1527) );
  INVX1 U711 ( .A(n1528), .Y(n1934) );
  INVX1 U712 ( .A(n1529), .Y(n1945) );
  AOI22XL U713 ( .A0(n144), .A1(N810), .B0(N802), .B1(n112), .Y(n1529) );
  INVX1 U715 ( .A(n1530), .Y(n1956) );
  AOI22XL U717 ( .A0(n146), .A1(N809), .B0(N801), .B1(n111), .Y(n1530) );
  INVX1 U718 ( .A(n1531), .Y(n1967) );
  AOI22XL U720 ( .A0(n147), .A1(N808), .B0(N800), .B1(n113), .Y(n1531) );
  INVX1 U721 ( .A(n1532), .Y(n1978) );
  AOI22XL U723 ( .A0(n142), .A1(N807), .B0(N799), .B1(n111), .Y(n1532) );
  INVX1 U724 ( .A(n1533), .Y(n1989) );
  INVX1 U725 ( .A(n1534), .Y(n2000) );
  AOI22XL U726 ( .A0(n144), .A1(N805), .B0(N797), .B1(n111), .Y(n1534) );
  INVX1 U727 ( .A(n1535), .Y(n2011) );
  AOI22XL U728 ( .A0(n141), .A1(N804), .B0(N796), .B1(n111), .Y(n1535) );
  INVX1 U729 ( .A(n1536), .Y(n2022) );
  INVX1 U730 ( .A(n1537), .Y(n2033) );
  AOI22XL U731 ( .A0(n146), .A1(N802), .B0(N794), .B1(n111), .Y(n1537) );
  AOI22XL U732 ( .A0(n141), .A1(N801), .B0(data[7]), .B1(n113), .Y(n1538) );
  INVX1 U733 ( .A(n1539), .Y(n1813) );
  AOI22XL U734 ( .A0(n144), .A1(N800), .B0(data[6]), .B1(n113), .Y(n1539) );
  INVX1 U735 ( .A(n1540), .Y(n1814) );
  AOI22XL U736 ( .A0(n142), .A1(N799), .B0(data[5]), .B1(n111), .Y(n1540) );
  INVX1 U737 ( .A(n1542), .Y(n1815) );
  INVX1 U738 ( .A(n1543), .Y(n1824) );
  AOI22XL U739 ( .A0(n147), .A1(N796), .B0(data[2]), .B1(n113), .Y(n1543) );
  INVX1 U740 ( .A(n1544), .Y(n1825) );
  AOI22XL U741 ( .A0(n142), .A1(N795), .B0(data[1]), .B1(n112), .Y(n1544) );
  INVX1 U742 ( .A(n1545), .Y(n2202) );
  AOI22XL U743 ( .A0(n141), .A1(N794), .B0(data[0]), .B1(n111), .Y(n1545) );
  INVX1 U744 ( .A(n1452), .Y(n1473) );
  INVX1 U745 ( .A(n1453), .Y(n1474) );
  AOI22XL U746 ( .A0(n694), .A1(N752), .B0(N744), .B1(n690), .Y(n1453) );
  INVX1 U747 ( .A(n1454), .Y(n1478) );
  AOI22XL U748 ( .A0(n693), .A1(N751), .B0(N743), .B1(n690), .Y(n1454) );
  INVX1 U749 ( .A(n1455), .Y(n1541) );
  AOI22XL U750 ( .A0(n694), .A1(N750), .B0(N742), .B1(n690), .Y(n1455) );
  INVX1 U751 ( .A(n1456), .Y(n1625) );
  AOI22XL U752 ( .A0(n694), .A1(N749), .B0(N741), .B1(n690), .Y(n1456) );
  INVX1 U753 ( .A(n1457), .Y(n1626) );
  AOI22XL U754 ( .A0(n693), .A1(N748), .B0(N740), .B1(n690), .Y(n1457) );
  INVX1 U755 ( .A(n1458), .Y(n1627) );
  AOI22XL U756 ( .A0(n694), .A1(N747), .B0(N739), .B1(n690), .Y(n1458) );
  INVX1 U757 ( .A(n1459), .Y(n1639) );
  INVX1 U758 ( .A(n1460), .Y(n1656) );
  AOI22XL U759 ( .A0(n693), .A1(N745), .B0(N737), .B1(n690), .Y(n1460) );
  INVX1 U760 ( .A(n1461), .Y(n1660) );
  AOI22XL U761 ( .A0(n694), .A1(N744), .B0(N736), .B1(n690), .Y(n1461) );
  INVX1 U762 ( .A(n1462), .Y(n1661) );
  AOI22XL U763 ( .A0(n693), .A1(N743), .B0(N735), .B1(n690), .Y(n1462) );
  INVX1 U764 ( .A(n1463), .Y(n1663) );
  AOI22XL U765 ( .A0(n694), .A1(N742), .B0(N734), .B1(n690), .Y(n1463) );
  INVX1 U766 ( .A(n1464), .Y(n1669) );
  INVX1 U767 ( .A(n1465), .Y(n1672) );
  AOI22XL U768 ( .A0(n693), .A1(N740), .B0(N732), .B1(n691), .Y(n1465) );
  INVX1 U769 ( .A(n1466), .Y(n1673) );
  AOI22XL U770 ( .A0(n694), .A1(N739), .B0(N731), .B1(n691), .Y(n1466) );
  INVX1 U771 ( .A(n1467), .Y(n1681) );
  AOI22XL U772 ( .A0(n694), .A1(N738), .B0(N730), .B1(n690), .Y(n1467) );
  INVX1 U773 ( .A(n1468), .Y(n1109) );
  AOI22XL U774 ( .A0(n693), .A1(N737), .B0(data[7]), .B1(n691), .Y(n1468) );
  INVX1 U775 ( .A(n1469), .Y(n1110) );
  AOI22XL U776 ( .A0(n694), .A1(N736), .B0(data[6]), .B1(n690), .Y(n1469) );
  INVX1 U777 ( .A(n1470), .Y(n1111) );
  AOI22XL U778 ( .A0(n693), .A1(N735), .B0(data[5]), .B1(n691), .Y(n1470) );
  INVX1 U779 ( .A(n1471), .Y(n1112) );
  AOI22XL U780 ( .A0(n694), .A1(N734), .B0(data[4]), .B1(n1444), .Y(n1471) );
  INVX1 U781 ( .A(n1472), .Y(n1113) );
  AOI22XL U782 ( .A0(n693), .A1(N733), .B0(data[3]), .B1(n691), .Y(n1472) );
  AOI22XL U783 ( .A0(n694), .A1(N730), .B0(data[0]), .B1(n1444), .Y(n1475) );
  INVX1 U784 ( .A(n1381), .Y(n1066) );
  INVX1 U785 ( .A(n1382), .Y(n1067) );
  INVX1 U786 ( .A(n1383), .Y(n1068) );
  INVX1 U787 ( .A(n1384), .Y(n1069) );
  INVX1 U788 ( .A(n1385), .Y(n1070) );
  INVX1 U789 ( .A(n1386), .Y(n1071) );
  INVX1 U790 ( .A(n1387), .Y(n1072) );
  INVX1 U791 ( .A(n1388), .Y(n1073) );
  INVX1 U792 ( .A(n1389), .Y(n1074) );
  INVX1 U793 ( .A(n1390), .Y(n1075) );
  INVX1 U794 ( .A(n1391), .Y(n1076) );
  AOI22XL U795 ( .A0(n707), .A1(N679), .B0(N671), .B1(n704), .Y(n1391) );
  INVX1 U796 ( .A(n1392), .Y(n1077) );
  AOI22XL U797 ( .A0(n707), .A1(N678), .B0(N670), .B1(n704), .Y(n1392) );
  INVX1 U798 ( .A(n1393), .Y(n1078) );
  INVX1 U799 ( .A(n1394), .Y(n1079) );
  AOI22XL U800 ( .A0(n707), .A1(N676), .B0(N668), .B1(n703), .Y(n1394) );
  INVX1 U801 ( .A(n1395), .Y(n1080) );
  AOI22XL U802 ( .A0(n707), .A1(N675), .B0(N667), .B1(n703), .Y(n1395) );
  INVX1 U803 ( .A(n1396), .Y(n1081) );
  AOI22XL U804 ( .A0(n707), .A1(N674), .B0(N666), .B1(n703), .Y(n1396) );
  INVX1 U805 ( .A(n1397), .Y(n1042) );
  AOI22XL U806 ( .A0(n708), .A1(N673), .B0(data[7]), .B1(n703), .Y(n1397) );
  INVX1 U807 ( .A(n1398), .Y(n1043) );
  AOI22XL U808 ( .A0(n708), .A1(N672), .B0(data[6]), .B1(n703), .Y(n1398) );
  INVX1 U809 ( .A(n1399), .Y(n1044) );
  AOI22XL U810 ( .A0(n708), .A1(N671), .B0(data[5]), .B1(n703), .Y(n1399) );
  INVX1 U811 ( .A(n1400), .Y(n1045) );
  AOI22XL U812 ( .A0(n708), .A1(N670), .B0(data[4]), .B1(n703), .Y(n1400) );
  INVX1 U813 ( .A(n1401), .Y(n1046) );
  AOI22XL U814 ( .A0(n708), .A1(N669), .B0(data[3]), .B1(n703), .Y(n1401) );
  INVX1 U815 ( .A(n1402), .Y(n1047) );
  AOI22XL U816 ( .A0(n708), .A1(N668), .B0(data[2]), .B1(n703), .Y(n1402) );
  INVX1 U817 ( .A(n1403), .Y(n1048) );
  AOI22XL U818 ( .A0(n708), .A1(N667), .B0(data[1]), .B1(n703), .Y(n1403) );
  INVX1 U819 ( .A(n1404), .Y(n2206) );
  AOI22XL U820 ( .A0(n708), .A1(N666), .B0(data[0]), .B1(n703), .Y(n1404) );
  INVX1 U821 ( .A(n1309), .Y(n995) );
  INVX1 U822 ( .A(n1310), .Y(n996) );
  INVX1 U823 ( .A(n1311), .Y(n997) );
  AOI22XL U824 ( .A0(n718), .A1(N623), .B0(N615), .B1(n161), .Y(n1311) );
  INVX1 U825 ( .A(n1312), .Y(n998) );
  AOI22XL U826 ( .A0(n718), .A1(N622), .B0(N614), .B1(n162), .Y(n1312) );
  INVX1 U827 ( .A(n1313), .Y(n999) );
  AOI22XL U828 ( .A0(n718), .A1(N621), .B0(N613), .B1(n159), .Y(n1313) );
  INVX1 U829 ( .A(n1314), .Y(n1000) );
  AOI22XL U830 ( .A0(n718), .A1(N620), .B0(N612), .B1(n160), .Y(n1314) );
  INVX1 U831 ( .A(n1315), .Y(n1001) );
  AOI22XL U832 ( .A0(n718), .A1(N619), .B0(N611), .B1(n159), .Y(n1315) );
  INVX1 U833 ( .A(n1316), .Y(n1002) );
  AOI22XL U834 ( .A0(n718), .A1(N618), .B0(N610), .B1(n160), .Y(n1316) );
  INVX1 U835 ( .A(n1317), .Y(n1003) );
  AOI22XL U836 ( .A0(n718), .A1(N617), .B0(N609), .B1(n162), .Y(n1317) );
  INVX1 U837 ( .A(n1318), .Y(n1004) );
  AOI22XL U838 ( .A0(n718), .A1(N616), .B0(N608), .B1(n161), .Y(n1318) );
  INVX1 U839 ( .A(n1319), .Y(n1005) );
  AOI22XL U840 ( .A0(n718), .A1(N615), .B0(N607), .B1(n161), .Y(n1319) );
  INVX1 U841 ( .A(n1320), .Y(n1006) );
  AOI22XL U842 ( .A0(n718), .A1(N614), .B0(N606), .B1(n162), .Y(n1320) );
  INVX1 U843 ( .A(n1321), .Y(n1007) );
  INVX1 U844 ( .A(n1322), .Y(n1008) );
  AOI22XL U845 ( .A0(n718), .A1(N612), .B0(N604), .B1(n160), .Y(n1322) );
  INVX1 U846 ( .A(n1323), .Y(n1009) );
  AOI22XL U847 ( .A0(n718), .A1(N611), .B0(N603), .B1(n161), .Y(n1323) );
  INVX1 U848 ( .A(n1324), .Y(n1010) );
  AOI22XL U849 ( .A0(n718), .A1(N610), .B0(N602), .B1(n162), .Y(n1324) );
  INVX1 U850 ( .A(n1325), .Y(n980) );
  AOI22XL U851 ( .A0(n718), .A1(N609), .B0(data[7]), .B1(n156), .Y(n1325) );
  INVX1 U852 ( .A(n1326), .Y(n981) );
  AOI22XL U853 ( .A0(n718), .A1(N608), .B0(data[6]), .B1(n159), .Y(n1326) );
  INVX1 U854 ( .A(n1327), .Y(n982) );
  AOI22XL U855 ( .A0(n718), .A1(N607), .B0(data[5]), .B1(n156), .Y(n1327) );
  INVX1 U856 ( .A(n1328), .Y(n983) );
  AOI22XL U857 ( .A0(n718), .A1(N606), .B0(data[4]), .B1(n159), .Y(n1328) );
  INVX1 U858 ( .A(n1329), .Y(n984) );
  AOI22XL U859 ( .A0(n718), .A1(N605), .B0(data[3]), .B1(n159), .Y(n1329) );
  INVX1 U860 ( .A(n1330), .Y(n985) );
  AOI22XL U861 ( .A0(n718), .A1(N604), .B0(data[2]), .B1(n156), .Y(n1330) );
  INVX1 U862 ( .A(n1331), .Y(n986) );
  AOI22XL U863 ( .A0(n718), .A1(N603), .B0(data[1]), .B1(n159), .Y(n1331) );
  INVX1 U864 ( .A(n1332), .Y(n2208) );
  AOI22XL U865 ( .A0(n718), .A1(N602), .B0(data[0]), .B1(n160), .Y(n1332) );
  INVX1 U866 ( .A(n1167), .Y(n871) );
  AOI22X1 U867 ( .A0(n733), .A1(N497), .B0(N489), .B1(n731), .Y(n1167) );
  INVX1 U868 ( .A(n1168), .Y(n872) );
  AOI22X1 U869 ( .A0(n733), .A1(N496), .B0(N488), .B1(n731), .Y(n1168) );
  INVX1 U870 ( .A(n1169), .Y(n873) );
  AOI22X1 U871 ( .A0(n733), .A1(N495), .B0(N487), .B1(n731), .Y(n1169) );
  INVX1 U872 ( .A(n1170), .Y(n874) );
  AOI22X1 U873 ( .A0(n733), .A1(N494), .B0(N486), .B1(n731), .Y(n1170) );
  INVX1 U874 ( .A(n1171), .Y(n875) );
  AOI22X1 U875 ( .A0(n733), .A1(N493), .B0(N485), .B1(n731), .Y(n1171) );
  INVX1 U876 ( .A(n1172), .Y(n876) );
  AOI22X1 U877 ( .A0(n733), .A1(N492), .B0(N484), .B1(n731), .Y(n1172) );
  INVX1 U878 ( .A(n1173), .Y(n877) );
  AOI22X1 U879 ( .A0(n733), .A1(N491), .B0(N483), .B1(n731), .Y(n1173) );
  INVX1 U880 ( .A(n1174), .Y(n878) );
  AOI22X1 U881 ( .A0(n733), .A1(N490), .B0(N482), .B1(n731), .Y(n1174) );
  INVX1 U882 ( .A(n1175), .Y(n879) );
  AOI22X1 U883 ( .A0(n733), .A1(N489), .B0(N481), .B1(n731), .Y(n1175) );
  INVX1 U884 ( .A(n1176), .Y(n880) );
  AOI22X1 U885 ( .A0(n733), .A1(N488), .B0(N480), .B1(n731), .Y(n1176) );
  INVX1 U886 ( .A(n1177), .Y(n881) );
  AOI22X1 U887 ( .A0(n733), .A1(N487), .B0(N479), .B1(n731), .Y(n1177) );
  INVX1 U888 ( .A(n1178), .Y(n882) );
  AOI22X1 U889 ( .A0(n733), .A1(N486), .B0(N478), .B1(n731), .Y(n1178) );
  INVX1 U890 ( .A(n1179), .Y(n883) );
  INVX1 U891 ( .A(n1180), .Y(n884) );
  AOI22X1 U892 ( .A0(n733), .A1(N484), .B0(N476), .B1(n732), .Y(n1180) );
  INVX1 U893 ( .A(n1181), .Y(n885) );
  AOI22X1 U894 ( .A0(n733), .A1(N483), .B0(N475), .B1(n732), .Y(n1181) );
  INVX1 U895 ( .A(n1182), .Y(n886) );
  AOI22X1 U896 ( .A0(n733), .A1(N482), .B0(N474), .B1(n732), .Y(n1182) );
  INVX1 U897 ( .A(n1183), .Y(n856) );
  INVX1 U898 ( .A(n1184), .Y(n857) );
  INVX1 U899 ( .A(n1185), .Y(n858) );
  INVX1 U900 ( .A(n1186), .Y(n859) );
  INVX1 U901 ( .A(n1187), .Y(n860) );
  INVX1 U902 ( .A(n1188), .Y(n861) );
  INVX1 U903 ( .A(n1189), .Y(n862) );
  INVX1 U904 ( .A(n1697), .Y(n2197) );
  INVX1 U905 ( .A(n1236), .Y(n933) );
  AOI22X1 U906 ( .A0(n725), .A1(N561), .B0(N553), .B1(n723), .Y(n1236) );
  INVX1 U907 ( .A(n1237), .Y(n934) );
  AOI22X1 U908 ( .A0(n725), .A1(N560), .B0(N552), .B1(n723), .Y(n1237) );
  INVX1 U909 ( .A(n1238), .Y(n935) );
  AOI22X1 U910 ( .A0(n725), .A1(N559), .B0(N551), .B1(n723), .Y(n1238) );
  INVX1 U911 ( .A(n1239), .Y(n936) );
  AOI22X1 U912 ( .A0(n725), .A1(N558), .B0(N550), .B1(n723), .Y(n1239) );
  INVX1 U913 ( .A(n1240), .Y(n937) );
  AOI22X1 U914 ( .A0(n725), .A1(N557), .B0(N549), .B1(n723), .Y(n1240) );
  INVX1 U915 ( .A(n1241), .Y(n938) );
  AOI22X1 U916 ( .A0(n725), .A1(N556), .B0(N548), .B1(n723), .Y(n1241) );
  INVX1 U917 ( .A(n1242), .Y(n939) );
  AOI22X1 U918 ( .A0(n725), .A1(N555), .B0(N547), .B1(n723), .Y(n1242) );
  INVX1 U919 ( .A(n1243), .Y(n940) );
  AOI22X1 U920 ( .A0(n725), .A1(N554), .B0(N546), .B1(n723), .Y(n1243) );
  INVX1 U921 ( .A(n1244), .Y(n941) );
  AOI22X1 U922 ( .A0(n725), .A1(N553), .B0(N545), .B1(n723), .Y(n1244) );
  INVX1 U923 ( .A(n1245), .Y(n942) );
  AOI22X1 U924 ( .A0(n725), .A1(N552), .B0(N544), .B1(n723), .Y(n1245) );
  INVX1 U925 ( .A(n1246), .Y(n943) );
  AOI22X1 U926 ( .A0(n725), .A1(N551), .B0(N543), .B1(n723), .Y(n1246) );
  INVX1 U927 ( .A(n1247), .Y(n944) );
  AOI22X1 U928 ( .A0(n725), .A1(N550), .B0(N542), .B1(n723), .Y(n1247) );
  INVX1 U929 ( .A(n1248), .Y(n945) );
  AOI22X1 U930 ( .A0(n725), .A1(N549), .B0(N541), .B1(n724), .Y(n1248) );
  INVX1 U931 ( .A(n1249), .Y(n946) );
  AOI22X1 U932 ( .A0(n725), .A1(N548), .B0(N540), .B1(n724), .Y(n1249) );
  INVX1 U933 ( .A(n1250), .Y(n947) );
  AOI22X1 U934 ( .A0(n725), .A1(N547), .B0(N539), .B1(n723), .Y(n1250) );
  INVX1 U935 ( .A(n1251), .Y(n948) );
  AOI22X1 U936 ( .A0(n725), .A1(N546), .B0(N538), .B1(n724), .Y(n1251) );
  INVX1 U937 ( .A(n1252), .Y(n918) );
  INVX1 U938 ( .A(n1253), .Y(n919) );
  INVX1 U939 ( .A(n1254), .Y(n920) );
  INVX1 U940 ( .A(n1255), .Y(n921) );
  INVX1 U941 ( .A(n1256), .Y(n922) );
  INVX1 U942 ( .A(n1257), .Y(n923) );
  INVX1 U943 ( .A(n1258), .Y(n924) );
  INVX1 U944 ( .A(n1259), .Y(n2211) );
  INVX1 U945 ( .A(n1631), .Y(n2161) );
  AOI22XL U946 ( .A0(n154), .A1(N912), .B0(N904), .B1(n75), .Y(n1631) );
  INVX1 U947 ( .A(n1633), .Y(n2163) );
  AOI22XL U948 ( .A0(n154), .A1(N910), .B0(N902), .B1(n75), .Y(n1633) );
  INVX1 U949 ( .A(n1634), .Y(n2164) );
  INVX1 U950 ( .A(n1635), .Y(n2165) );
  AOI22XL U951 ( .A0(n154), .A1(N908), .B0(N900), .B1(n75), .Y(n1635) );
  AOI22XL U952 ( .A0(n154), .A1(N906), .B0(N898), .B1(n72), .Y(n1637) );
  INVX1 U953 ( .A(n1638), .Y(n2168) );
  AOI22XL U954 ( .A0(n154), .A1(N905), .B0(N897), .B1(n72), .Y(n1638) );
  INVX1 U955 ( .A(n1640), .Y(n2169) );
  INVX1 U956 ( .A(n1641), .Y(n2170) );
  INVX1 U957 ( .A(n1642), .Y(n2171) );
  AOI22XL U958 ( .A0(n154), .A1(N901), .B0(N893), .B1(n75), .Y(n1642) );
  INVX1 U959 ( .A(n1643), .Y(n2172) );
  AOI22XL U960 ( .A0(n154), .A1(N900), .B0(N892), .B1(n75), .Y(n1643) );
  INVX1 U961 ( .A(n1644), .Y(n2173) );
  INVX1 U962 ( .A(n1645), .Y(n2174) );
  AOI22XL U963 ( .A0(n154), .A1(N897), .B0(data[7]), .B1(n75), .Y(n1646) );
  INVX1 U964 ( .A(n1647), .Y(n2149) );
  INVX1 U965 ( .A(n1648), .Y(n2150) );
  INVX1 U966 ( .A(n1649), .Y(n2151) );
  AOI22XL U967 ( .A0(n155), .A1(N893), .B0(data[3]), .B1(n75), .Y(n1650) );
  INVX1 U968 ( .A(n1651), .Y(n2153) );
  INVX1 U969 ( .A(n1652), .Y(n2154) );
  AOI22XL U970 ( .A0(n154), .A1(N891), .B0(data[1]), .B1(n72), .Y(n1652) );
  INVX1 U971 ( .A(n1653), .Y(n2199) );
  AOI22XL U972 ( .A0(n154), .A1(N890), .B0(data[0]), .B1(n75), .Y(n1653) );
  INVX1 U973 ( .A(n1559), .Y(n2101) );
  INVX1 U974 ( .A(n1560), .Y(n2102) );
  AOI22XL U975 ( .A0(n686), .A1(N848), .B0(N840), .B1(n170), .Y(n1560) );
  INVX1 U976 ( .A(n1561), .Y(n2103) );
  AOI22XL U977 ( .A0(n686), .A1(N847), .B0(N839), .B1(n170), .Y(n1561) );
  INVX1 U978 ( .A(n1562), .Y(n2104) );
  AOI22XL U979 ( .A0(n151), .A1(N846), .B0(N838), .B1(n170), .Y(n1562) );
  INVX1 U980 ( .A(n1563), .Y(n2105) );
  AOI22XL U981 ( .A0(n151), .A1(N845), .B0(N837), .B1(n170), .Y(n1563) );
  INVX1 U982 ( .A(n1564), .Y(n2106) );
  AOI22XL U983 ( .A0(n152), .A1(N844), .B0(N836), .B1(n170), .Y(n1564) );
  INVX1 U984 ( .A(n1565), .Y(n2107) );
  AOI22XL U985 ( .A0(n686), .A1(N843), .B0(N835), .B1(n170), .Y(n1565) );
  INVX1 U986 ( .A(n1566), .Y(n2108) );
  AOI22XL U987 ( .A0(n152), .A1(N842), .B0(N834), .B1(n170), .Y(n1566) );
  INVX1 U988 ( .A(n1567), .Y(n2109) );
  AOI22XL U989 ( .A0(n686), .A1(N841), .B0(N833), .B1(n170), .Y(n1567) );
  INVX1 U990 ( .A(n1568), .Y(n2110) );
  AOI22XL U991 ( .A0(n151), .A1(N840), .B0(N832), .B1(n170), .Y(n1568) );
  INVX1 U992 ( .A(n1569), .Y(n2111) );
  AOI22XL U993 ( .A0(n152), .A1(N839), .B0(N831), .B1(n170), .Y(n1569) );
  INVX1 U994 ( .A(n1570), .Y(n2112) );
  AOI22XL U995 ( .A0(n686), .A1(N838), .B0(N830), .B1(n170), .Y(n1570) );
  INVX1 U996 ( .A(n1571), .Y(n2113) );
  AOI22XL U997 ( .A0(n686), .A1(N837), .B0(N829), .B1(n170), .Y(n1571) );
  INVX1 U998 ( .A(n1572), .Y(n2114) );
  AOI22XL U999 ( .A0(n686), .A1(N836), .B0(N828), .B1(n170), .Y(n1572) );
  INVX1 U1000 ( .A(n1573), .Y(n2115) );
  AOI22XL U1001 ( .A0(n151), .A1(N835), .B0(N827), .B1(n170), .Y(n1573) );
  INVX1 U1002 ( .A(n1574), .Y(n2116) );
  AOI22XL U1003 ( .A0(n152), .A1(N834), .B0(N826), .B1(n170), .Y(n1574) );
  INVX1 U1004 ( .A(n1575), .Y(n2044) );
  AOI22XL U1005 ( .A0(n686), .A1(N833), .B0(data[7]), .B1(n170), .Y(n1575) );
  INVX1 U1006 ( .A(n1576), .Y(n2055) );
  AOI22XL U1007 ( .A0(n151), .A1(N832), .B0(data[6]), .B1(n170), .Y(n1576) );
  INVX1 U1008 ( .A(n1577), .Y(n2066) );
  AOI22XL U1009 ( .A0(n152), .A1(N831), .B0(data[5]), .B1(n170), .Y(n1577) );
  INVX1 U1010 ( .A(n1578), .Y(n2069) );
  AOI22XL U1011 ( .A0(n686), .A1(N830), .B0(data[4]), .B1(n170), .Y(n1578) );
  INVX1 U1012 ( .A(n1579), .Y(n2090) );
  AOI22XL U1013 ( .A0(n152), .A1(N829), .B0(data[3]), .B1(n170), .Y(n1579) );
  INVX1 U1014 ( .A(n1580), .Y(n2091) );
  AOI22XL U1015 ( .A0(n686), .A1(N828), .B0(data[2]), .B1(n170), .Y(n1580) );
  INVX1 U1016 ( .A(n1581), .Y(n2092) );
  AOI22XL U1017 ( .A0(n686), .A1(N827), .B0(data[1]), .B1(n170), .Y(n1581) );
  INVX1 U1018 ( .A(n1582), .Y(n2201) );
  AOI22XL U1019 ( .A0(n151), .A1(N826), .B0(data[0]), .B1(n170), .Y(n1582) );
  INVX1 U1020 ( .A(n1486), .Y(n1748) );
  INVX1 U1021 ( .A(n1487), .Y(n1749) );
  AOI22XL U1022 ( .A0(n688), .A1(N784), .B0(N776), .B1(n172), .Y(n1487) );
  INVX1 U1023 ( .A(n1488), .Y(n1758) );
  AOI22XL U1024 ( .A0(n688), .A1(N783), .B0(N775), .B1(n172), .Y(n1488) );
  INVX1 U1025 ( .A(n1489), .Y(n1759) );
  AOI22XL U1026 ( .A0(n688), .A1(N782), .B0(N774), .B1(n172), .Y(n1489) );
  INVX1 U1027 ( .A(n1490), .Y(n1760) );
  AOI22XL U1028 ( .A0(n688), .A1(N781), .B0(N773), .B1(n172), .Y(n1490) );
  INVX1 U1029 ( .A(n1491), .Y(n1769) );
  AOI22XL U1030 ( .A0(n688), .A1(N780), .B0(N772), .B1(n172), .Y(n1491) );
  INVX1 U1031 ( .A(n1492), .Y(n1770) );
  AOI22XL U1032 ( .A0(n688), .A1(N779), .B0(N771), .B1(n172), .Y(n1492) );
  INVX1 U1033 ( .A(n1493), .Y(n1771) );
  AOI22XL U1034 ( .A0(n688), .A1(N778), .B0(N770), .B1(n172), .Y(n1493) );
  INVX1 U1035 ( .A(n1494), .Y(n1780) );
  AOI22XL U1036 ( .A0(n688), .A1(N777), .B0(N769), .B1(n172), .Y(n1494) );
  INVX1 U1037 ( .A(n1495), .Y(n1781) );
  AOI22XL U1038 ( .A0(n688), .A1(N776), .B0(N768), .B1(n172), .Y(n1495) );
  INVX1 U1039 ( .A(n1496), .Y(n1782) );
  AOI22XL U1040 ( .A0(n688), .A1(N775), .B0(N767), .B1(n172), .Y(n1496) );
  INVX1 U1041 ( .A(n1497), .Y(n1791) );
  AOI22XL U1042 ( .A0(n688), .A1(N774), .B0(N766), .B1(n172), .Y(n1497) );
  INVX1 U1043 ( .A(n1498), .Y(n1792) );
  AOI22XL U1044 ( .A0(n688), .A1(N773), .B0(N765), .B1(n172), .Y(n1498) );
  INVX1 U1045 ( .A(n1499), .Y(n1793) );
  AOI22XL U1046 ( .A0(n688), .A1(N772), .B0(N764), .B1(n172), .Y(n1499) );
  INVX1 U1047 ( .A(n1500), .Y(n1802) );
  AOI22XL U1048 ( .A0(n688), .A1(N771), .B0(N763), .B1(n172), .Y(n1500) );
  INVX1 U1049 ( .A(n1501), .Y(n1803) );
  AOI22XL U1050 ( .A0(n688), .A1(N770), .B0(N762), .B1(n172), .Y(n1501) );
  INVX1 U1051 ( .A(n1502), .Y(n1682) );
  AOI22XL U1052 ( .A0(n688), .A1(N769), .B0(data[7]), .B1(n172), .Y(n1502) );
  INVX1 U1053 ( .A(n1503), .Y(n1686) );
  AOI22XL U1054 ( .A0(n688), .A1(N768), .B0(data[6]), .B1(n172), .Y(n1503) );
  INVX1 U1055 ( .A(n1504), .Y(n1707) );
  AOI22XL U1056 ( .A0(n688), .A1(N767), .B0(data[5]), .B1(n172), .Y(n1504) );
  INVX1 U1057 ( .A(n1505), .Y(n1708) );
  AOI22XL U1058 ( .A0(n688), .A1(N766), .B0(data[4]), .B1(n172), .Y(n1505) );
  INVX1 U1059 ( .A(n1506), .Y(n1709) );
  AOI22XL U1060 ( .A0(n688), .A1(N765), .B0(data[3]), .B1(n172), .Y(n1506) );
  INVX1 U1061 ( .A(n1507), .Y(n1710) );
  AOI22XL U1062 ( .A0(n688), .A1(N764), .B0(data[2]), .B1(n172), .Y(n1507) );
  INVX1 U1063 ( .A(n1508), .Y(n1711) );
  AOI22XL U1064 ( .A0(n688), .A1(N763), .B0(data[1]), .B1(n172), .Y(n1508) );
  INVX1 U1065 ( .A(n1509), .Y(n2203) );
  AOI22XL U1066 ( .A0(n688), .A1(N762), .B0(data[0]), .B1(n172), .Y(n1509) );
  INVX1 U1067 ( .A(n1417), .Y(n1094) );
  INVX1 U1068 ( .A(n1418), .Y(n1095) );
  AOI22XL U1069 ( .A0(n699), .A1(N720), .B0(N712), .B1(n696), .Y(n1418) );
  INVX1 U1070 ( .A(n1419), .Y(n1096) );
  AOI22XL U1071 ( .A0(n699), .A1(N719), .B0(N711), .B1(n696), .Y(n1419) );
  INVX1 U1072 ( .A(n1420), .Y(n1097) );
  AOI22XL U1073 ( .A0(n699), .A1(N718), .B0(N710), .B1(n696), .Y(n1420) );
  INVX1 U1074 ( .A(n1421), .Y(n1098) );
  AOI22XL U1075 ( .A0(n700), .A1(N717), .B0(N709), .B1(n696), .Y(n1421) );
  INVX1 U1076 ( .A(n1422), .Y(n1099) );
  AOI22XL U1077 ( .A0(n700), .A1(N716), .B0(N708), .B1(n696), .Y(n1422) );
  INVX1 U1078 ( .A(n1423), .Y(n1100) );
  AOI22XL U1079 ( .A0(n700), .A1(N715), .B0(N707), .B1(n696), .Y(n1423) );
  INVX1 U1080 ( .A(n1424), .Y(n1101) );
  INVX1 U1081 ( .A(n1425), .Y(n1102) );
  AOI22XL U1082 ( .A0(n700), .A1(N713), .B0(N705), .B1(n696), .Y(n1425) );
  INVX1 U1083 ( .A(n1426), .Y(n1103) );
  AOI22XL U1084 ( .A0(n700), .A1(N712), .B0(N704), .B1(n696), .Y(n1426) );
  INVX1 U1085 ( .A(n1427), .Y(n1104) );
  AOI22XL U1086 ( .A0(n700), .A1(N711), .B0(N703), .B1(n696), .Y(n1427) );
  INVX1 U1087 ( .A(n1428), .Y(n1105) );
  AOI22XL U1088 ( .A0(n700), .A1(N710), .B0(N702), .B1(n696), .Y(n1428) );
  INVX1 U1089 ( .A(n1429), .Y(n1106) );
  INVX1 U1090 ( .A(n1430), .Y(n1107) );
  AOI22XL U1091 ( .A0(n700), .A1(N708), .B0(N700), .B1(n697), .Y(n1430) );
  INVX1 U1092 ( .A(n1431), .Y(n1108) );
  AOI22XL U1093 ( .A0(n701), .A1(N705), .B0(data[7]), .B1(n697), .Y(n1433) );
  INVX1 U1094 ( .A(n1434), .Y(n1083) );
  INVX1 U1095 ( .A(n1435), .Y(n1084) );
  INVX1 U1096 ( .A(n1436), .Y(n1085) );
  AOI22XL U1097 ( .A0(n701), .A1(N698), .B0(data[0]), .B1(n697), .Y(n1440) );
  INVX1 U1098 ( .A(n1274), .Y(n964) );
  AOI22X1 U1099 ( .A0(n721), .A1(N593), .B0(N585), .B1(n138), .Y(n1274) );
  INVX1 U1100 ( .A(n1275), .Y(n965) );
  AOI22X1 U1101 ( .A0(n721), .A1(N592), .B0(N584), .B1(n139), .Y(n1275) );
  INVX1 U1102 ( .A(n1276), .Y(n966) );
  AOI22X1 U1103 ( .A0(n721), .A1(N591), .B0(N583), .B1(n140), .Y(n1276) );
  INVX1 U1104 ( .A(n1277), .Y(n967) );
  AOI22X1 U1107 ( .A0(n721), .A1(N590), .B0(N582), .B1(n139), .Y(n1277) );
  INVX1 U1110 ( .A(n1278), .Y(n968) );
  AOI22X1 U1111 ( .A0(n720), .A1(N589), .B0(N581), .B1(n138), .Y(n1278) );
  INVX1 U1113 ( .A(n1279), .Y(n969) );
  AOI22X1 U1115 ( .A0(n720), .A1(N588), .B0(N580), .B1(n139), .Y(n1279) );
  INVX1 U1116 ( .A(n1280), .Y(n970) );
  AOI22X1 U1117 ( .A0(n720), .A1(N587), .B0(N579), .B1(n138), .Y(n1280) );
  INVX1 U1118 ( .A(n1281), .Y(n971) );
  AOI22X1 U1119 ( .A0(n720), .A1(N586), .B0(N578), .B1(n139), .Y(n1281) );
  INVX1 U1123 ( .A(n1282), .Y(n972) );
  AOI22X1 U1127 ( .A0(n720), .A1(N585), .B0(N577), .B1(n140), .Y(n1282) );
  INVX1 U1129 ( .A(n1283), .Y(n973) );
  AOI22X1 U1130 ( .A0(n720), .A1(N584), .B0(N576), .B1(n138), .Y(n1283) );
  INVX1 U1131 ( .A(n1284), .Y(n974) );
  AOI22X1 U1133 ( .A0(n720), .A1(N583), .B0(N575), .B1(n140), .Y(n1284) );
  INVX1 U1134 ( .A(n1285), .Y(n975) );
  AOI22X1 U1135 ( .A0(n720), .A1(N582), .B0(N574), .B1(n140), .Y(n1285) );
  INVX1 U1136 ( .A(n1286), .Y(n976) );
  AOI22X1 U1137 ( .A0(n720), .A1(N581), .B0(N573), .B1(n140), .Y(n1286) );
  INVX1 U1138 ( .A(n1287), .Y(n977) );
  AOI22X1 U1139 ( .A0(n720), .A1(N580), .B0(N572), .B1(n140), .Y(n1287) );
  INVX1 U1140 ( .A(n1288), .Y(n978) );
  AOI22X1 U1141 ( .A0(n720), .A1(N579), .B0(N571), .B1(n138), .Y(n1288) );
  INVX1 U1143 ( .A(n1289), .Y(n979) );
  AOI22X1 U1144 ( .A0(n720), .A1(N578), .B0(N570), .B1(n139), .Y(n1289) );
  INVX1 U1145 ( .A(n1290), .Y(n949) );
  INVX1 U1146 ( .A(n1291), .Y(n950) );
  INVX1 U1147 ( .A(n1292), .Y(n951) );
  INVX1 U1148 ( .A(n1293), .Y(n952) );
  INVX1 U1149 ( .A(n1294), .Y(n953) );
  INVX1 U1150 ( .A(n1295), .Y(n954) );
  INVX1 U1151 ( .A(n1296), .Y(n955) );
  INVX1 U1152 ( .A(n1297), .Y(n2209) );
  INVX1 U1153 ( .A(n1345), .Y(n1026) );
  INVX1 U1154 ( .A(n1346), .Y(n1027) );
  AOI22XL U1155 ( .A0(n715), .A1(N656), .B0(N648), .B1(n711), .Y(n1346) );
  INVX1 U1156 ( .A(n1347), .Y(n1028) );
  AOI22XL U1157 ( .A0(n715), .A1(N655), .B0(N647), .B1(n711), .Y(n1347) );
  INVX1 U1158 ( .A(n1348), .Y(n1029) );
  AOI22XL U1159 ( .A0(n715), .A1(N654), .B0(N646), .B1(n711), .Y(n1348) );
  INVX1 U1160 ( .A(n1349), .Y(n1030) );
  INVX1 U1161 ( .A(n1350), .Y(n1031) );
  INVX1 U1162 ( .A(n1351), .Y(n1032) );
  INVX1 U1163 ( .A(n1352), .Y(n1033) );
  INVX1 U1164 ( .A(n1353), .Y(n1034) );
  INVX1 U1165 ( .A(n1354), .Y(n1035) );
  INVX1 U1166 ( .A(n1355), .Y(n1036) );
  AOI22XL U1167 ( .A0(n715), .A1(N647), .B0(N639), .B1(n711), .Y(n1355) );
  INVX1 U1168 ( .A(n1356), .Y(n1037) );
  AOI22XL U1169 ( .A0(n715), .A1(N646), .B0(N638), .B1(n711), .Y(n1356) );
  INVX1 U1170 ( .A(n1357), .Y(n1038) );
  INVX1 U1171 ( .A(n1358), .Y(n1039) );
  AOI22XL U1172 ( .A0(n715), .A1(N644), .B0(N636), .B1(n710), .Y(n1358) );
  INVX1 U1173 ( .A(n1359), .Y(n1040) );
  AOI22XL U1174 ( .A0(n715), .A1(N643), .B0(N635), .B1(n710), .Y(n1359) );
  INVX1 U1175 ( .A(n1360), .Y(n1041) );
  AOI22XL U1176 ( .A0(n715), .A1(N642), .B0(N634), .B1(n710), .Y(n1360) );
  INVX1 U1177 ( .A(n1361), .Y(n1011) );
  AOI22XL U1178 ( .A0(n716), .A1(N641), .B0(data[7]), .B1(n710), .Y(n1361) );
  INVX1 U1179 ( .A(n1362), .Y(n1012) );
  AOI22XL U1180 ( .A0(n716), .A1(N640), .B0(data[6]), .B1(n710), .Y(n1362) );
  INVX1 U1181 ( .A(n1363), .Y(n1013) );
  AOI22XL U1182 ( .A0(n716), .A1(N639), .B0(data[5]), .B1(n710), .Y(n1363) );
  INVX1 U1183 ( .A(n1364), .Y(n1014) );
  AOI22XL U1184 ( .A0(n716), .A1(N638), .B0(data[4]), .B1(n710), .Y(n1364) );
  INVX1 U1185 ( .A(n1365), .Y(n1015) );
  AOI22XL U1186 ( .A0(n716), .A1(N637), .B0(data[3]), .B1(n710), .Y(n1365) );
  INVX1 U1187 ( .A(n1366), .Y(n1016) );
  AOI22XL U1188 ( .A0(n716), .A1(N636), .B0(data[2]), .B1(n710), .Y(n1366) );
  INVX1 U1189 ( .A(n1367), .Y(n1017) );
  AOI22XL U1190 ( .A0(n716), .A1(N635), .B0(data[1]), .B1(n710), .Y(n1367) );
  INVX1 U1191 ( .A(n1368), .Y(n2207) );
  AOI22XL U1192 ( .A0(n716), .A1(N634), .B0(data[0]), .B1(n710), .Y(n1368) );
  INVX1 U1193 ( .A(n1200), .Y(n902) );
  AOI22X1 U1194 ( .A0(n728), .A1(N529), .B0(N521), .B1(n727), .Y(n1200) );
  INVX1 U1195 ( .A(n1201), .Y(n903) );
  AOI22X1 U1196 ( .A0(n728), .A1(N528), .B0(N520), .B1(n727), .Y(n1201) );
  INVX1 U1197 ( .A(n1202), .Y(n904) );
  AOI22X1 U1198 ( .A0(n728), .A1(N527), .B0(N519), .B1(n727), .Y(n1202) );
  INVX1 U1199 ( .A(n1203), .Y(n905) );
  AOI22X1 U1200 ( .A0(n728), .A1(N526), .B0(N518), .B1(n727), .Y(n1203) );
  INVX1 U1201 ( .A(n1204), .Y(n906) );
  AOI22X1 U1202 ( .A0(n729), .A1(N525), .B0(N517), .B1(n727), .Y(n1204) );
  INVX1 U1203 ( .A(n1205), .Y(n907) );
  AOI22X1 U1204 ( .A0(n729), .A1(N524), .B0(N516), .B1(n727), .Y(n1205) );
  INVX1 U1205 ( .A(n1206), .Y(n908) );
  AOI22X1 U1206 ( .A0(n729), .A1(N523), .B0(N515), .B1(n727), .Y(n1206) );
  INVX1 U1207 ( .A(n1207), .Y(n909) );
  AOI22X1 U1208 ( .A0(n729), .A1(N522), .B0(N514), .B1(n727), .Y(n1207) );
  INVX1 U1209 ( .A(n1208), .Y(n910) );
  AOI22X1 U1210 ( .A0(n729), .A1(N521), .B0(N513), .B1(n727), .Y(n1208) );
  INVX1 U1211 ( .A(n1209), .Y(n911) );
  AOI22X1 U1212 ( .A0(n729), .A1(N520), .B0(N512), .B1(n727), .Y(n1209) );
  INVX1 U1213 ( .A(n1210), .Y(n912) );
  AOI22X1 U1214 ( .A0(n729), .A1(N519), .B0(N511), .B1(n727), .Y(n1210) );
  INVX1 U1215 ( .A(n1211), .Y(n913) );
  AOI22X1 U1216 ( .A0(n729), .A1(N518), .B0(N510), .B1(n727), .Y(n1211) );
  INVX1 U1217 ( .A(n1212), .Y(n914) );
  INVX1 U1218 ( .A(n1213), .Y(n915) );
  AOI22X1 U1219 ( .A0(n729), .A1(N516), .B0(N508), .B1(n727), .Y(n1213) );
  INVX1 U1220 ( .A(n1214), .Y(n916) );
  AOI22X1 U1221 ( .A0(n729), .A1(N515), .B0(N507), .B1(n727), .Y(n1214) );
  INVX1 U1222 ( .A(n1215), .Y(n917) );
  AOI22X1 U1223 ( .A0(n729), .A1(N514), .B0(N506), .B1(n727), .Y(n1215) );
  INVX1 U1224 ( .A(n1216), .Y(n887) );
  INVX1 U1225 ( .A(n1217), .Y(n888) );
  INVX1 U1226 ( .A(n1218), .Y(n889) );
  INVX1 U1227 ( .A(n1219), .Y(n890) );
  INVX1 U1228 ( .A(n1220), .Y(n891) );
  INVX1 U1229 ( .A(n1221), .Y(n892) );
  INVX1 U1230 ( .A(n1222), .Y(n893) );
  INVX1 U1231 ( .A(n1223), .Y(n2212) );
  INVX1 U1232 ( .A(n1124), .Y(n840) );
  AOI22X1 U1233 ( .A0(n739), .A1(N465), .B0(N457), .B1(n1116), .Y(n1124) );
  INVX1 U1234 ( .A(n1125), .Y(n841) );
  AOI22X1 U1235 ( .A0(n739), .A1(N464), .B0(N456), .B1(n1116), .Y(n1125) );
  INVX1 U1236 ( .A(n1126), .Y(n842) );
  AOI22X1 U1237 ( .A0(n739), .A1(N463), .B0(N455), .B1(n1116), .Y(n1126) );
  INVX1 U1238 ( .A(n1127), .Y(n843) );
  AOI22X1 U1239 ( .A0(n739), .A1(N462), .B0(N454), .B1(n1116), .Y(n1127) );
  INVX1 U1240 ( .A(n1128), .Y(n844) );
  AOI22X1 U1241 ( .A0(n740), .A1(N461), .B0(N453), .B1(n736), .Y(n1128) );
  INVX1 U1242 ( .A(n1129), .Y(n845) );
  AOI22X1 U1243 ( .A0(n740), .A1(N460), .B0(N452), .B1(n736), .Y(n1129) );
  INVX1 U1244 ( .A(n1130), .Y(n846) );
  AOI22X1 U1245 ( .A0(n740), .A1(N459), .B0(N451), .B1(n736), .Y(n1130) );
  INVX1 U1246 ( .A(n1131), .Y(n847) );
  AOI22X1 U1247 ( .A0(n740), .A1(N458), .B0(N450), .B1(n736), .Y(n1131) );
  INVX1 U1248 ( .A(n1132), .Y(n848) );
  AOI22X1 U1249 ( .A0(n740), .A1(N457), .B0(N449), .B1(n736), .Y(n1132) );
  INVX1 U1250 ( .A(n1133), .Y(n849) );
  AOI22X1 U1251 ( .A0(n740), .A1(N456), .B0(N448), .B1(n735), .Y(n1133) );
  INVX1 U1252 ( .A(n1134), .Y(n850) );
  AOI22X1 U1253 ( .A0(n740), .A1(N455), .B0(N447), .B1(n1116), .Y(n1134) );
  INVX1 U1254 ( .A(n1135), .Y(n851) );
  AOI22X1 U1255 ( .A0(n740), .A1(N454), .B0(N446), .B1(n1116), .Y(n1135) );
  INVX1 U1256 ( .A(n1136), .Y(n852) );
  INVX1 U1257 ( .A(n1137), .Y(n853) );
  AOI22X1 U1258 ( .A0(n740), .A1(N452), .B0(N444), .B1(n735), .Y(n1137) );
  INVX1 U1259 ( .A(n1138), .Y(n854) );
  AOI22X1 U1260 ( .A0(n740), .A1(N451), .B0(N443), .B1(n735), .Y(n1138) );
  INVX1 U1261 ( .A(n1139), .Y(n855) );
  AOI22X1 U1262 ( .A0(n740), .A1(N450), .B0(N442), .B1(n735), .Y(n1139) );
  INVX1 U1263 ( .A(n1140), .Y(n825) );
  INVX1 U1264 ( .A(n1141), .Y(n826) );
  INVX1 U1265 ( .A(n1142), .Y(n827) );
  INVX1 U1266 ( .A(n1143), .Y(n828) );
  INVX1 U1267 ( .A(n1144), .Y(n829) );
  INVX1 U1268 ( .A(n1145), .Y(n830) );
  INVX1 U1269 ( .A(n1146), .Y(n831) );
  INVX1 U1270 ( .A(n1147), .Y(n2210) );
  INVX1 U1271 ( .A(n1659), .Y(n2180) );
  INVX1 U1272 ( .A(n1662), .Y(n2181) );
  INVX1 U1273 ( .A(n1664), .Y(n2182) );
  INVX1 U1274 ( .A(n1665), .Y(n2183) );
  AOI22XL U1275 ( .A0(n154), .A1(buffer[15]), .B0(N913), .B1(n72), .Y(n1620)
         );
  INVX1 U1276 ( .A(n1623), .Y(n2156) );
  INVX1 U1277 ( .A(n1624), .Y(n2157) );
  AOI22XL U1278 ( .A0(n154), .A1(buffer[13]), .B0(N911), .B1(n72), .Y(n1624)
         );
  INVX1 U1279 ( .A(n1629), .Y(n2159) );
  INVX1 U1280 ( .A(n1585), .Y(n2124) );
  AOI22XL U1281 ( .A0(n150), .A1(buffer[23]), .B0(N881), .B1(n169), .Y(n1585)
         );
  INVX1 U1282 ( .A(n1588), .Y(n2125) );
  AOI22XL U1283 ( .A0(n683), .A1(buffer[22]), .B0(N880), .B1(n169), .Y(n1588)
         );
  INVX1 U1284 ( .A(n1589), .Y(n2126) );
  AOI22XL U1285 ( .A0(n683), .A1(buffer[21]), .B0(N879), .B1(n169), .Y(n1589)
         );
  INVX1 U1286 ( .A(n1590), .Y(n2127) );
  AOI22XL U1287 ( .A0(n683), .A1(buffer[20]), .B0(N878), .B1(n169), .Y(n1590)
         );
  INVX1 U1288 ( .A(n1591), .Y(n2128) );
  AOI22XL U1289 ( .A0(n149), .A1(buffer[19]), .B0(N877), .B1(n169), .Y(n1591)
         );
  INVX1 U1290 ( .A(n1592), .Y(n2129) );
  AOI22XL U1291 ( .A0(n150), .A1(buffer[18]), .B0(N876), .B1(n169), .Y(n1592)
         );
  INVX1 U1292 ( .A(n1593), .Y(n2130) );
  AOI22XL U1293 ( .A0(n683), .A1(buffer[17]), .B0(N875), .B1(n169), .Y(n1593)
         );
  INVX1 U1294 ( .A(n1594), .Y(n2131) );
  AOI22XL U1295 ( .A0(n149), .A1(buffer[16]), .B0(N874), .B1(n169), .Y(n1594)
         );
  INVX1 U1296 ( .A(n1549), .Y(n2093) );
  AOI22XL U1297 ( .A0(n152), .A1(buffer[31]), .B0(N849), .B1(n170), .Y(n1549)
         );
  INVX1 U1298 ( .A(n1552), .Y(n2094) );
  AOI22XL U1299 ( .A0(n686), .A1(buffer[30]), .B0(N848), .B1(n170), .Y(n1552)
         );
  INVX1 U1300 ( .A(n1553), .Y(n2095) );
  AOI22XL U1301 ( .A0(n686), .A1(buffer[29]), .B0(N847), .B1(n170), .Y(n1553)
         );
  INVX1 U1302 ( .A(n1554), .Y(n2096) );
  AOI22XL U1303 ( .A0(n686), .A1(buffer[28]), .B0(N846), .B1(n170), .Y(n1554)
         );
  INVX1 U1304 ( .A(n1555), .Y(n2097) );
  AOI22XL U1305 ( .A0(n151), .A1(buffer[27]), .B0(N845), .B1(n170), .Y(n1555)
         );
  INVX1 U1306 ( .A(n1556), .Y(n2098) );
  AOI22XL U1307 ( .A0(n152), .A1(buffer[26]), .B0(N844), .B1(n170), .Y(n1556)
         );
  INVX1 U1308 ( .A(n1557), .Y(n2099) );
  AOI22XL U1309 ( .A0(n686), .A1(buffer[25]), .B0(N843), .B1(n170), .Y(n1557)
         );
  INVX1 U1310 ( .A(n1558), .Y(n2100) );
  AOI22XL U1311 ( .A0(n151), .A1(buffer[24]), .B0(N842), .B1(n170), .Y(n1558)
         );
  INVX1 U1312 ( .A(n1512), .Y(n1826) );
  AOI22XL U1313 ( .A0(n141), .A1(buffer[39]), .B0(N817), .B1(n113), .Y(n1512)
         );
  INVX1 U1314 ( .A(n1515), .Y(n1835) );
  AOI22XL U1315 ( .A0(n141), .A1(buffer[38]), .B0(N816), .B1(n111), .Y(n1515)
         );
  INVX1 U1316 ( .A(n1516), .Y(n1836) );
  INVX1 U1317 ( .A(n1517), .Y(n1837) );
  AOI22XL U1318 ( .A0(n141), .A1(buffer[36]), .B0(N814), .B1(n113), .Y(n1517)
         );
  INVX1 U1319 ( .A(n1518), .Y(n1846) );
  AOI22XL U1320 ( .A0(n146), .A1(buffer[35]), .B0(N813), .B1(n112), .Y(n1518)
         );
  INVX1 U1321 ( .A(n1519), .Y(n1847) );
  AOI22XL U1322 ( .A0(n147), .A1(buffer[34]), .B0(N812), .B1(n112), .Y(n1519)
         );
  INVX1 U1323 ( .A(n1520), .Y(n1848) );
  INVX1 U1324 ( .A(n1521), .Y(n1857) );
  AOI22XL U1325 ( .A0(n144), .A1(buffer[32]), .B0(N810), .B1(n113), .Y(n1521)
         );
  INVX1 U1326 ( .A(n1476), .Y(n1712) );
  AOI22XL U1327 ( .A0(n688), .A1(buffer[47]), .B0(N785), .B1(n172), .Y(n1476)
         );
  INVX1 U1328 ( .A(n1479), .Y(n1722) );
  AOI22XL U1329 ( .A0(n688), .A1(buffer[46]), .B0(N784), .B1(n172), .Y(n1479)
         );
  INVX1 U1330 ( .A(n1480), .Y(n1732) );
  AOI22XL U1331 ( .A0(n688), .A1(buffer[45]), .B0(N783), .B1(n172), .Y(n1480)
         );
  INVX1 U1332 ( .A(n1481), .Y(n1734) );
  AOI22XL U1333 ( .A0(n688), .A1(buffer[44]), .B0(N782), .B1(n172), .Y(n1481)
         );
  INVX1 U1334 ( .A(n1482), .Y(n1736) );
  AOI22XL U1335 ( .A0(n688), .A1(buffer[43]), .B0(N781), .B1(n172), .Y(n1482)
         );
  INVX1 U1336 ( .A(n1483), .Y(n1737) );
  AOI22XL U1337 ( .A0(n688), .A1(buffer[42]), .B0(N780), .B1(n172), .Y(n1483)
         );
  INVX1 U1338 ( .A(n1484), .Y(n1738) );
  AOI22XL U1339 ( .A0(n688), .A1(buffer[41]), .B0(N779), .B1(n172), .Y(n1484)
         );
  INVX1 U1340 ( .A(n1485), .Y(n1747) );
  AOI22XL U1341 ( .A0(n688), .A1(buffer[40]), .B0(N778), .B1(n172), .Y(n1485)
         );
  INVX1 U1342 ( .A(n1442), .Y(n1150) );
  INVX1 U1343 ( .A(n1445), .Y(n1159) );
  AOI22XL U1344 ( .A0(n694), .A1(buffer[54]), .B0(N752), .B1(n691), .Y(n1445)
         );
  INVX1 U1345 ( .A(n1446), .Y(n1192) );
  AOI22XL U1346 ( .A0(n693), .A1(buffer[53]), .B0(N751), .B1(n691), .Y(n1446)
         );
  INVX1 U1347 ( .A(n1447), .Y(n1228) );
  AOI22XL U1348 ( .A0(n694), .A1(buffer[52]), .B0(N750), .B1(n691), .Y(n1447)
         );
  INVX1 U1349 ( .A(n1448), .Y(n1432) );
  AOI22XL U1350 ( .A0(n693), .A1(buffer[51]), .B0(N749), .B1(n691), .Y(n1448)
         );
  INVX1 U1351 ( .A(n1449), .Y(n1437) );
  AOI22XL U1352 ( .A0(n694), .A1(buffer[50]), .B0(N748), .B1(n691), .Y(n1449)
         );
  INVX1 U1353 ( .A(n1450), .Y(n1438) );
  AOI22XL U1354 ( .A0(n693), .A1(buffer[49]), .B0(N747), .B1(n691), .Y(n1450)
         );
  INVX1 U1355 ( .A(n1451), .Y(n1439) );
  INVX1 U1356 ( .A(n1407), .Y(n1086) );
  INVX1 U1357 ( .A(n1410), .Y(n1087) );
  AOI22XL U1358 ( .A0(n699), .A1(buffer[62]), .B0(N720), .B1(n697), .Y(n1410)
         );
  INVX1 U1359 ( .A(n1411), .Y(n1088) );
  AOI22XL U1360 ( .A0(n699), .A1(buffer[61]), .B0(N719), .B1(n697), .Y(n1411)
         );
  INVX1 U1361 ( .A(n1412), .Y(n1089) );
  AOI22XL U1362 ( .A0(n699), .A1(buffer[60]), .B0(N718), .B1(n697), .Y(n1412)
         );
  INVX1 U1363 ( .A(n1413), .Y(n1090) );
  AOI22XL U1364 ( .A0(n699), .A1(buffer[59]), .B0(N717), .B1(n697), .Y(n1413)
         );
  INVX1 U1365 ( .A(n1414), .Y(n1091) );
  AOI22XL U1366 ( .A0(n699), .A1(buffer[58]), .B0(N716), .B1(n697), .Y(n1414)
         );
  INVX1 U1367 ( .A(n1415), .Y(n1092) );
  AOI22XL U1368 ( .A0(n699), .A1(buffer[57]), .B0(N715), .B1(n697), .Y(n1415)
         );
  INVX1 U1369 ( .A(n1416), .Y(n1093) );
  INVX1 U1370 ( .A(n1299), .Y(n987) );
  AOI22X1 U1371 ( .A0(n718), .A1(buffer[87]), .B0(N625), .B1(n159), .Y(n1299)
         );
  INVX1 U1372 ( .A(n1302), .Y(n988) );
  AOI22X1 U1373 ( .A0(n718), .A1(buffer[86]), .B0(N624), .B1(n160), .Y(n1302)
         );
  INVX1 U1374 ( .A(n1303), .Y(n989) );
  AOI22X1 U1375 ( .A0(n718), .A1(buffer[85]), .B0(N623), .B1(n162), .Y(n1303)
         );
  INVX1 U1376 ( .A(n1304), .Y(n990) );
  AOI22X1 U1377 ( .A0(n718), .A1(buffer[84]), .B0(N622), .B1(n156), .Y(n1304)
         );
  INVX1 U1378 ( .A(n1305), .Y(n991) );
  AOI22X1 U1379 ( .A0(n718), .A1(buffer[83]), .B0(N621), .B1(n160), .Y(n1305)
         );
  INVX1 U1380 ( .A(n1306), .Y(n992) );
  AOI22X1 U1381 ( .A0(n718), .A1(buffer[82]), .B0(N620), .B1(n161), .Y(n1306)
         );
  INVX1 U1382 ( .A(n1307), .Y(n993) );
  AOI22X1 U1383 ( .A0(n718), .A1(buffer[81]), .B0(N619), .B1(n161), .Y(n1307)
         );
  INVX1 U1384 ( .A(n1308), .Y(n994) );
  AOI22X1 U1385 ( .A0(n718), .A1(buffer[80]), .B0(N618), .B1(n162), .Y(n1308)
         );
  INVX1 U1386 ( .A(n1264), .Y(n956) );
  AOI22X1 U1387 ( .A0(n721), .A1(buffer[95]), .B0(N593), .B1(n139), .Y(n1264)
         );
  INVX1 U1388 ( .A(n1267), .Y(n957) );
  AOI22X1 U1389 ( .A0(n721), .A1(buffer[94]), .B0(N592), .B1(n139), .Y(n1267)
         );
  INVX1 U1390 ( .A(n1268), .Y(n958) );
  AOI22X1 U1391 ( .A0(n721), .A1(buffer[93]), .B0(N591), .B1(n138), .Y(n1268)
         );
  INVX1 U1392 ( .A(n1269), .Y(n959) );
  AOI22X1 U1393 ( .A0(n721), .A1(buffer[92]), .B0(N590), .B1(n139), .Y(n1269)
         );
  INVX1 U1394 ( .A(n1270), .Y(n960) );
  AOI22X1 U1395 ( .A0(n721), .A1(buffer[91]), .B0(N589), .B1(n139), .Y(n1270)
         );
  INVX1 U1396 ( .A(n1271), .Y(n961) );
  AOI22X1 U1397 ( .A0(n721), .A1(buffer[90]), .B0(N588), .B1(n140), .Y(n1271)
         );
  INVX1 U1398 ( .A(n1272), .Y(n962) );
  AOI22X1 U1399 ( .A0(n721), .A1(buffer[89]), .B0(N587), .B1(n138), .Y(n1272)
         );
  INVX1 U1400 ( .A(n1273), .Y(n963) );
  AOI22X1 U1401 ( .A0(n721), .A1(buffer[88]), .B0(N586), .B1(n139), .Y(n1273)
         );
  INVX1 U1402 ( .A(n1335), .Y(n1018) );
  INVX1 U1403 ( .A(n1338), .Y(n1019) );
  AOI22XL U1404 ( .A0(n715), .A1(buffer[78]), .B0(N656), .B1(n712), .Y(n1338)
         );
  INVX1 U1405 ( .A(n1339), .Y(n1020) );
  AOI22XL U1406 ( .A0(n715), .A1(buffer[77]), .B0(N655), .B1(n712), .Y(n1339)
         );
  INVX1 U1407 ( .A(n1340), .Y(n1021) );
  AOI22XL U1408 ( .A0(n715), .A1(buffer[76]), .B0(N654), .B1(n712), .Y(n1340)
         );
  INVX1 U1409 ( .A(n1341), .Y(n1022) );
  AOI22XL U1410 ( .A0(n715), .A1(buffer[75]), .B0(N653), .B1(n712), .Y(n1341)
         );
  INVX1 U1411 ( .A(n1342), .Y(n1023) );
  AOI22XL U1412 ( .A0(n715), .A1(buffer[74]), .B0(N652), .B1(n712), .Y(n1342)
         );
  INVX1 U1413 ( .A(n1343), .Y(n1024) );
  AOI22XL U1414 ( .A0(n715), .A1(buffer[73]), .B0(N651), .B1(n712), .Y(n1343)
         );
  INVX1 U1415 ( .A(n1344), .Y(n1025) );
  AOI22XL U1416 ( .A0(n715), .A1(buffer[72]), .B0(N650), .B1(n712), .Y(n1344)
         );
  INVX1 U1417 ( .A(n1371), .Y(n1049) );
  INVX1 U1418 ( .A(n1374), .Y(n1050) );
  AOI22XL U1419 ( .A0(n707), .A1(buffer[70]), .B0(N688), .B1(n703), .Y(n1374)
         );
  INVX1 U1420 ( .A(n1375), .Y(n1051) );
  AOI22XL U1421 ( .A0(n707), .A1(buffer[69]), .B0(N687), .B1(n704), .Y(n1375)
         );
  INVX1 U1422 ( .A(n1376), .Y(n1052) );
  AOI22XL U1423 ( .A0(n707), .A1(buffer[68]), .B0(N686), .B1(n703), .Y(n1376)
         );
  INVX1 U1424 ( .A(n1377), .Y(n1053) );
  AOI22XL U1425 ( .A0(n707), .A1(buffer[67]), .B0(N685), .B1(n704), .Y(n1377)
         );
  INVX1 U1426 ( .A(n1378), .Y(n1063) );
  AOI22XL U1427 ( .A0(n707), .A1(buffer[66]), .B0(N684), .B1(n703), .Y(n1378)
         );
  INVX1 U1428 ( .A(n1379), .Y(n1064) );
  AOI22XL U1429 ( .A0(n707), .A1(buffer[65]), .B0(N683), .B1(n1373), .Y(n1379)
         );
  INVX1 U1430 ( .A(n1380), .Y(n1065) );
  AOI22XL U1431 ( .A0(n707), .A1(buffer[64]), .B0(N682), .B1(n1373), .Y(n1380)
         );
  INVX1 U1432 ( .A(n1157), .Y(n863) );
  AOI22X1 U1433 ( .A0(n733), .A1(buffer[119]), .B0(N497), .B1(n732), .Y(n1157)
         );
  INVX1 U1434 ( .A(n1160), .Y(n864) );
  AOI22X1 U1435 ( .A0(n733), .A1(buffer[118]), .B0(N496), .B1(n732), .Y(n1160)
         );
  INVX1 U1436 ( .A(n1161), .Y(n865) );
  AOI22X1 U1437 ( .A0(n733), .A1(buffer[117]), .B0(N495), .B1(n732), .Y(n1161)
         );
  INVX1 U1438 ( .A(n1162), .Y(n866) );
  AOI22X1 U1439 ( .A0(n733), .A1(buffer[116]), .B0(N494), .B1(n732), .Y(n1162)
         );
  INVX1 U1440 ( .A(n1163), .Y(n867) );
  AOI22X1 U1441 ( .A0(n733), .A1(buffer[115]), .B0(N493), .B1(n732), .Y(n1163)
         );
  INVX1 U1442 ( .A(n1164), .Y(n868) );
  AOI22X1 U1443 ( .A0(n733), .A1(buffer[114]), .B0(N492), .B1(n732), .Y(n1164)
         );
  INVX1 U1444 ( .A(n1165), .Y(n869) );
  AOI22X1 U1445 ( .A0(n733), .A1(buffer[113]), .B0(N491), .B1(n732), .Y(n1165)
         );
  INVX1 U1446 ( .A(n1166), .Y(n870) );
  INVX1 U1447 ( .A(n1226), .Y(n925) );
  AOI22X1 U1448 ( .A0(n725), .A1(buffer[103]), .B0(N561), .B1(n724), .Y(n1226)
         );
  INVX1 U1449 ( .A(n1229), .Y(n926) );
  AOI22X1 U1450 ( .A0(n725), .A1(buffer[102]), .B0(N560), .B1(n724), .Y(n1229)
         );
  INVX1 U1451 ( .A(n1230), .Y(n927) );
  AOI22X1 U1452 ( .A0(n725), .A1(buffer[101]), .B0(N559), .B1(n724), .Y(n1230)
         );
  INVX1 U1453 ( .A(n1231), .Y(n928) );
  AOI22X1 U1454 ( .A0(n725), .A1(buffer[100]), .B0(N558), .B1(n724), .Y(n1231)
         );
  INVX1 U1455 ( .A(n1232), .Y(n929) );
  AOI22X1 U1456 ( .A0(n725), .A1(buffer[99]), .B0(N557), .B1(n724), .Y(n1232)
         );
  INVX1 U1457 ( .A(n1233), .Y(n930) );
  AOI22X1 U1458 ( .A0(n725), .A1(buffer[98]), .B0(N556), .B1(n724), .Y(n1233)
         );
  INVX1 U1459 ( .A(n1234), .Y(n931) );
  AOI22X1 U1460 ( .A0(n725), .A1(buffer[97]), .B0(N555), .B1(n724), .Y(n1234)
         );
  INVX1 U1461 ( .A(n1235), .Y(n932) );
  INVX1 U1462 ( .A(n1190), .Y(n894) );
  AOI22X1 U1463 ( .A0(n728), .A1(buffer[111]), .B0(N529), .B1(n727), .Y(n1190)
         );
  INVX1 U1464 ( .A(n1193), .Y(n895) );
  AOI22X1 U1465 ( .A0(n728), .A1(buffer[110]), .B0(N528), .B1(n727), .Y(n1193)
         );
  INVX1 U1466 ( .A(n1194), .Y(n896) );
  AOI22X1 U1467 ( .A0(n728), .A1(buffer[109]), .B0(N527), .B1(n727), .Y(n1194)
         );
  INVX1 U1468 ( .A(n1195), .Y(n897) );
  AOI22X1 U1469 ( .A0(n728), .A1(buffer[108]), .B0(N526), .B1(n727), .Y(n1195)
         );
  INVX1 U1470 ( .A(n1196), .Y(n898) );
  AOI22X1 U1471 ( .A0(n728), .A1(buffer[107]), .B0(N525), .B1(n727), .Y(n1196)
         );
  INVX1 U1472 ( .A(n1197), .Y(n899) );
  AOI22X1 U1473 ( .A0(n728), .A1(buffer[106]), .B0(N524), .B1(n727), .Y(n1197)
         );
  INVX1 U1474 ( .A(n1198), .Y(n900) );
  AOI22X1 U1475 ( .A0(n728), .A1(buffer[105]), .B0(N523), .B1(n727), .Y(n1198)
         );
  INVX1 U1476 ( .A(n1199), .Y(n901) );
  INVX1 U1477 ( .A(n1114), .Y(n832) );
  AOI22X1 U1478 ( .A0(n739), .A1(buffer[127]), .B0(N465), .B1(n736), .Y(n1114)
         );
  INVX1 U1479 ( .A(n1117), .Y(n833) );
  AOI22X1 U1480 ( .A0(n739), .A1(buffer[126]), .B0(N464), .B1(n736), .Y(n1117)
         );
  INVX1 U1481 ( .A(n1118), .Y(n834) );
  AOI22X1 U1482 ( .A0(n739), .A1(buffer[125]), .B0(N463), .B1(n736), .Y(n1118)
         );
  INVX1 U1483 ( .A(n1119), .Y(n835) );
  AOI22X1 U1484 ( .A0(n739), .A1(buffer[124]), .B0(N462), .B1(n736), .Y(n1119)
         );
  INVX1 U1485 ( .A(n1120), .Y(n836) );
  AOI22X1 U1486 ( .A0(n739), .A1(buffer[123]), .B0(N461), .B1(n736), .Y(n1120)
         );
  INVX1 U1487 ( .A(n1121), .Y(n837) );
  AOI22X1 U1488 ( .A0(n739), .A1(buffer[122]), .B0(N460), .B1(n736), .Y(n1121)
         );
  INVX1 U1489 ( .A(n1122), .Y(n838) );
  AOI22X1 U1490 ( .A0(n739), .A1(buffer[121]), .B0(N459), .B1(n736), .Y(n1122)
         );
  INVX1 U1491 ( .A(n1123), .Y(n839) );
  XOR3X2 U1492 ( .A(R14[25]), .B(R14[29]), .C(R14[8]), .Y(sigma0[22]) );
  XOR3X2 U1493 ( .A(R14[24]), .B(R14[28]), .C(R14[7]), .Y(sigma0[21]) );
  XOR3X2 U1494 ( .A(R14[20]), .B(R14[24]), .C(R14[3]), .Y(sigma0[17]) );
  XOR3X2 U1495 ( .A(R14[19]), .B(R14[23]), .C(R14[2]), .Y(sigma0[16]) );
  XOR3X2 U1496 ( .A(R14[21]), .B(R14[25]), .C(R14[4]), .Y(sigma0[18]) );
  XOR3X2 U1497 ( .A(R14[22]), .B(R14[26]), .C(R14[5]), .Y(sigma0[19]) );
  XOR3X2 U1498 ( .A(R14[23]), .B(R14[27]), .C(R14[6]), .Y(sigma0[20]) );
  XOR3X2 U1499 ( .A(R1[30]), .B(R1[7]), .C(R1[5]), .Y(sigma1[20]) );
  XOR3X2 U1500 ( .A(R1[31]), .B(R1[8]), .C(R1[6]), .Y(sigma1[21]) );
  XOR3X2 U1501 ( .A(R1[27]), .B(R1[4]), .C(R1[2]), .Y(sigma1[17]) );
  XOR3X2 U1502 ( .A(R1[26]), .B(R1[3]), .C(R1[1]), .Y(sigma1[16]) );
  XOR3X2 U1503 ( .A(R1[28]), .B(R1[5]), .C(R1[3]), .Y(sigma1[18]) );
  XOR3X2 U1504 ( .A(R1[29]), .B(R1[6]), .C(R1[4]), .Y(sigma1[19]) );
  NAND4X1 U1505 ( .A(n1058), .B(n1057), .C(n1059), .D(n2088), .Y(n2087) );
  AOI211X1 U1506 ( .A0(counter2[0]), .A1(counter2[1]), .B0(n1056), .C0(
        counter2[2]), .Y(n2088) );
  XOR3X2 U1507 ( .A(R14[26]), .B(R14[30]), .C(R14[9]), .Y(sigma0[23]) );
  XOR3X2 U1508 ( .A(R14[12]), .B(R14[29]), .C(R14[1]), .Y(sigma0[26]) );
  XOR3X2 U1509 ( .A(R14[27]), .B(R14[31]), .C(R14[10]), .Y(sigma0[24]) );
  XOR3X2 U1510 ( .A(R14[11]), .B(R14[28]), .C(R14[0]), .Y(sigma0[25]) );
  XOR2X1 U1511 ( .A(R1[7]), .B(R1[9]), .Y(sigma1[22]) );
  NAND4X1 U1512 ( .A(counter2[6]), .B(n673), .C(n1058), .D(n1057), .Y(n1706)
         );
  XOR3X2 U1513 ( .A(R14[13]), .B(R14[30]), .C(R14[2]), .Y(sigma0[27]) );
  XOR3X2 U1514 ( .A(R14[14]), .B(R14[31]), .C(R14[3]), .Y(sigma0[28]) );
  XOR2X1 U1515 ( .A(R1[11]), .B(R1[13]), .Y(sigma1[26]) );
  NOR2X1 U1516 ( .A(counter2[2]), .B(counter2[1]), .Y(n2080) );
  NOR2X1 U1517 ( .A(n1060), .B(counter2[2]), .Y(n2079) );
  NOR2X1 U1518 ( .A(counter2[3]), .B(counter2[0]), .Y(n2076) );
  NOR2X1 U1519 ( .A(n1059), .B(counter2[0]), .Y(n2085) );
  NOR2X1 U1520 ( .A(n1061), .B(counter2[3]), .Y(n2077) );
  NOR2X1 U1521 ( .A(n1059), .B(n1061), .Y(n2086) );
  NAND4X1 U1522 ( .A(n1952), .B(n1953), .C(n1954), .D(n1955), .Y(n1946) );
  AOI22X1 U1523 ( .A0(n667), .A1(N741), .B0(n1735), .B1(N709), .Y(n1952) );
  AOI22X1 U1524 ( .A0(n669), .A1(N805), .B0(n1733), .B1(N773), .Y(n1953) );
  AOI22X1 U1525 ( .A0(n1730), .A1(N869), .B0(n1731), .B1(N837), .Y(n1954) );
  NAND4X1 U1526 ( .A(n1930), .B(n1931), .C(n1932), .D(n1933), .Y(n1924) );
  AOI22X1 U1527 ( .A0(n668), .A1(N743), .B0(n1735), .B1(N711), .Y(n1930) );
  AOI22X1 U1528 ( .A0(n670), .A1(N807), .B0(n1733), .B1(N775), .Y(n1931) );
  AOI22X1 U1529 ( .A0(n1730), .A1(N871), .B0(n1731), .B1(N839), .Y(n1932) );
  NAND4X1 U1530 ( .A(n1919), .B(n1920), .C(n1921), .D(n1922), .Y(n1913) );
  AOI22X1 U1531 ( .A0(n668), .A1(N744), .B0(n1735), .B1(N712), .Y(n1919) );
  AOI22X1 U1532 ( .A0(n670), .A1(N808), .B0(n1733), .B1(N776), .Y(n1920) );
  AOI22X1 U1533 ( .A0(n1730), .A1(N872), .B0(n1731), .B1(N840), .Y(n1921) );
  NAND4X1 U1534 ( .A(n1908), .B(n1909), .C(n1910), .D(n1911), .Y(n1902) );
  AOI22X1 U1535 ( .A0(n668), .A1(N745), .B0(n1735), .B1(N713), .Y(n1908) );
  AOI22X1 U1536 ( .A0(n670), .A1(N809), .B0(n1733), .B1(N777), .Y(n1909) );
  AOI22X1 U1537 ( .A0(n1730), .A1(N873), .B0(n1731), .B1(N841), .Y(n1910) );
  NAND4X1 U1538 ( .A(n1897), .B(n1898), .C(n1899), .D(n1900), .Y(n1891) );
  AOI22X1 U1539 ( .A0(n668), .A1(N746), .B0(n1735), .B1(N714), .Y(n1897) );
  AOI22X1 U1540 ( .A0(n670), .A1(N810), .B0(n1733), .B1(N778), .Y(n1898) );
  AOI22X1 U1541 ( .A0(n1730), .A1(N874), .B0(n1731), .B1(N842), .Y(n1899) );
  NAND4X1 U1542 ( .A(n1886), .B(n1887), .C(n1888), .D(n1889), .Y(n1880) );
  AOI22X1 U1543 ( .A0(n668), .A1(N747), .B0(n1735), .B1(N715), .Y(n1886) );
  AOI22X1 U1544 ( .A0(n670), .A1(N811), .B0(n1733), .B1(N779), .Y(n1887) );
  AOI22X1 U1545 ( .A0(n1730), .A1(N875), .B0(n1731), .B1(N843), .Y(n1888) );
  NAND4X1 U1546 ( .A(n1875), .B(n1876), .C(n1877), .D(n1878), .Y(n1869) );
  AOI22X1 U1547 ( .A0(n668), .A1(N748), .B0(n1735), .B1(N716), .Y(n1875) );
  AOI22X1 U1548 ( .A0(n670), .A1(N812), .B0(n1733), .B1(N780), .Y(n1876) );
  AOI22X1 U1549 ( .A0(n1730), .A1(N876), .B0(n1731), .B1(N844), .Y(n1877) );
  NAND4X1 U1550 ( .A(n1864), .B(n1865), .C(n1866), .D(n1867), .Y(n1858) );
  AOI22X1 U1551 ( .A0(n668), .A1(N749), .B0(n1735), .B1(N717), .Y(n1864) );
  AOI22X1 U1552 ( .A0(n670), .A1(N813), .B0(n1733), .B1(N781), .Y(n1865) );
  AOI22X1 U1553 ( .A0(n1730), .A1(N877), .B0(n1731), .B1(N845), .Y(n1866) );
  NAND4X1 U1554 ( .A(n1855), .B(n1856), .C(n1853), .D(n1854), .Y(n776) );
  AOI22X1 U1555 ( .A0(n668), .A1(N750), .B0(n1735), .B1(N718), .Y(n1853) );
  AOI22X1 U1556 ( .A0(n670), .A1(N814), .B0(n1733), .B1(N782), .Y(n1854) );
  AOI22X1 U1557 ( .A0(n1730), .A1(N878), .B0(n1731), .B1(N846), .Y(n1855) );
  NAND4X1 U1558 ( .A(n1844), .B(n1845), .C(n1842), .D(n1843), .Y(n780) );
  AOI22X1 U1559 ( .A0(n668), .A1(N751), .B0(n1735), .B1(N719), .Y(n1842) );
  AOI22X1 U1560 ( .A0(n670), .A1(N815), .B0(n1733), .B1(N783), .Y(n1843) );
  AOI22X1 U1561 ( .A0(n1730), .A1(N879), .B0(n1731), .B1(N847), .Y(n1844) );
  NAND4X1 U1562 ( .A(n1833), .B(n1834), .C(n1831), .D(n1832), .Y(n784) );
  AOI22X1 U1563 ( .A0(n668), .A1(N752), .B0(n1735), .B1(N720), .Y(n1831) );
  AOI22X1 U1564 ( .A0(n670), .A1(N816), .B0(n1733), .B1(N784), .Y(n1832) );
  AOI22X1 U1565 ( .A0(n1730), .A1(N880), .B0(n1731), .B1(N848), .Y(n1833) );
  NAND4X1 U1566 ( .A(n1822), .B(n1823), .C(n1820), .D(n1821), .Y(n788) );
  AOI22X1 U1567 ( .A0(n668), .A1(N753), .B0(n1735), .B1(N721), .Y(n1820) );
  AOI22X1 U1568 ( .A0(n670), .A1(N817), .B0(n1733), .B1(N785), .Y(n1821) );
  AOI22X1 U1569 ( .A0(n1730), .A1(N881), .B0(n1731), .B1(N849), .Y(n1822) );
  NAND4X1 U1570 ( .A(n1811), .B(n1812), .C(n1809), .D(n1810), .Y(n792) );
  AOI22X1 U1571 ( .A0(n668), .A1(buffer[48]), .B0(n1735), .B1(buffer[56]), .Y(
        n1809) );
  AOI22X1 U1572 ( .A0(n669), .A1(buffer[32]), .B0(n1733), .B1(buffer[40]), .Y(
        n1810) );
  AOI22X1 U1573 ( .A0(n1730), .A1(buffer[16]), .B0(n1731), .B1(buffer[24]), 
        .Y(n1811) );
  NAND4X1 U1574 ( .A(n1800), .B(n1801), .C(n1798), .D(n1799), .Y(n796) );
  AOI22X1 U1575 ( .A0(n667), .A1(buffer[49]), .B0(n1735), .B1(buffer[57]), .Y(
        n1798) );
  AOI22X1 U1576 ( .A0(n670), .A1(buffer[33]), .B0(n1733), .B1(buffer[41]), .Y(
        n1799) );
  AOI22X1 U1577 ( .A0(n1730), .A1(buffer[17]), .B0(n1731), .B1(buffer[25]), 
        .Y(n1800) );
  NAND4X1 U1578 ( .A(n1789), .B(n1790), .C(n1787), .D(n1788), .Y(n800) );
  AOI22X1 U1579 ( .A0(n668), .A1(buffer[50]), .B0(n1735), .B1(buffer[58]), .Y(
        n1787) );
  AOI22X1 U1580 ( .A0(n670), .A1(buffer[34]), .B0(n1733), .B1(buffer[42]), .Y(
        n1788) );
  AOI22X1 U1581 ( .A0(n1730), .A1(buffer[18]), .B0(n1731), .B1(buffer[26]), 
        .Y(n1789) );
  NAND4X1 U1582 ( .A(n1778), .B(n1779), .C(n1776), .D(n1777), .Y(n804) );
  AOI22X1 U1583 ( .A0(n668), .A1(buffer[51]), .B0(n1735), .B1(buffer[59]), .Y(
        n1776) );
  AOI22X1 U1584 ( .A0(n670), .A1(buffer[35]), .B0(n1733), .B1(buffer[43]), .Y(
        n1777) );
  AOI22X1 U1585 ( .A0(n1730), .A1(buffer[19]), .B0(n1731), .B1(buffer[27]), 
        .Y(n1778) );
  NAND4X1 U1586 ( .A(n1767), .B(n1768), .C(n1765), .D(n1766), .Y(n808) );
  AOI22X1 U1587 ( .A0(n667), .A1(buffer[52]), .B0(n1735), .B1(buffer[60]), .Y(
        n1765) );
  AOI22X1 U1588 ( .A0(n669), .A1(buffer[36]), .B0(n1733), .B1(buffer[44]), .Y(
        n1766) );
  AOI22X1 U1589 ( .A0(n1730), .A1(buffer[20]), .B0(n1731), .B1(buffer[28]), 
        .Y(n1767) );
  NAND4X1 U1590 ( .A(n1756), .B(n1757), .C(n1754), .D(n1755), .Y(n812) );
  AOI22X1 U1591 ( .A0(n668), .A1(buffer[53]), .B0(n1735), .B1(buffer[61]), .Y(
        n1754) );
  AOI22X1 U1592 ( .A0(n669), .A1(buffer[37]), .B0(n1733), .B1(buffer[45]), .Y(
        n1755) );
  AOI22X1 U1593 ( .A0(n1730), .A1(buffer[21]), .B0(n1731), .B1(buffer[29]), 
        .Y(n1756) );
  NAND4X1 U1594 ( .A(n1745), .B(n1746), .C(n1743), .D(n1744), .Y(n816) );
  AOI22X1 U1595 ( .A0(n667), .A1(buffer[54]), .B0(n1735), .B1(buffer[62]), .Y(
        n1743) );
  AOI22X1 U1596 ( .A0(n669), .A1(buffer[38]), .B0(n1733), .B1(buffer[46]), .Y(
        n1744) );
  AOI22X1 U1597 ( .A0(n1730), .A1(buffer[22]), .B0(n1731), .B1(buffer[30]), 
        .Y(n1745) );
  NAND4X1 U1598 ( .A(n1726), .B(n1727), .C(n1724), .D(n1725), .Y(n821) );
  AOI22X1 U1599 ( .A0(n667), .A1(buffer[55]), .B0(n1735), .B1(buffer[63]), .Y(
        n1724) );
  AOI22X1 U1600 ( .A0(n670), .A1(buffer[39]), .B0(n1733), .B1(buffer[47]), .Y(
        n1725) );
  AOI22X1 U1601 ( .A0(n1730), .A1(buffer[23]), .B0(n1731), .B1(buffer[31]), 
        .Y(n1726) );
  NAND4X1 U1602 ( .A(n2081), .B(n2082), .C(n2083), .D(n2084), .Y(n2067) );
  AOI22X1 U1603 ( .A0(n667), .A1(N730), .B0(n1735), .B1(N698), .Y(n2081) );
  AOI22X1 U1604 ( .A0(n669), .A1(N794), .B0(n1733), .B1(N762), .Y(n2082) );
  AOI22X1 U1605 ( .A0(n1730), .A1(N858), .B0(n1731), .B1(N826), .Y(n2083) );
  NAND4X1 U1606 ( .A(n2062), .B(n2063), .C(n2064), .D(n2065), .Y(n2056) );
  AOI22X1 U1607 ( .A0(n667), .A1(N731), .B0(n1735), .B1(N699), .Y(n2062) );
  AOI22X1 U1608 ( .A0(n669), .A1(N795), .B0(n1733), .B1(N763), .Y(n2063) );
  AOI22X1 U1609 ( .A0(n1730), .A1(N859), .B0(n1731), .B1(N827), .Y(n2064) );
  NAND4X1 U1610 ( .A(n2051), .B(n2052), .C(n2053), .D(n2054), .Y(n2045) );
  AOI22X1 U1611 ( .A0(n667), .A1(N732), .B0(n1735), .B1(N700), .Y(n2051) );
  AOI22X1 U1612 ( .A0(n669), .A1(N796), .B0(n1733), .B1(N764), .Y(n2052) );
  AOI22X1 U1613 ( .A0(n1730), .A1(N860), .B0(n1731), .B1(N828), .Y(n2053) );
  NAND4X1 U1614 ( .A(n2040), .B(n2041), .C(n2042), .D(n2043), .Y(n2034) );
  AOI22X1 U1615 ( .A0(n667), .A1(N733), .B0(n1735), .B1(N701), .Y(n2040) );
  AOI22X1 U1616 ( .A0(n669), .A1(N797), .B0(n1733), .B1(N765), .Y(n2041) );
  AOI22X1 U1617 ( .A0(n1730), .A1(N861), .B0(n1731), .B1(N829), .Y(n2042) );
  NAND4X1 U1618 ( .A(n2029), .B(n2030), .C(n2031), .D(n2032), .Y(n2023) );
  AOI22X1 U1619 ( .A0(n667), .A1(N734), .B0(n1735), .B1(N702), .Y(n2029) );
  AOI22X1 U1620 ( .A0(n669), .A1(N798), .B0(n1733), .B1(N766), .Y(n2030) );
  AOI22X1 U1621 ( .A0(n1730), .A1(N862), .B0(n1731), .B1(N830), .Y(n2031) );
  NAND4X1 U1622 ( .A(n2018), .B(n2019), .C(n2020), .D(n2021), .Y(n2012) );
  AOI22X1 U1623 ( .A0(n667), .A1(N735), .B0(n1735), .B1(N703), .Y(n2018) );
  AOI22X1 U1624 ( .A0(n669), .A1(N799), .B0(n1733), .B1(N767), .Y(n2019) );
  AOI22X1 U1625 ( .A0(n1730), .A1(N863), .B0(n1731), .B1(N831), .Y(n2020) );
  NAND4X1 U1626 ( .A(n2007), .B(n2008), .C(n2009), .D(n2010), .Y(n2001) );
  AOI22X1 U1627 ( .A0(n667), .A1(N736), .B0(n1735), .B1(N704), .Y(n2007) );
  AOI22X1 U1628 ( .A0(n669), .A1(N800), .B0(n1733), .B1(N768), .Y(n2008) );
  AOI22X1 U1629 ( .A0(n1730), .A1(N864), .B0(n1731), .B1(N832), .Y(n2009) );
  NAND4X1 U1630 ( .A(n1996), .B(n1997), .C(n1998), .D(n1999), .Y(n1990) );
  AOI22X1 U1631 ( .A0(n667), .A1(N737), .B0(n1735), .B1(N705), .Y(n1996) );
  AOI22X1 U1632 ( .A0(n669), .A1(N801), .B0(n1733), .B1(N769), .Y(n1997) );
  AOI22X1 U1633 ( .A0(n1730), .A1(N865), .B0(n1731), .B1(N833), .Y(n1998) );
  NAND4X1 U1634 ( .A(n1985), .B(n1986), .C(n1987), .D(n1988), .Y(n1979) );
  AOI22X1 U1635 ( .A0(n667), .A1(N738), .B0(n1735), .B1(N706), .Y(n1985) );
  AOI22X1 U1636 ( .A0(n669), .A1(N802), .B0(n1733), .B1(N770), .Y(n1986) );
  AOI22X1 U1637 ( .A0(n1730), .A1(N866), .B0(n1731), .B1(N834), .Y(n1987) );
  NAND4X1 U1638 ( .A(n1974), .B(n1975), .C(n1976), .D(n1977), .Y(n1968) );
  AOI22X1 U1639 ( .A0(n667), .A1(N739), .B0(n1735), .B1(N707), .Y(n1974) );
  AOI22X1 U1640 ( .A0(n669), .A1(N803), .B0(n1733), .B1(N771), .Y(n1975) );
  AOI22X1 U1641 ( .A0(n1730), .A1(N867), .B0(n1731), .B1(N835), .Y(n1976) );
  NAND4X1 U1642 ( .A(n1963), .B(n1964), .C(n1965), .D(n1966), .Y(n1957) );
  AOI22X1 U1643 ( .A0(n667), .A1(N740), .B0(n1735), .B1(N708), .Y(n1963) );
  AOI22X1 U1644 ( .A0(n669), .A1(N804), .B0(n1733), .B1(N772), .Y(n1964) );
  AOI22X1 U1645 ( .A0(n1730), .A1(N868), .B0(n1731), .B1(N836), .Y(n1965) );
  NAND4X1 U1646 ( .A(n1941), .B(n1942), .C(n1943), .D(n1944), .Y(n1935) );
  AOI22X1 U1647 ( .A0(n668), .A1(N742), .B0(n1735), .B1(N710), .Y(n1941) );
  AOI22X1 U1648 ( .A0(n670), .A1(N806), .B0(n1733), .B1(N774), .Y(n1942) );
  AOI22X1 U1649 ( .A0(n1730), .A1(N870), .B0(n1731), .B1(N838), .Y(n1943) );
  NAND4X1 U1650 ( .A(n2071), .B(n2072), .C(n2073), .D(n2074), .Y(n2068) );
  AOI22X1 U1651 ( .A0(n671), .A1(N474), .B0(n1723), .B1(N442), .Y(n2071) );
  AOI22X1 U1652 ( .A0(n1721), .A1(N538), .B0(n673), .B1(N506), .Y(n2072) );
  AOI22X1 U1653 ( .A0(n1717), .A1(N666), .B0(n1718), .B1(N634), .Y(n2074) );
  AOI22X1 U1654 ( .A0(n1728), .A1(N922), .B0(n1729), .B1(N890), .Y(n2084) );
  AOI22X1 U1656 ( .A0(n1728), .A1(N923), .B0(n1729), .B1(N891), .Y(n2065) );
  AOI22X1 U1657 ( .A0(n1717), .A1(N667), .B0(n1718), .B1(N635), .Y(n2061) );
  AOI22X1 U1658 ( .A0(n1728), .A1(N924), .B0(n1729), .B1(N892), .Y(n2054) );
  AOI22X1 U1659 ( .A0(n1717), .A1(N668), .B0(n1718), .B1(N636), .Y(n2050) );
  AOI22X1 U1660 ( .A0(n1728), .A1(N925), .B0(n1729), .B1(N893), .Y(n2043) );
  AOI22X1 U1661 ( .A0(n1717), .A1(N669), .B0(n1718), .B1(N637), .Y(n2039) );
  AOI22X1 U1662 ( .A0(n1728), .A1(N926), .B0(n1729), .B1(N894), .Y(n2032) );
  AOI22X1 U1663 ( .A0(n1717), .A1(N670), .B0(n1718), .B1(N638), .Y(n2028) );
  AOI22X1 U1664 ( .A0(n1728), .A1(N927), .B0(n1729), .B1(N895), .Y(n2021) );
  AOI22X1 U1665 ( .A0(n1717), .A1(N671), .B0(n1718), .B1(N639), .Y(n2017) );
  AOI22X1 U1666 ( .A0(n1728), .A1(N928), .B0(n1729), .B1(N896), .Y(n2010) );
  AOI22X1 U1667 ( .A0(n1717), .A1(N672), .B0(n1718), .B1(N640), .Y(n2006) );
  AOI22X1 U1668 ( .A0(n1728), .A1(N929), .B0(n1729), .B1(N897), .Y(n1999) );
  AOI22X1 U1669 ( .A0(n1717), .A1(N673), .B0(n1718), .B1(N641), .Y(n1995) );
  AOI22X1 U1670 ( .A0(n1728), .A1(N930), .B0(n1729), .B1(N898), .Y(n1988) );
  AOI22X1 U1671 ( .A0(n1717), .A1(N674), .B0(n1718), .B1(N642), .Y(n1984) );
  AOI22X1 U1672 ( .A0(n1728), .A1(N931), .B0(n1729), .B1(N899), .Y(n1977) );
  AOI22X1 U1673 ( .A0(n1717), .A1(N675), .B0(n1718), .B1(N643), .Y(n1973) );
  AOI22X1 U1674 ( .A0(n1728), .A1(N932), .B0(n1729), .B1(N900), .Y(n1966) );
  AOI22X1 U1675 ( .A0(n1717), .A1(N676), .B0(n1718), .B1(N644), .Y(n1962) );
  AOI22X1 U1676 ( .A0(n1728), .A1(N933), .B0(n1729), .B1(N901), .Y(n1955) );
  AOI22X1 U1677 ( .A0(n1717), .A1(N677), .B0(n1718), .B1(N645), .Y(n1951) );
  AOI22X1 U1678 ( .A0(n1728), .A1(N934), .B0(n1729), .B1(N902), .Y(n1944) );
  AOI22X1 U1679 ( .A0(n1717), .A1(N678), .B0(n1718), .B1(N646), .Y(n1940) );
  AOI22X1 U1680 ( .A0(n1728), .A1(N935), .B0(n1729), .B1(N903), .Y(n1933) );
  AOI22X1 U1681 ( .A0(n1717), .A1(N679), .B0(n1718), .B1(N647), .Y(n1929) );
  AOI22X1 U1682 ( .A0(n1728), .A1(N936), .B0(n1729), .B1(N904), .Y(n1922) );
  AOI22X1 U1683 ( .A0(n1717), .A1(N680), .B0(n1718), .B1(N648), .Y(n1918) );
  AOI22X1 U1684 ( .A0(n1728), .A1(N937), .B0(n1729), .B1(N905), .Y(n1911) );
  AOI22X1 U1685 ( .A0(n1717), .A1(N681), .B0(n1718), .B1(N649), .Y(n1907) );
  AOI22X1 U1686 ( .A0(n1728), .A1(N938), .B0(n1729), .B1(N906), .Y(n1900) );
  AOI22X1 U1687 ( .A0(n1717), .A1(N682), .B0(n1718), .B1(N650), .Y(n1896) );
  AOI22X1 U1688 ( .A0(n1728), .A1(N939), .B0(n1729), .B1(N907), .Y(n1889) );
  AOI22X1 U1689 ( .A0(n1717), .A1(N683), .B0(n1718), .B1(N651), .Y(n1885) );
  AOI22X1 U1690 ( .A0(n1728), .A1(N940), .B0(n1729), .B1(N908), .Y(n1878) );
  AOI22X1 U1691 ( .A0(n1717), .A1(N684), .B0(n1718), .B1(N652), .Y(n1874) );
  AOI22X1 U1692 ( .A0(n1728), .A1(N941), .B0(n1729), .B1(N909), .Y(n1867) );
  AOI22X1 U1693 ( .A0(n1717), .A1(N685), .B0(n1718), .B1(N653), .Y(n1863) );
  AOI22X1 U1694 ( .A0(n1721), .A1(N558), .B0(n674), .B1(N526), .Y(n1850) );
  AOI22X1 U1695 ( .A0(n1721), .A1(N559), .B0(n674), .B1(N527), .Y(n1839) );
  AOI22X1 U1696 ( .A0(n1721), .A1(N560), .B0(n674), .B1(N528), .Y(n1828) );
  AOI22X1 U1697 ( .A0(n1721), .A1(N561), .B0(n674), .B1(N529), .Y(n1817) );
  AOI22X1 U1698 ( .A0(n1719), .A1(N602), .B0(n1720), .B1(N570), .Y(n2073) );
  AOI22X1 U1699 ( .A0(n1719), .A1(N603), .B0(n1720), .B1(N571), .Y(n2060) );
  AOI22X1 U1700 ( .A0(n1719), .A1(N604), .B0(n1720), .B1(N572), .Y(n2049) );
  AOI22X1 U1701 ( .A0(n1719), .A1(N605), .B0(n1720), .B1(N573), .Y(n2038) );
  AOI22X1 U1702 ( .A0(n1719), .A1(N606), .B0(n1720), .B1(N574), .Y(n2027) );
  AOI22X1 U1703 ( .A0(n1719), .A1(N607), .B0(n1720), .B1(N575), .Y(n2016) );
  AOI22X1 U1704 ( .A0(n1719), .A1(N608), .B0(n1720), .B1(N576), .Y(n2005) );
  AOI22X1 U1705 ( .A0(n1719), .A1(N609), .B0(n1720), .B1(N577), .Y(n1994) );
  AOI22X1 U1706 ( .A0(n1719), .A1(N610), .B0(n1720), .B1(N578), .Y(n1983) );
  AOI22X1 U1707 ( .A0(n1719), .A1(N611), .B0(n1720), .B1(N579), .Y(n1972) );
  AOI22X1 U1708 ( .A0(n1719), .A1(N612), .B0(n1720), .B1(N580), .Y(n1961) );
  AOI22X1 U1709 ( .A0(n1719), .A1(N613), .B0(n1720), .B1(N581), .Y(n1950) );
  AOI22X1 U1710 ( .A0(n1719), .A1(N614), .B0(n1720), .B1(N582), .Y(n1939) );
  AOI22X1 U1711 ( .A0(n1719), .A1(N615), .B0(n1720), .B1(N583), .Y(n1928) );
  AOI22X1 U1712 ( .A0(n1719), .A1(N616), .B0(n1720), .B1(N584), .Y(n1917) );
  AOI22X1 U1713 ( .A0(n1719), .A1(N617), .B0(n1720), .B1(N585), .Y(n1906) );
  AOI22X1 U1714 ( .A0(n1719), .A1(N618), .B0(n1720), .B1(N586), .Y(n1895) );
  AOI22X1 U1715 ( .A0(n1719), .A1(N619), .B0(n1720), .B1(N587), .Y(n1884) );
  AOI22X1 U1716 ( .A0(n1719), .A1(N620), .B0(n1720), .B1(N588), .Y(n1873) );
  AOI22X1 U1717 ( .A0(n1719), .A1(N621), .B0(n1720), .B1(N589), .Y(n1862) );
  AOI22X1 U1718 ( .A0(n672), .A1(N494), .B0(n1723), .B1(N462), .Y(n1849) );
  AOI22X1 U1719 ( .A0(n672), .A1(N495), .B0(n1723), .B1(N463), .Y(n1838) );
  AOI22X1 U1720 ( .A0(n672), .A1(N496), .B0(n1723), .B1(N464), .Y(n1827) );
  AOI22X1 U1721 ( .A0(n672), .A1(N497), .B0(n1723), .B1(N465), .Y(n1816) );
  AOI22X1 U1722 ( .A0(n1721), .A1(buffer[96]), .B0(n673), .B1(buffer[104]), 
        .Y(n1806) );
  AOI22X1 U1723 ( .A0(n1721), .A1(buffer[97]), .B0(n674), .B1(buffer[105]), 
        .Y(n1795) );
  AOI22X1 U1724 ( .A0(n1721), .A1(buffer[98]), .B0(n673), .B1(buffer[106]), 
        .Y(n1784) );
  AOI22X1 U1725 ( .A0(n1721), .A1(buffer[99]), .B0(n674), .B1(buffer[107]), 
        .Y(n1773) );
  AOI22X1 U1726 ( .A0(n1721), .A1(buffer[100]), .B0(n673), .B1(buffer[108]), 
        .Y(n1762) );
  AOI22X1 U1727 ( .A0(n1721), .A1(buffer[101]), .B0(n674), .B1(buffer[109]), 
        .Y(n1751) );
  AOI22X1 U1728 ( .A0(n1721), .A1(buffer[102]), .B0(n674), .B1(buffer[110]), 
        .Y(n1740) );
  AOI22X1 U1729 ( .A0(n1721), .A1(buffer[103]), .B0(n674), .B1(buffer[111]), 
        .Y(n1714) );
  AOI22X1 U1730 ( .A0(n1721), .A1(N539), .B0(n673), .B1(N507), .Y(n2059) );
  AOI22X1 U1731 ( .A0(n1721), .A1(N540), .B0(n673), .B1(N508), .Y(n2048) );
  AOI22X1 U1732 ( .A0(n1721), .A1(N541), .B0(n673), .B1(N509), .Y(n2037) );
  AOI22X1 U1733 ( .A0(n1721), .A1(N542), .B0(n673), .B1(N510), .Y(n2026) );
  AOI22X1 U1734 ( .A0(n1721), .A1(N543), .B0(n673), .B1(N511), .Y(n2015) );
  AOI22X1 U1735 ( .A0(n1721), .A1(N544), .B0(n673), .B1(N512), .Y(n2004) );
  AOI22X1 U1736 ( .A0(n1721), .A1(N545), .B0(n673), .B1(N513), .Y(n1993) );
  AOI22X1 U1737 ( .A0(n1721), .A1(N546), .B0(n673), .B1(N514), .Y(n1982) );
  AOI22X1 U1738 ( .A0(n1721), .A1(N547), .B0(n673), .B1(N515), .Y(n1971) );
  AOI22X1 U1739 ( .A0(n1721), .A1(N548), .B0(n673), .B1(N516), .Y(n1960) );
  AOI22X1 U1740 ( .A0(n1721), .A1(N549), .B0(n673), .B1(N517), .Y(n1949) );
  AOI22X1 U1741 ( .A0(n1721), .A1(N550), .B0(n674), .B1(N518), .Y(n1938) );
  AOI22X1 U1742 ( .A0(n1721), .A1(N551), .B0(n674), .B1(N519), .Y(n1927) );
  AOI22X1 U1743 ( .A0(n1721), .A1(N552), .B0(n674), .B1(N520), .Y(n1916) );
  AOI22X1 U1744 ( .A0(n1721), .A1(N553), .B0(n674), .B1(N521), .Y(n1905) );
  AOI22X1 U1745 ( .A0(n1721), .A1(N554), .B0(n674), .B1(N522), .Y(n1894) );
  AOI22X1 U1746 ( .A0(n1721), .A1(N555), .B0(n674), .B1(N523), .Y(n1883) );
  AOI22X1 U1747 ( .A0(n1721), .A1(N556), .B0(n674), .B1(N524), .Y(n1872) );
  AOI22X1 U1748 ( .A0(n1721), .A1(N557), .B0(n674), .B1(N525), .Y(n1861) );
  AOI22X1 U1749 ( .A0(n1728), .A1(N942), .B0(n1729), .B1(N910), .Y(n1856) );
  AOI22X1 U1750 ( .A0(n1717), .A1(N686), .B0(n1718), .B1(N654), .Y(n1852) );
  AOI22X1 U1751 ( .A0(n1728), .A1(N943), .B0(n1729), .B1(N911), .Y(n1845) );
  AOI22X1 U1752 ( .A0(n1717), .A1(N687), .B0(n1718), .B1(N655), .Y(n1841) );
  AOI22X1 U1753 ( .A0(n1728), .A1(N944), .B0(n1729), .B1(N912), .Y(n1834) );
  AOI22X1 U1754 ( .A0(n1717), .A1(N688), .B0(n1718), .B1(N656), .Y(n1830) );
  AOI22X1 U1755 ( .A0(n1728), .A1(N945), .B0(n1729), .B1(N913), .Y(n1823) );
  AOI22X1 U1756 ( .A0(n1717), .A1(N689), .B0(n1718), .B1(N657), .Y(n1819) );
  AOI22X1 U1757 ( .A0(n671), .A1(N475), .B0(n1723), .B1(N443), .Y(n2058) );
  AOI22X1 U1758 ( .A0(n671), .A1(N476), .B0(n1723), .B1(N444), .Y(n2047) );
  AOI22X1 U1759 ( .A0(n671), .A1(N477), .B0(n1723), .B1(N445), .Y(n2036) );
  AOI22X1 U1760 ( .A0(n671), .A1(N478), .B0(n1723), .B1(N446), .Y(n2025) );
  AOI22X1 U1761 ( .A0(n671), .A1(N479), .B0(n1723), .B1(N447), .Y(n2014) );
  AOI22X1 U1762 ( .A0(n671), .A1(N480), .B0(n1723), .B1(N448), .Y(n2003) );
  AOI22X1 U1763 ( .A0(n671), .A1(N481), .B0(n1723), .B1(N449), .Y(n1992) );
  AOI22X1 U1764 ( .A0(n671), .A1(N482), .B0(n1723), .B1(N450), .Y(n1981) );
  AOI22X1 U1765 ( .A0(n671), .A1(N483), .B0(n1723), .B1(N451), .Y(n1970) );
  AOI22X1 U1766 ( .A0(n671), .A1(N484), .B0(n1723), .B1(N452), .Y(n1959) );
  AOI22X1 U1767 ( .A0(n671), .A1(N485), .B0(n1723), .B1(N453), .Y(n1948) );
  AOI22X1 U1768 ( .A0(n672), .A1(N486), .B0(n1723), .B1(N454), .Y(n1937) );
  AOI22X1 U1769 ( .A0(n672), .A1(N487), .B0(n1723), .B1(N455), .Y(n1926) );
  AOI22X1 U1770 ( .A0(n672), .A1(N488), .B0(n1723), .B1(N456), .Y(n1915) );
  AOI22X1 U1771 ( .A0(n672), .A1(N489), .B0(n1723), .B1(N457), .Y(n1904) );
  AOI22X1 U1772 ( .A0(n672), .A1(N490), .B0(n1723), .B1(N458), .Y(n1893) );
  AOI22X1 U1773 ( .A0(n672), .A1(N491), .B0(n1723), .B1(N459), .Y(n1882) );
  AOI22X1 U1774 ( .A0(n672), .A1(N492), .B0(n1723), .B1(N460), .Y(n1871) );
  AOI22X1 U1775 ( .A0(n672), .A1(N493), .B0(n1723), .B1(N461), .Y(n1860) );
  AOI22X1 U1776 ( .A0(n1719), .A1(N622), .B0(n1720), .B1(N590), .Y(n1851) );
  AOI22X1 U1777 ( .A0(n1719), .A1(N623), .B0(n1720), .B1(N591), .Y(n1840) );
  AOI22X1 U1778 ( .A0(n1719), .A1(N624), .B0(n1720), .B1(N592), .Y(n1829) );
  AOI22X1 U1779 ( .A0(n1719), .A1(N625), .B0(n1720), .B1(N593), .Y(n1818) );
  AOI22X1 U1780 ( .A0(n671), .A1(buffer[112]), .B0(n1723), .B1(buffer[120]), 
        .Y(n1805) );
  AOI22X1 U1781 ( .A0(n672), .A1(buffer[113]), .B0(n1723), .B1(buffer[121]), 
        .Y(n1794) );
  AOI22X1 U1782 ( .A0(n672), .A1(buffer[114]), .B0(n1723), .B1(buffer[122]), 
        .Y(n1783) );
  AOI22X1 U1783 ( .A0(n672), .A1(buffer[115]), .B0(n1723), .B1(buffer[123]), 
        .Y(n1772) );
  AOI22X1 U1784 ( .A0(n671), .A1(buffer[116]), .B0(n1723), .B1(buffer[124]), 
        .Y(n1761) );
  AOI22X1 U1785 ( .A0(n671), .A1(buffer[117]), .B0(n1723), .B1(buffer[125]), 
        .Y(n1750) );
  AOI22X1 U1786 ( .A0(n671), .A1(buffer[118]), .B0(n1723), .B1(buffer[126]), 
        .Y(n1739) );
  AOI22X1 U1787 ( .A0(n672), .A1(buffer[119]), .B0(n1723), .B1(buffer[127]), 
        .Y(n1713) );
  AOI22X1 U1788 ( .A0(n1728), .A1(buffer[0]), .B0(n1729), .B1(buffer[8]), .Y(
        n1812) );
  AOI22X1 U1789 ( .A0(n1717), .A1(buffer[64]), .B0(n1718), .B1(buffer[72]), 
        .Y(n1808) );
  AOI22X1 U1790 ( .A0(n1728), .A1(buffer[1]), .B0(n1729), .B1(buffer[9]), .Y(
        n1801) );
  AOI22X1 U1791 ( .A0(n1717), .A1(buffer[65]), .B0(n1718), .B1(buffer[73]), 
        .Y(n1797) );
  AOI22X1 U1792 ( .A0(n1728), .A1(buffer[2]), .B0(n1729), .B1(buffer[10]), .Y(
        n1790) );
  AOI22X1 U1793 ( .A0(n1717), .A1(buffer[66]), .B0(n1718), .B1(buffer[74]), 
        .Y(n1786) );
  AOI22X1 U1794 ( .A0(n1728), .A1(buffer[3]), .B0(n1729), .B1(buffer[11]), .Y(
        n1779) );
  AOI22X1 U1795 ( .A0(n1717), .A1(buffer[67]), .B0(n1718), .B1(buffer[75]), 
        .Y(n1775) );
  AOI22X1 U1796 ( .A0(n1728), .A1(buffer[4]), .B0(n1729), .B1(buffer[12]), .Y(
        n1768) );
  AOI22X1 U1797 ( .A0(n1717), .A1(buffer[68]), .B0(n1718), .B1(buffer[76]), 
        .Y(n1764) );
  AOI22X1 U1798 ( .A0(n1728), .A1(buffer[5]), .B0(n1729), .B1(buffer[13]), .Y(
        n1757) );
  AOI22X1 U1799 ( .A0(n1717), .A1(buffer[69]), .B0(n1718), .B1(buffer[77]), 
        .Y(n1753) );
  AOI22X1 U1800 ( .A0(n1728), .A1(buffer[6]), .B0(n1729), .B1(buffer[14]), .Y(
        n1746) );
  AOI22X1 U1801 ( .A0(n1717), .A1(buffer[70]), .B0(n1718), .B1(buffer[78]), 
        .Y(n1742) );
  AOI22X1 U1802 ( .A0(n1728), .A1(buffer[7]), .B0(n1729), .B1(buffer[15]), .Y(
        n1727) );
  AOI22X1 U1803 ( .A0(n1717), .A1(buffer[71]), .B0(n1718), .B1(buffer[79]), 
        .Y(n1716) );
  AOI22X1 U1804 ( .A0(n1719), .A1(buffer[80]), .B0(n1720), .B1(buffer[88]), 
        .Y(n1807) );
  AOI22X1 U1805 ( .A0(n1719), .A1(buffer[81]), .B0(n1720), .B1(buffer[89]), 
        .Y(n1796) );
  AOI22X1 U1806 ( .A0(n1719), .A1(buffer[82]), .B0(n1720), .B1(buffer[90]), 
        .Y(n1785) );
  AOI22X1 U1807 ( .A0(n1719), .A1(buffer[83]), .B0(n1720), .B1(buffer[91]), 
        .Y(n1774) );
  AOI22X1 U1808 ( .A0(n1719), .A1(buffer[84]), .B0(n1720), .B1(buffer[92]), 
        .Y(n1763) );
  AOI22X1 U1809 ( .A0(n1719), .A1(buffer[85]), .B0(n1720), .B1(buffer[93]), 
        .Y(n1752) );
  AOI22X1 U1810 ( .A0(n1719), .A1(buffer[86]), .B0(n1720), .B1(buffer[94]), 
        .Y(n1741) );
  AOI22X1 U1811 ( .A0(n1719), .A1(buffer[87]), .B0(n1720), .B1(buffer[95]), 
        .Y(n1715) );
  OR2X2 U1812 ( .A(n546), .B(counter2[4]), .Y(n746) );
  OR2X2 U1813 ( .A(counter2[5]), .B(counter2[6]), .Y(n546) );
endmodule


module hash_core_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
endmodule


module hash_core_DW01_add_16 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223;

  OAI21X2 U2 ( .A0(n195), .A1(n171), .B0(n176), .Y(n193) );
  INVX2 U3 ( .A(n204), .Y(n203) );
  CLKINVX3 U4 ( .A(n155), .Y(n154) );
  INVX2 U5 ( .A(n27), .Y(n24) );
  INVX2 U6 ( .A(n33), .Y(n30) );
  AOI21X4 U7 ( .A0(n172), .A1(n177), .B0(n178), .Y(n175) );
  INVX4 U8 ( .A(n150), .Y(n132) );
  NOR2X4 U9 ( .A(n82), .B(n83), .Y(n75) );
  CLKINVX3 U10 ( .A(n215), .Y(n31) );
  NOR2X1 U11 ( .A(n218), .B(n180), .Y(n7) );
  CLKINVX8 U12 ( .A(n179), .Y(n178) );
  OAI21X4 U13 ( .A0(n186), .A1(n170), .B0(n168), .Y(n184) );
  INVX4 U14 ( .A(n187), .Y(n186) );
  NOR2X4 U15 ( .A(n169), .B(n170), .Y(n162) );
  XOR2X2 U16 ( .A(n148), .B(n149), .Y(SUM[19]) );
  NOR2X4 U17 ( .A(n51), .B(n52), .Y(n47) );
  NOR2X2 U18 ( .A(A[30]), .B(B[30]), .Y(n52) );
  OAI21X4 U19 ( .A0(n89), .A1(n83), .B0(n90), .Y(n87) );
  NAND2X2 U20 ( .A(B[13]), .B(A[13]), .Y(n167) );
  INVX4 U21 ( .A(n16), .Y(n195) );
  NAND3BX4 U22 ( .AN(n129), .B(n130), .C(n131), .Y(n128) );
  NOR2X2 U23 ( .A(n132), .B(n133), .Y(n131) );
  NOR2X2 U24 ( .A(n133), .B(n132), .Y(n136) );
  INVX4 U25 ( .A(n144), .Y(n133) );
  INVX4 U26 ( .A(n177), .Y(n218) );
  OAI21X4 U27 ( .A0(n220), .A1(n221), .B0(n39), .Y(n177) );
  OAI21X2 U28 ( .A0(n118), .A1(n113), .B0(n111), .Y(n116) );
  NAND2X2 U29 ( .A(B[8]), .B(A[8]), .Y(n18) );
  NOR2BX1 U30 ( .AN(n111), .B(n113), .Y(n120) );
  OR2X2 U31 ( .A(A[5]), .B(B[5]), .Y(n215) );
  OR2X2 U32 ( .A(A[1]), .B(B[1]), .Y(n64) );
  CLKINVX3 U33 ( .A(n86), .Y(n82) );
  OR2X2 U34 ( .A(A[19]), .B(B[19]), .Y(n144) );
  INVX1 U35 ( .A(n53), .Y(n51) );
  NAND2X1 U36 ( .A(B[29]), .B(A[29]), .Y(n57) );
  NAND2X1 U37 ( .A(n157), .B(n141), .Y(n155) );
  OAI2BB1X1 U38 ( .A0N(n189), .A1N(n6), .B0(n167), .Y(n187) );
  INVX2 U39 ( .A(n182), .Y(n170) );
  NAND2X2 U40 ( .A(B[12]), .B(A[12]), .Y(n166) );
  NAND2X2 U41 ( .A(B[11]), .B(A[11]), .Y(n204) );
  CLKINVX3 U42 ( .A(n200), .Y(n15) );
  OAI21XL U43 ( .A0(n11), .A1(n218), .B0(n35), .Y(n33) );
  OAI21XL U44 ( .A0(n24), .A1(n25), .B0(n26), .Y(n20) );
  INVX1 U45 ( .A(n107), .Y(n106) );
  AOI21X1 U46 ( .A0(n199), .A1(n208), .B0(n209), .Y(n207) );
  XOR2X1 U47 ( .A(n119), .B(n120), .Y(SUM[22]) );
  NAND2X2 U48 ( .A(n14), .B(n18), .Y(n201) );
  NAND2X2 U49 ( .A(B[18]), .B(A[18]), .Y(n143) );
  NAND2X1 U50 ( .A(B[17]), .B(A[17]), .Y(n142) );
  INVX1 U51 ( .A(n78), .Y(n77) );
  AOI21X4 U52 ( .A0(n162), .A1(n163), .B0(n164), .Y(n161) );
  INVX2 U53 ( .A(n135), .Y(n140) );
  INVX4 U54 ( .A(n94), .Y(n84) );
  AOI21X4 U55 ( .A0(n75), .A1(n76), .B0(n77), .Y(n74) );
  NAND2BX4 U56 ( .AN(n173), .B(n174), .Y(n160) );
  OAI2BB1X2 U57 ( .A0N(n12), .A1N(n200), .B0(n14), .Y(n208) );
  NAND2XL U58 ( .A(n212), .B(n18), .Y(n12) );
  XOR2X4 U59 ( .A(n184), .B(n185), .Y(SUM[15]) );
  NAND2X2 U60 ( .A(B[6]), .B(A[6]), .Y(n26) );
  XOR2X2 U61 ( .A(n91), .B(n92), .Y(SUM[26]) );
  XNOR2X2 U62 ( .A(B[31]), .B(A[31]), .Y(n45) );
  OAI2BB1X4 U63 ( .A0N(n1), .A1N(n2), .B0(n50), .Y(n49) );
  OR2X4 U64 ( .A(A[30]), .B(B[30]), .Y(n1) );
  AND2X1 U65 ( .A(A[29]), .B(B[29]), .Y(n2) );
  NAND2X1 U66 ( .A(B[3]), .B(n5), .Y(n39) );
  OAI21X4 U67 ( .A0(n58), .A1(n59), .B0(n60), .Y(n3) );
  OR2X2 U68 ( .A(A[8]), .B(B[8]), .Y(n205) );
  INVX8 U69 ( .A(n121), .Y(n108) );
  BUFX4 U70 ( .A(n110), .Y(n8) );
  BUFX4 U71 ( .A(n125), .Y(n4) );
  AND2X1 U72 ( .A(n109), .B(n4), .Y(n126) );
  NAND2X4 U73 ( .A(B[22]), .B(A[22]), .Y(n111) );
  XNOR2X1 U74 ( .A(B[30]), .B(A[30]), .Y(n54) );
  INVX4 U75 ( .A(n91), .Y(n89) );
  NAND3BX2 U76 ( .AN(n108), .B(n114), .C(n115), .Y(n102) );
  NAND2X1 U77 ( .A(B[21]), .B(A[21]), .Y(n110) );
  INVX8 U78 ( .A(n69), .Y(n59) );
  NAND2X4 U79 ( .A(n93), .B(n80), .Y(n91) );
  NAND2X4 U80 ( .A(n94), .B(n95), .Y(n93) );
  NAND4BBX4 U81 ( .AN(n19), .BN(n15), .C(n199), .D(n198), .Y(n171) );
  AOI21X2 U82 ( .A0(n61), .A1(n69), .B0(n70), .Y(n68) );
  NAND2X4 U83 ( .A(B[28]), .B(A[28]), .Y(n60) );
  AOI21X4 U84 ( .A0(n47), .A1(n3), .B0(n49), .Y(n46) );
  NAND3X1 U85 ( .A(n215), .B(n29), .C(n216), .Y(n214) );
  OAI21X4 U86 ( .A0(n72), .A1(n73), .B0(n74), .Y(n69) );
  OAI2BB1X4 U87 ( .A0N(n196), .A1N(n197), .B0(n198), .Y(n176) );
  NOR2BX2 U88 ( .AN(n202), .B(n203), .Y(n196) );
  NAND3X1 U89 ( .A(n199), .B(n200), .C(n201), .Y(n197) );
  NAND2X4 U90 ( .A(B[24]), .B(A[24]), .Y(n97) );
  AOI21X2 U91 ( .A0(n136), .A1(n137), .B0(n138), .Y(n127) );
  INVX4 U92 ( .A(n193), .Y(n192) );
  OAI211X2 U93 ( .A0(n140), .A1(n141), .B0(n142), .C0(n143), .Y(n137) );
  NAND2X4 U94 ( .A(n160), .B(n161), .Y(n130) );
  NAND3BX1 U95 ( .AN(n84), .B(n85), .C(n86), .Y(n73) );
  CLKINVX2 U96 ( .A(n180), .Y(n172) );
  NAND2X4 U97 ( .A(B[23]), .B(A[23]), .Y(n107) );
  NAND2X2 U98 ( .A(A[24]), .B(B[24]), .Y(n79) );
  NAND2X2 U99 ( .A(B[25]), .B(A[25]), .Y(n80) );
  NOR2BX2 U100 ( .AN(n26), .B(n217), .Y(n213) );
  AOI21X4 U101 ( .A0(n53), .A1(n48), .B0(n56), .Y(n55) );
  NOR2BXL U102 ( .AN(n168), .B(n170), .Y(n188) );
  NAND2X2 U103 ( .A(B[14]), .B(A[14]), .Y(n168) );
  XOR2X4 U104 ( .A(n46), .B(n45), .Y(SUM[31]) );
  XOR2X2 U105 ( .A(n206), .B(n207), .Y(SUM[11]) );
  OAI21X4 U106 ( .A0(n175), .A1(n171), .B0(n176), .Y(n174) );
  AOI21X2 U107 ( .A0(n150), .A1(n151), .B0(n152), .Y(n149) );
  OAI211X2 U108 ( .A0(n84), .A1(n79), .B0(n80), .C0(n81), .Y(n76) );
  XOR2X1 U109 ( .A(n71), .B(n59), .Y(SUM[28]) );
  OAI211X2 U110 ( .A0(n108), .A1(n109), .B0(n8), .C0(n111), .Y(n105) );
  AOI21X4 U111 ( .A0(n104), .A1(n105), .B0(n106), .Y(n103) );
  NOR2X4 U112 ( .A(n112), .B(n113), .Y(n104) );
  INVX4 U113 ( .A(n114), .Y(n113) );
  INVX4 U114 ( .A(n115), .Y(n112) );
  XOR2X4 U115 ( .A(n54), .B(n55), .Y(SUM[30]) );
  XOR2X2 U116 ( .A(n116), .B(n117), .Y(SUM[23]) );
  XOR2X4 U117 ( .A(n87), .B(n88), .Y(SUM[27]) );
  OAI21X2 U118 ( .A0(n154), .A1(n140), .B0(n142), .Y(n151) );
  OAI21X4 U119 ( .A0(n191), .A1(n192), .B0(n166), .Y(n189) );
  CLKBUFXL U120 ( .A(A[3]), .Y(n5) );
  NAND2X1 U121 ( .A(n101), .B(n109), .Y(n122) );
  NAND2X4 U122 ( .A(n124), .B(n4), .Y(n101) );
  INVX2 U123 ( .A(n119), .Y(n118) );
  OAI21X4 U124 ( .A0(n58), .A1(n59), .B0(n60), .Y(n48) );
  OAI2BB1XL U125 ( .A0N(n64), .A1N(n65), .B0(n66), .Y(n44) );
  NOR2BX1 U126 ( .AN(n66), .B(n146), .Y(n145) );
  OAI21X2 U127 ( .A0(n146), .A1(n147), .B0(n66), .Y(n223) );
  NAND2X4 U128 ( .A(B[20]), .B(A[20]), .Y(n109) );
  NAND2X2 U129 ( .A(n72), .B(n97), .Y(n95) );
  NAND2X4 U130 ( .A(n98), .B(n99), .Y(n72) );
  NAND2X2 U131 ( .A(B[2]), .B(A[2]), .Y(n43) );
  OR2XL U132 ( .A(A[2]), .B(B[2]), .Y(n63) );
  NOR2X4 U133 ( .A(A[13]), .B(B[13]), .Y(n10) );
  OR2X2 U134 ( .A(n7), .B(n178), .Y(n16) );
  OAI21X4 U135 ( .A0(n101), .A1(n102), .B0(n103), .Y(n98) );
  NAND2XL U136 ( .A(n16), .B(n205), .Y(n212) );
  OAI2BB1X2 U137 ( .A0N(n121), .A1N(n122), .B0(n8), .Y(n119) );
  XOR2X1 U138 ( .A(n16), .B(n17), .Y(SUM[8]) );
  INVX1 U139 ( .A(n10), .Y(n6) );
  OAI2BB1X4 U140 ( .A0N(n213), .A1N(n214), .B0(n23), .Y(n179) );
  CLKINVX3 U141 ( .A(n139), .Y(n138) );
  INVX2 U142 ( .A(n61), .Y(n58) );
  NAND2X2 U143 ( .A(B[7]), .B(A[7]), .Y(n22) );
  NAND2XL U144 ( .A(B[1]), .B(A[1]), .Y(n66) );
  OR2XL U145 ( .A(A[20]), .B(B[20]), .Y(n125) );
  INVX1 U146 ( .A(n64), .Y(n146) );
  OR2X2 U147 ( .A(A[24]), .B(B[24]), .Y(n99) );
  NOR2X1 U148 ( .A(A[4]), .B(B[4]), .Y(n11) );
  NAND2X4 U149 ( .A(B[9]), .B(A[9]), .Y(n14) );
  NAND2X2 U150 ( .A(B[5]), .B(A[5]), .Y(n32) );
  NAND4BX1 U151 ( .AN(n10), .B(n181), .C(n182), .D(n183), .Y(n173) );
  NAND2XL U152 ( .A(n53), .B(n57), .Y(n67) );
  NAND2X1 U153 ( .A(n134), .B(n135), .Y(n129) );
  CLKINVX3 U154 ( .A(n165), .Y(n164) );
  INVXL U155 ( .A(n202), .Y(n209) );
  NAND2XL U156 ( .A(n60), .B(n61), .Y(n71) );
  INVXL U157 ( .A(n181), .Y(n191) );
  INVXL U158 ( .A(n134), .Y(n159) );
  AND2X1 U159 ( .A(n97), .B(n99), .Y(n100) );
  INVXL U160 ( .A(n29), .Y(n25) );
  INVXL U161 ( .A(n219), .Y(n40) );
  AND2X1 U162 ( .A(n22), .B(n23), .Y(n21) );
  INVXL U163 ( .A(n147), .Y(n65) );
  NAND2X2 U164 ( .A(B[4]), .B(A[4]), .Y(n35) );
  NAND2XL U165 ( .A(B[27]), .B(A[27]), .Y(n78) );
  NAND2XL U166 ( .A(B[30]), .B(A[30]), .Y(n50) );
  NOR2BX1 U167 ( .AN(n147), .B(n9), .Y(SUM[0]) );
  NOR2XL U168 ( .A(A[0]), .B(B[0]), .Y(n9) );
  NAND2X1 U169 ( .A(n63), .B(n219), .Y(n221) );
  NOR2X1 U170 ( .A(n222), .B(n223), .Y(n220) );
  INVX1 U171 ( .A(n43), .Y(n222) );
  NAND4BBX2 U172 ( .AN(n31), .BN(n11), .C(n29), .D(n23), .Y(n180) );
  NOR2BXL U173 ( .AN(n90), .B(n83), .Y(n92) );
  NOR2BXL U174 ( .AN(n143), .B(n132), .Y(n153) );
  NOR2BXL U175 ( .AN(n8), .B(n108), .Y(n123) );
  NOR2BXL U176 ( .AN(n107), .B(n112), .Y(n117) );
  NAND2XL U177 ( .A(n130), .B(n134), .Y(n157) );
  XOR2X1 U178 ( .A(n155), .B(n156), .Y(SUM[17]) );
  NOR2BXL U179 ( .AN(n142), .B(n140), .Y(n156) );
  XOR2X1 U180 ( .A(n208), .B(n210), .Y(SUM[10]) );
  NOR2BX1 U181 ( .AN(n202), .B(n211), .Y(n210) );
  INVXL U182 ( .A(n199), .Y(n211) );
  XOR2X1 U183 ( .A(n187), .B(n188), .Y(SUM[14]) );
  XOR2X1 U184 ( .A(n189), .B(n190), .Y(SUM[13]) );
  NOR2BX1 U185 ( .AN(n167), .B(n10), .Y(n190) );
  XOR2X1 U186 ( .A(n130), .B(n158), .Y(SUM[16]) );
  NOR2BX1 U187 ( .AN(n141), .B(n159), .Y(n158) );
  XOR2X1 U188 ( .A(n67), .B(n68), .Y(SUM[29]) );
  INVX1 U189 ( .A(n60), .Y(n70) );
  NAND2XL U190 ( .A(n139), .B(n144), .Y(n148) );
  INVX1 U191 ( .A(n143), .Y(n152) );
  NOR2BXL U192 ( .AN(n78), .B(n82), .Y(n88) );
  XOR2X1 U193 ( .A(n95), .B(n96), .Y(SUM[25]) );
  NOR2BXL U194 ( .AN(n80), .B(n84), .Y(n96) );
  NOR2BXL U195 ( .AN(n165), .B(n169), .Y(n185) );
  XOR2X1 U196 ( .A(n33), .B(n34), .Y(SUM[5]) );
  NOR2BXL U197 ( .AN(n32), .B(n31), .Y(n34) );
  XOR2X1 U198 ( .A(n12), .B(n13), .Y(SUM[9]) );
  NOR2BXL U199 ( .AN(n14), .B(n15), .Y(n13) );
  XOR2X1 U200 ( .A(n27), .B(n28), .Y(SUM[6]) );
  NOR2BX1 U201 ( .AN(n26), .B(n25), .Y(n28) );
  XOR2X1 U202 ( .A(n44), .B(n62), .Y(SUM[2]) );
  NOR2BX1 U203 ( .AN(n43), .B(n42), .Y(n62) );
  XOR2X1 U204 ( .A(n65), .B(n145), .Y(SUM[1]) );
  INVX1 U205 ( .A(n22), .Y(n217) );
  NAND2X1 U206 ( .A(n32), .B(n35), .Y(n216) );
  XOR2X1 U207 ( .A(n193), .B(n194), .Y(SUM[12]) );
  NOR2BX1 U208 ( .AN(n166), .B(n191), .Y(n194) );
  XOR2X1 U209 ( .A(n98), .B(n100), .Y(SUM[24]) );
  XOR2X1 U210 ( .A(n151), .B(n153), .Y(SUM[18]) );
  XOR2X1 U211 ( .A(n122), .B(n123), .Y(SUM[21]) );
  XOR2X1 U212 ( .A(n124), .B(n126), .Y(SUM[20]) );
  XOR2X1 U213 ( .A(n20), .B(n21), .Y(SUM[7]) );
  XOR2X1 U214 ( .A(n177), .B(n36), .Y(SUM[4]) );
  OAI21XL U215 ( .A0(n30), .A1(n31), .B0(n32), .Y(n27) );
  NOR2BXL U216 ( .AN(n18), .B(n19), .Y(n17) );
  NAND2XL U217 ( .A(n198), .B(n204), .Y(n206) );
  INVX1 U218 ( .A(n63), .Y(n42) );
  NOR2BX1 U219 ( .AN(n35), .B(n11), .Y(n36) );
  XOR2X1 U220 ( .A(n37), .B(n38), .Y(SUM[3]) );
  OAI21XL U221 ( .A0(n41), .A1(n42), .B0(n43), .Y(n37) );
  NOR2BX1 U222 ( .AN(n39), .B(n40), .Y(n38) );
  INVX1 U223 ( .A(n44), .Y(n41) );
  INVX1 U224 ( .A(n57), .Y(n56) );
  NAND2XL U225 ( .A(B[26]), .B(A[26]), .Y(n81) );
  OR2X2 U226 ( .A(A[6]), .B(B[6]), .Y(n29) );
  OR2X2 U227 ( .A(A[29]), .B(B[29]), .Y(n53) );
  NAND2X2 U228 ( .A(B[10]), .B(A[10]), .Y(n202) );
  NAND2XL U229 ( .A(B[19]), .B(A[19]), .Y(n139) );
  NAND2XL U230 ( .A(B[26]), .B(A[26]), .Y(n90) );
  NAND2XL U231 ( .A(B[15]), .B(A[15]), .Y(n165) );
  OR2X2 U232 ( .A(A[12]), .B(B[12]), .Y(n181) );
  OR2X2 U233 ( .A(A[3]), .B(B[3]), .Y(n219) );
  OR2X2 U234 ( .A(A[27]), .B(B[27]), .Y(n86) );
  NAND2X1 U235 ( .A(B[0]), .B(A[0]), .Y(n147) );
  OR2X4 U236 ( .A(A[28]), .B(B[28]), .Y(n61) );
  CLKINVX3 U237 ( .A(n85), .Y(n83) );
  OR2X4 U238 ( .A(A[26]), .B(B[26]), .Y(n85) );
  OR2X4 U239 ( .A(A[25]), .B(B[25]), .Y(n94) );
  OR2X4 U240 ( .A(A[23]), .B(B[23]), .Y(n115) );
  OR2X4 U241 ( .A(A[22]), .B(B[22]), .Y(n114) );
  OR2X4 U242 ( .A(A[21]), .B(B[21]), .Y(n121) );
  NAND2X4 U243 ( .A(n127), .B(n128), .Y(n124) );
  OR2X4 U244 ( .A(A[18]), .B(B[18]), .Y(n150) );
  OR2X4 U245 ( .A(A[17]), .B(B[17]), .Y(n135) );
  OR2X4 U246 ( .A(A[16]), .B(B[16]), .Y(n134) );
  NAND2X4 U247 ( .A(B[16]), .B(A[16]), .Y(n141) );
  OAI211X2 U248 ( .A0(n10), .A1(n166), .B0(n167), .C0(n168), .Y(n163) );
  CLKINVX3 U249 ( .A(n183), .Y(n169) );
  OR2X4 U250 ( .A(A[15]), .B(B[15]), .Y(n183) );
  OR2X4 U251 ( .A(A[14]), .B(B[14]), .Y(n182) );
  CLKINVX3 U252 ( .A(n205), .Y(n19) );
  OR2X4 U253 ( .A(A[11]), .B(B[11]), .Y(n198) );
  OR2X4 U254 ( .A(A[10]), .B(B[10]), .Y(n199) );
  OR2X4 U255 ( .A(A[9]), .B(B[9]), .Y(n200) );
  OR2X4 U256 ( .A(A[7]), .B(B[7]), .Y(n23) );
endmodule


module hash_core_DW01_add_24 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n301, n302, n303, n1, n2, n3, n4, n5, n6, n7, n9, n12, n13, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300;

  NAND3X1 U2 ( .A(n243), .B(n244), .C(n245), .Y(n15) );
  NAND4BBX2 U3 ( .AN(n246), .BN(n249), .C(n247), .D(n248), .Y(n245) );
  XNOR2X2 U4 ( .A(n280), .B(n281), .Y(SUM[11]) );
  OR2X4 U5 ( .A(n241), .B(n58), .Y(n39) );
  OR3X4 U6 ( .A(n288), .B(n58), .C(n241), .Y(n287) );
  NAND2X2 U7 ( .A(n255), .B(n210), .Y(n246) );
  INVX4 U8 ( .A(n237), .Y(n277) );
  INVX8 U9 ( .A(n229), .Y(n219) );
  OR2X4 U10 ( .A(A[1]), .B(B[1]), .Y(n78) );
  BUFX8 U11 ( .A(n302), .Y(SUM[16]) );
  NAND2X4 U12 ( .A(n247), .B(n255), .Y(n220) );
  OAI21X4 U13 ( .A0(n195), .A1(n188), .B0(n196), .Y(n193) );
  NOR3X4 U14 ( .A(n4), .B(n189), .C(n191), .Y(n195) );
  AOI21XL U15 ( .A0(n111), .A1(n106), .B0(n112), .Y(n110) );
  NOR2BX1 U16 ( .AN(n49), .B(n55), .Y(n57) );
  NAND2X2 U17 ( .A(n143), .B(n144), .Y(n136) );
  AOI21X4 U18 ( .A0(n38), .A1(n295), .B0(n296), .Y(n286) );
  NAND2X2 U19 ( .A(B[27]), .B(A[27]), .Y(n99) );
  CLKINVX3 U20 ( .A(n207), .Y(n206) );
  OAI21X2 U21 ( .A0(n208), .A1(n209), .B0(n192), .Y(n207) );
  NOR2BX2 U22 ( .AN(n37), .B(n288), .Y(n295) );
  NAND2X2 U23 ( .A(n297), .B(n298), .Y(n7) );
  NAND2XL U24 ( .A(n105), .B(n122), .Y(n113) );
  OR2X2 U25 ( .A(A[24]), .B(B[24]), .Y(n105) );
  BUFX8 U26 ( .A(n301), .Y(SUM[30]) );
  BUFX8 U27 ( .A(n45), .Y(n1) );
  OAI21X2 U28 ( .A0(n219), .A1(n253), .B0(n213), .Y(n267) );
  NAND2X4 U29 ( .A(n247), .B(n230), .Y(n253) );
  NAND2X2 U30 ( .A(n230), .B(n210), .Y(n221) );
  OR2X4 U31 ( .A(A[11]), .B(B[11]), .Y(n230) );
  BUFX8 U32 ( .A(n303), .Y(SUM[13]) );
  CLKINVX8 U33 ( .A(n135), .Y(n134) );
  NAND2X4 U34 ( .A(B[22]), .B(A[22]), .Y(n141) );
  XOR2X4 U35 ( .A(n152), .B(n153), .Y(SUM[22]) );
  OAI21X2 U36 ( .A0(n95), .A1(n85), .B0(n91), .Y(n92) );
  NAND4BX2 U37 ( .AN(n104), .B(n105), .C(n106), .D(n98), .Y(n85) );
  NAND4BX1 U38 ( .AN(n151), .B(n144), .C(n131), .D(n115), .Y(n146) );
  NAND2X4 U39 ( .A(n134), .B(n143), .Y(n151) );
  NAND3BX4 U40 ( .AN(n85), .B(n86), .C(n87), .Y(n84) );
  OAI21X4 U41 ( .A0(n96), .A1(n97), .B0(n98), .Y(n91) );
  NAND2X2 U42 ( .A(n99), .B(n100), .Y(n97) );
  NAND2X2 U43 ( .A(n31), .B(n35), .Y(n278) );
  NAND3BX2 U44 ( .AN(n205), .B(n200), .C(n206), .Y(n203) );
  INVX2 U45 ( .A(n259), .Y(n13) );
  NAND2X2 U46 ( .A(B[4]), .B(A[4]), .Y(n54) );
  NOR2X1 U47 ( .A(n151), .B(n157), .Y(n154) );
  OAI21X2 U48 ( .A0(n183), .A1(n184), .B0(n185), .Y(n180) );
  INVXL U49 ( .A(n175), .Y(n182) );
  AND2X1 U50 ( .A(n192), .B(n211), .Y(n16) );
  NOR2BX1 U51 ( .AN(n31), .B(n32), .Y(n30) );
  NAND2XL U52 ( .A(n36), .B(n37), .Y(n34) );
  CLKINVX4 U53 ( .A(n3), .Y(SUM[6]) );
  NOR2BX2 U54 ( .AN(n65), .B(n27), .Y(n77) );
  NAND2X1 U55 ( .A(n37), .B(n210), .Y(n234) );
  NAND4BBX2 U56 ( .AN(n170), .BN(n176), .C(n174), .D(n175), .Y(n135) );
  INVX1 U57 ( .A(n253), .Y(n263) );
  INVX1 U58 ( .A(n35), .Y(n5) );
  NAND2X1 U59 ( .A(B[0]), .B(A[0]), .Y(n179) );
  INVX1 U60 ( .A(n137), .Y(n167) );
  INVX1 U61 ( .A(n131), .Y(n148) );
  NAND2X2 U62 ( .A(n140), .B(n149), .Y(n155) );
  NAND3X2 U63 ( .A(n163), .B(n162), .C(n145), .Y(n161) );
  AOI21X1 U64 ( .A0(n186), .A1(n174), .B0(n187), .Y(n185) );
  INVX1 U65 ( .A(n173), .Y(n187) );
  NAND2X2 U66 ( .A(n83), .B(n84), .Y(n75) );
  OR2X2 U67 ( .A(A[29]), .B(B[29]), .Y(n76) );
  NAND2X1 U68 ( .A(B[9]), .B(A[9]), .Y(n31) );
  CLKINVX3 U69 ( .A(n235), .Y(n32) );
  NOR2BX2 U70 ( .AN(n39), .B(n6), .Y(n33) );
  NOR2X2 U71 ( .A(A[2]), .B(B[2]), .Y(n27) );
  NAND2X1 U72 ( .A(B[2]), .B(A[2]), .Y(n65) );
  INVX1 U73 ( .A(n78), .Y(n178) );
  NOR2BX1 U74 ( .AN(n171), .B(n176), .Y(n222) );
  NOR2BX1 U75 ( .AN(n102), .B(n104), .Y(n124) );
  XOR2X2 U76 ( .A(n87), .B(n128), .Y(SUM[24]) );
  AND2X2 U77 ( .A(n173), .B(n174), .Y(n194) );
  INVX1 U78 ( .A(n186), .Y(n196) );
  NOR2BX1 U79 ( .AN(n70), .B(n23), .Y(n72) );
  NAND2X1 U80 ( .A(n197), .B(n172), .Y(n201) );
  INVX1 U81 ( .A(n171), .Y(n204) );
  NAND2X1 U82 ( .A(n210), .B(n9), .Y(n256) );
  XOR2X2 U83 ( .A(n283), .B(n285), .Y(SUM[10]) );
  NAND2X1 U84 ( .A(n35), .B(n36), .Y(n40) );
  NOR2BX1 U85 ( .AN(n54), .B(n59), .Y(n60) );
  NAND2X4 U86 ( .A(n146), .B(n147), .Y(n17) );
  AND2X4 U87 ( .A(n174), .B(n175), .Y(n25) );
  NAND2X1 U88 ( .A(B[23]), .B(A[23]), .Y(n2) );
  NAND2X1 U89 ( .A(B[20]), .B(A[20]), .Y(n145) );
  NAND2X1 U90 ( .A(B[6]), .B(A[6]), .Y(n45) );
  XNOR2X1 U91 ( .A(n46), .B(n47), .Y(n3) );
  OR2X2 U92 ( .A(n199), .B(n190), .Y(n4) );
  NAND2X1 U93 ( .A(B[15]), .B(A[15]), .Y(n192) );
  INVX1 U94 ( .A(n192), .Y(n199) );
  OR2X2 U95 ( .A(A[7]), .B(B[7]), .Y(n37) );
  NOR2X1 U96 ( .A(A[7]), .B(B[7]), .Y(n289) );
  NAND2X1 U97 ( .A(n198), .B(n197), .Y(n188) );
  OR2X2 U98 ( .A(n221), .B(n220), .Y(n217) );
  NAND2X4 U99 ( .A(n131), .B(n132), .Y(n142) );
  INVX3 U100 ( .A(n197), .Y(n170) );
  NAND2X2 U101 ( .A(B[17]), .B(A[17]), .Y(n172) );
  AOI21X2 U102 ( .A0(n154), .A1(n115), .B0(n155), .Y(n152) );
  AOI21X2 U103 ( .A0(n114), .A1(n115), .B0(n116), .Y(n120) );
  NAND2XL U104 ( .A(n114), .B(n115), .Y(n130) );
  XOR2X1 U105 ( .A(B[26]), .B(A[26]), .Y(n119) );
  NAND2X1 U106 ( .A(n258), .B(n248), .Y(n12) );
  AND2X2 U107 ( .A(n272), .B(n228), .Y(n258) );
  INVX4 U108 ( .A(n220), .Y(n228) );
  NOR3X4 U109 ( .A(n44), .B(n54), .C(n55), .Y(n300) );
  CLKINVX3 U110 ( .A(n1), .Y(n299) );
  NAND3BX4 U111 ( .AN(n48), .B(n49), .C(n50), .Y(n46) );
  AOI2BB2X4 U112 ( .B0(B[7]), .B1(A[7]), .A0N(n44), .A1N(n49), .Y(n297) );
  NAND2X1 U113 ( .A(B[5]), .B(A[5]), .Y(n49) );
  INVX8 U114 ( .A(n53), .Y(n58) );
  OAI2BB1XL U115 ( .A0N(n235), .A1N(n5), .B0(n31), .Y(n296) );
  INVX8 U116 ( .A(n290), .Y(n44) );
  INVX1 U117 ( .A(n111), .Y(n121) );
  OAI21X1 U118 ( .A0(n104), .A1(n101), .B0(n102), .Y(n111) );
  CLKINVX2 U119 ( .A(n249), .Y(n272) );
  NAND2XL U120 ( .A(n297), .B(n298), .Y(n6) );
  NOR2X4 U121 ( .A(n299), .B(n300), .Y(n298) );
  NOR2BX1 U122 ( .AN(n63), .B(n24), .Y(n62) );
  NOR2X4 U123 ( .A(A[3]), .B(B[3]), .Y(n24) );
  NAND2X2 U124 ( .A(B[3]), .B(A[3]), .Y(n63) );
  NOR3X2 U125 ( .A(n217), .B(n218), .C(n219), .Y(n205) );
  NAND2X2 U126 ( .A(n117), .B(n2), .Y(n116) );
  NAND2BX4 U127 ( .AN(n156), .B(n144), .Y(n149) );
  AOI21X2 U128 ( .A0(n88), .A1(n86), .B0(n89), .Y(n83) );
  INVX4 U129 ( .A(n91), .Y(n88) );
  AOI211X4 U130 ( .A0(n101), .A1(n102), .B0(n103), .C0(n104), .Y(n96) );
  INVX4 U131 ( .A(n106), .Y(n103) );
  NAND2X2 U132 ( .A(n210), .B(n211), .Y(n225) );
  NAND2X2 U133 ( .A(n263), .B(n255), .Y(n260) );
  NAND4X4 U134 ( .A(n21), .B(n211), .C(n231), .D(n232), .Y(n200) );
  OR2X4 U135 ( .A(n239), .B(n7), .Y(n21) );
  OR2X1 U136 ( .A(A[5]), .B(B[5]), .Y(n19) );
  NOR2X1 U137 ( .A(n269), .B(n249), .Y(n266) );
  INVX1 U138 ( .A(n87), .Y(n95) );
  XOR2X4 U139 ( .A(n92), .B(n93), .Y(SUM[28]) );
  OAI21X4 U140 ( .A0(n58), .A1(n59), .B0(n54), .Y(n56) );
  OAI21X2 U141 ( .A0(n170), .A1(n171), .B0(n172), .Y(n186) );
  XOR2X2 U142 ( .A(n66), .B(n77), .Y(SUM[2]) );
  OAI2BB1X2 U143 ( .A0N(n78), .A1N(n79), .B0(n80), .Y(n66) );
  AOI21X2 U144 ( .A0(B[13]), .A1(A[13]), .B0(n226), .Y(n224) );
  OR2X4 U145 ( .A(A[16]), .B(B[16]), .Y(n198) );
  NAND2X4 U146 ( .A(B[16]), .B(A[16]), .Y(n171) );
  NAND2X2 U147 ( .A(n279), .B(n282), .Y(n281) );
  OR2X4 U148 ( .A(A[27]), .B(B[27]), .Y(n98) );
  XOR2X4 U149 ( .A(n75), .B(n81), .Y(SUM[29]) );
  NOR2BX4 U150 ( .AN(n74), .B(n82), .Y(n81) );
  NOR2X2 U151 ( .A(n190), .B(n191), .Y(n223) );
  XOR2X4 U152 ( .A(n123), .B(n124), .Y(SUM[25]) );
  OAI2BB1X1 U153 ( .A0N(n160), .A1N(n115), .B0(n156), .Y(n158) );
  XOR2X4 U154 ( .A(n42), .B(n43), .Y(SUM[7]) );
  AND4X4 U155 ( .A(n131), .B(n132), .C(n133), .D(n134), .Y(n114) );
  AOI2BB1X2 U156 ( .A0N(n148), .A1N(n149), .B0(n150), .Y(n147) );
  NAND2X2 U157 ( .A(n235), .B(n36), .Y(n288) );
  AND2X4 U158 ( .A(n41), .B(n39), .Y(n22) );
  NAND2X1 U159 ( .A(n255), .B(n252), .Y(n264) );
  NAND2X1 U160 ( .A(B[13]), .B(A[13]), .Y(n252) );
  OR2X4 U161 ( .A(A[20]), .B(B[20]), .Y(n143) );
  INVX1 U162 ( .A(n198), .Y(n176) );
  NAND2X4 U163 ( .A(n286), .B(n287), .Y(n283) );
  NAND4BBX4 U164 ( .AN(n242), .BN(n32), .C(n237), .D(n238), .Y(n249) );
  AOI21X1 U165 ( .A0(n252), .A1(n213), .B0(n246), .Y(n250) );
  NOR2X2 U166 ( .A(n250), .B(n251), .Y(n244) );
  XOR2X2 U167 ( .A(n61), .B(n62), .Y(SUM[3]) );
  NOR2X2 U168 ( .A(A[13]), .B(B[13]), .Y(n28) );
  XOR2X2 U169 ( .A(n264), .B(n265), .Y(n303) );
  AOI21X2 U170 ( .A0(n266), .A1(n248), .B0(n267), .Y(n265) );
  BUFX8 U171 ( .A(n216), .Y(n9) );
  NAND2X1 U172 ( .A(n39), .B(n41), .Y(n273) );
  AOI21X4 U173 ( .A0(n224), .A1(n9), .B0(n225), .Y(n191) );
  OAI2BB1X1 U174 ( .A0N(B[2]), .A1N(A[2]), .B0(n80), .Y(n292) );
  NAND2X2 U175 ( .A(n163), .B(n168), .Y(n137) );
  NAND2X4 U176 ( .A(n25), .B(n169), .Y(n163) );
  XNOR2X4 U177 ( .A(n107), .B(n108), .Y(SUM[27]) );
  OAI21X2 U178 ( .A0(n120), .A1(n109), .B0(n110), .Y(n107) );
  NAND2X2 U179 ( .A(n161), .B(n143), .Y(n156) );
  OAI21X4 U180 ( .A0(n291), .A1(n292), .B0(n293), .Y(n240) );
  NAND2X1 U181 ( .A(n38), .B(n37), .Y(n41) );
  NAND4BX4 U182 ( .AN(n289), .B(n19), .C(n290), .D(n52), .Y(n241) );
  XOR2X2 U183 ( .A(n79), .B(n177), .Y(SUM[1]) );
  NOR4X2 U184 ( .A(n189), .B(n199), .C(n190), .D(n191), .Y(n183) );
  CLKINVX3 U185 ( .A(n151), .Y(n160) );
  INVX4 U186 ( .A(n51), .Y(n55) );
  XOR2X4 U187 ( .A(n164), .B(n165), .Y(SUM[20]) );
  OAI21X2 U188 ( .A0(n64), .A1(n27), .B0(n65), .Y(n61) );
  NAND2X4 U189 ( .A(B[18]), .B(A[18]), .Y(n173) );
  XOR2X4 U190 ( .A(n67), .B(n68), .Y(SUM[31]) );
  OAI21X4 U191 ( .A0(n23), .A1(n69), .B0(n70), .Y(n67) );
  OAI2BB1X1 U192 ( .A0N(n46), .A1N(n290), .B0(n1), .Y(n42) );
  CLKINVX4 U193 ( .A(n200), .Y(n189) );
  AND2X4 U194 ( .A(n12), .B(n13), .Y(n257) );
  OAI21X2 U195 ( .A0(n219), .A1(n260), .B0(n261), .Y(n259) );
  INVX4 U196 ( .A(n52), .Y(n59) );
  NAND3X2 U197 ( .A(n51), .B(n52), .C(n53), .Y(n50) );
  OR2X4 U198 ( .A(A[4]), .B(B[4]), .Y(n52) );
  NAND2X2 U199 ( .A(B[24]), .B(A[24]), .Y(n101) );
  NAND2X1 U200 ( .A(B[10]), .B(A[10]), .Y(n279) );
  INVX2 U201 ( .A(n66), .Y(n64) );
  NAND2X4 U202 ( .A(n63), .B(n240), .Y(n53) );
  NOR2X4 U203 ( .A(n24), .B(n27), .Y(n293) );
  XOR2X4 U204 ( .A(n180), .B(n181), .Y(SUM[19]) );
  NOR2BX1 U205 ( .AN(n80), .B(n178), .Y(n177) );
  NOR2XL U206 ( .A(n54), .B(n55), .Y(n48) );
  NAND2X2 U207 ( .A(n283), .B(n237), .Y(n282) );
  AND4X4 U208 ( .A(n227), .B(n228), .C(n211), .D(n229), .Y(n190) );
  OR2X4 U209 ( .A(A[8]), .B(B[8]), .Y(n36) );
  XOR2X4 U210 ( .A(n17), .B(n18), .Y(SUM[23]) );
  OAI21X2 U211 ( .A0(n125), .A1(n126), .B0(n101), .Y(n123) );
  OAI21X4 U212 ( .A0(n33), .A1(n34), .B0(n35), .Y(n29) );
  NAND2XL U213 ( .A(n213), .B(n247), .Y(n271) );
  AOI2BB1X1 U214 ( .A0N(n28), .A1N(n213), .B0(n262), .Y(n261) );
  INVXL U215 ( .A(n9), .Y(n251) );
  OAI21X2 U216 ( .A0(n120), .A1(n113), .B0(n121), .Y(n118) );
  AND2X1 U217 ( .A(n132), .B(n2), .Y(n18) );
  AND3X4 U218 ( .A(n192), .B(n200), .C(n223), .Y(n26) );
  INVX8 U219 ( .A(n26), .Y(n115) );
  NAND2X2 U220 ( .A(B[12]), .B(A[12]), .Y(n213) );
  INVXL U221 ( .A(A[13]), .Y(n214) );
  NAND2XL U222 ( .A(B[26]), .B(A[26]), .Y(n100) );
  XOR2X2 U223 ( .A(n115), .B(n222), .Y(n302) );
  INVX4 U224 ( .A(n122), .Y(n104) );
  INVXL U225 ( .A(n86), .Y(n94) );
  XOR2X4 U226 ( .A(n15), .B(n16), .Y(SUM[15]) );
  AOI21X2 U227 ( .A0(n114), .A1(n115), .B0(n127), .Y(n126) );
  XNOR2X4 U228 ( .A(n270), .B(n271), .Y(SUM[12]) );
  NAND2X2 U229 ( .A(n73), .B(n74), .Y(n71) );
  INVXL U230 ( .A(n144), .Y(n157) );
  INVXL U231 ( .A(n143), .Y(n166) );
  AOI21XL U232 ( .A0(B[7]), .A1(A[7]), .B0(n289), .Y(n43) );
  NAND2XL U233 ( .A(n99), .B(n98), .Y(n108) );
  OR2X4 U234 ( .A(A[12]), .B(B[12]), .Y(n247) );
  OR2X4 U235 ( .A(A[15]), .B(B[15]), .Y(n211) );
  AOI21XL U236 ( .A0(n63), .A1(n240), .B0(n241), .Y(n239) );
  OAI21XL U237 ( .A0(n140), .A1(n148), .B0(n141), .Y(n150) );
  OR2X4 U238 ( .A(A[23]), .B(B[23]), .Y(n132) );
  NOR2BX1 U239 ( .AN(n9), .B(n212), .Y(n208) );
  OR2X4 U240 ( .A(A[18]), .B(B[18]), .Y(n174) );
  OR2X4 U241 ( .A(A[26]), .B(B[26]), .Y(n106) );
  NOR2BX1 U242 ( .AN(n179), .B(n20), .Y(SUM[0]) );
  NOR2XL U243 ( .A(A[0]), .B(B[0]), .Y(n20) );
  INVX1 U244 ( .A(n71), .Y(n69) );
  XOR2X1 U245 ( .A(n71), .B(n72), .Y(n301) );
  INVX1 U246 ( .A(n36), .Y(n242) );
  INVX1 U247 ( .A(n76), .Y(n82) );
  NOR2BX1 U248 ( .AN(n101), .B(n125), .Y(n128) );
  NOR2BX1 U249 ( .AN(n90), .B(n94), .Y(n93) );
  NOR2BX1 U250 ( .AN(n140), .B(n157), .Y(n159) );
  NOR2BX1 U251 ( .AN(n145), .B(n166), .Y(n165) );
  OAI2BB1X1 U252 ( .A0N(n134), .A1N(n115), .B0(n167), .Y(n164) );
  XOR2X1 U253 ( .A(n53), .B(n60), .Y(SUM[4]) );
  XOR2X4 U254 ( .A(n40), .B(n22), .Y(SUM[8]) );
  NOR2BXL U255 ( .AN(n279), .B(n277), .Y(n285) );
  OAI2BB1X2 U256 ( .A0N(n272), .A1N(n273), .B0(n274), .Y(n270) );
  INVX1 U257 ( .A(n105), .Y(n125) );
  NAND3BXL U258 ( .AN(n253), .B(n254), .C(n229), .Y(n243) );
  INVX1 U259 ( .A(n246), .Y(n254) );
  INVX1 U260 ( .A(n90), .Y(n89) );
  INVX1 U261 ( .A(n247), .Y(n269) );
  INVX1 U262 ( .A(n211), .Y(n218) );
  NAND2XL U263 ( .A(n36), .B(n235), .Y(n233) );
  NAND2XL U264 ( .A(n230), .B(n229), .Y(n274) );
  NAND2XL U265 ( .A(n237), .B(n238), .Y(n236) );
  NAND2X1 U266 ( .A(n75), .B(n76), .Y(n73) );
  INVX1 U267 ( .A(n221), .Y(n227) );
  OAI2BB1X2 U268 ( .A0N(B[11]), .A1N(A[11]), .B0(n279), .Y(n275) );
  NAND3X1 U269 ( .A(n145), .B(n140), .C(n141), .Y(n138) );
  NAND2X1 U270 ( .A(B[21]), .B(A[21]), .Y(n140) );
  CLKINVX3 U271 ( .A(n136), .Y(n133) );
  OR2X2 U272 ( .A(A[21]), .B(B[21]), .Y(n144) );
  NAND2XL U273 ( .A(n141), .B(n131), .Y(n153) );
  NAND2XL U274 ( .A(n230), .B(n284), .Y(n280) );
  NAND2XL U275 ( .A(B[11]), .B(A[11]), .Y(n284) );
  NOR2BXL U276 ( .AN(n1), .B(n44), .Y(n47) );
  XOR2X2 U277 ( .A(n56), .B(n57), .Y(SUM[5]) );
  NAND2XL U278 ( .A(n2), .B(n117), .Y(n129) );
  NAND2X1 U279 ( .A(B[25]), .B(A[25]), .Y(n102) );
  NOR2X1 U280 ( .A(A[30]), .B(B[30]), .Y(n23) );
  INVX1 U281 ( .A(n100), .Y(n112) );
  NAND2XL U282 ( .A(B[19]), .B(A[19]), .Y(n168) );
  OR2X2 U283 ( .A(A[11]), .B(B[11]), .Y(n238) );
  NAND2XL U284 ( .A(B[19]), .B(A[19]), .Y(n162) );
  NAND2XL U285 ( .A(n210), .B(n211), .Y(n209) );
  INVX1 U286 ( .A(n179), .Y(n79) );
  NAND2X1 U287 ( .A(n117), .B(n2), .Y(n127) );
  NAND2BX1 U288 ( .AN(n188), .B(n174), .Y(n184) );
  NAND2BX1 U289 ( .AN(n113), .B(n106), .Y(n109) );
  OR2X2 U290 ( .A(A[25]), .B(B[25]), .Y(n122) );
  INVX1 U291 ( .A(n252), .Y(n262) );
  INVXL U292 ( .A(B[13]), .Y(n215) );
  OR2X2 U293 ( .A(A[28]), .B(B[28]), .Y(n86) );
  NAND2X1 U294 ( .A(B[29]), .B(A[29]), .Y(n74) );
  NAND2X1 U295 ( .A(B[30]), .B(A[30]), .Y(n70) );
  NAND2X1 U296 ( .A(B[28]), .B(A[28]), .Y(n90) );
  NOR2X1 U297 ( .A(n28), .B(n213), .Y(n226) );
  NOR2X2 U298 ( .A(n178), .B(n294), .Y(n291) );
  NAND2X1 U299 ( .A(B[14]), .B(A[14]), .Y(n216) );
  XOR2X1 U300 ( .A(B[31]), .B(A[31]), .Y(n68) );
  NAND2X1 U301 ( .A(B[1]), .B(A[1]), .Y(n80) );
  OAI22X1 U302 ( .A0(n28), .A1(n213), .B0(n214), .B1(n215), .Y(n212) );
  NAND2X1 U303 ( .A(A[0]), .B(B[0]), .Y(n294) );
  XOR2X4 U304 ( .A(n29), .B(n30), .Y(SUM[9]) );
  XOR2X4 U305 ( .A(n118), .B(n119), .Y(SUM[26]) );
  NAND2BX4 U306 ( .AN(n129), .B(n130), .Y(n87) );
  OAI21X4 U307 ( .A0(n137), .A1(n138), .B0(n139), .Y(n117) );
  AOI31X2 U308 ( .A0(n136), .A1(n140), .A2(n141), .B0(n142), .Y(n139) );
  OR2X4 U309 ( .A(A[22]), .B(B[22]), .Y(n131) );
  XOR2X4 U310 ( .A(n158), .B(n159), .Y(SUM[21]) );
  OAI211X2 U311 ( .A0(n170), .A1(n171), .B0(n172), .C0(n173), .Y(n169) );
  NOR2BX4 U312 ( .AN(n168), .B(n182), .Y(n181) );
  OR2X4 U313 ( .A(A[19]), .B(B[19]), .Y(n175) );
  XOR2X4 U314 ( .A(n193), .B(n194), .Y(SUM[18]) );
  XOR2X4 U315 ( .A(n201), .B(n202), .Y(SUM[17]) );
  AOI21X4 U316 ( .A0(n203), .A1(n198), .B0(n204), .Y(n202) );
  OR2X4 U317 ( .A(A[17]), .B(B[17]), .Y(n197) );
  NOR2X4 U318 ( .A(n233), .B(n234), .Y(n232) );
  NOR2X4 U319 ( .A(n220), .B(n236), .Y(n231) );
  XOR2X4 U320 ( .A(n256), .B(n257), .Y(SUM[14]) );
  OR2X4 U321 ( .A(A[14]), .B(B[14]), .Y(n210) );
  OAI21X4 U322 ( .A0(n58), .A1(n241), .B0(n268), .Y(n248) );
  NAND2X4 U323 ( .A(n7), .B(n37), .Y(n268) );
  OR2X4 U324 ( .A(A[13]), .B(B[13]), .Y(n255) );
  NAND2BX4 U325 ( .AN(n275), .B(n276), .Y(n229) );
  NAND3BX4 U326 ( .AN(n277), .B(n235), .C(n278), .Y(n276) );
  OR2X4 U327 ( .A(A[10]), .B(B[10]), .Y(n237) );
  NAND2X4 U328 ( .A(B[8]), .B(A[8]), .Y(n35) );
  NAND2X4 U329 ( .A(n297), .B(n298), .Y(n38) );
  OR2X4 U330 ( .A(A[5]), .B(B[5]), .Y(n51) );
  OR2X4 U331 ( .A(A[6]), .B(B[6]), .Y(n290) );
  OR2X4 U332 ( .A(A[9]), .B(B[9]), .Y(n235) );
endmodule


module hash_core_DW01_add_26 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n300, n301, n302, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299;

  NAND2X4 U2 ( .A(n53), .B(A[28]), .Y(n129) );
  BUFX3 U3 ( .A(B[28]), .Y(n53) );
  BUFX4 U4 ( .A(n219), .Y(n47) );
  NAND2X2 U5 ( .A(n18), .B(n223), .Y(n229) );
  BUFX3 U6 ( .A(n221), .Y(n18) );
  BUFX20 U7 ( .A(n300), .Y(SUM[18]) );
  NOR2X2 U8 ( .A(n283), .B(n282), .Y(n48) );
  NAND3BX4 U9 ( .AN(n167), .B(n165), .C(n156), .Y(n161) );
  OR2XL U10 ( .A(n219), .B(n20), .Y(n55) );
  CLKINVX3 U11 ( .A(n208), .Y(n184) );
  NOR2X4 U12 ( .A(B[17]), .B(A[17]), .Y(n217) );
  CLKINVX3 U13 ( .A(n175), .Y(n179) );
  INVX8 U14 ( .A(n38), .Y(n39) );
  NOR2X4 U15 ( .A(n143), .B(n32), .Y(n146) );
  XOR2X2 U16 ( .A(n95), .B(n96), .Y(n301) );
  CLKINVX3 U17 ( .A(n271), .Y(n24) );
  NAND3X2 U18 ( .A(n265), .B(n269), .C(n12), .Y(n271) );
  NAND2X2 U19 ( .A(n79), .B(A[19]), .Y(n203) );
  BUFX12 U20 ( .A(n200), .Y(n75) );
  NAND2X4 U21 ( .A(n74), .B(n144), .Y(n3) );
  BUFX20 U22 ( .A(n145), .Y(n74) );
  NAND3BX4 U23 ( .AN(n123), .B(n125), .C(n124), .Y(n117) );
  NAND2X4 U24 ( .A(B[5]), .B(A[5]), .Y(n100) );
  INVX12 U25 ( .A(n97), .Y(n93) );
  NAND2X4 U26 ( .A(n100), .B(n104), .Y(n294) );
  NAND2X4 U27 ( .A(B[21]), .B(A[21]), .Y(n191) );
  NAND2BX4 U28 ( .AN(n198), .B(n4), .Y(n196) );
  NAND2X4 U29 ( .A(n144), .B(n74), .Y(n165) );
  OR2X4 U30 ( .A(A[19]), .B(n79), .Y(n199) );
  BUFX8 U31 ( .A(B[19]), .Y(n79) );
  AND3X2 U32 ( .A(n221), .B(n222), .C(n223), .Y(n16) );
  OR2X4 U33 ( .A(B[18]), .B(A[18]), .Y(n223) );
  AND2X4 U34 ( .A(n202), .B(n203), .Y(n212) );
  OAI21X4 U35 ( .A0(n15), .A1(n190), .B0(n191), .Y(n187) );
  INVX8 U36 ( .A(n166), .Y(n144) );
  BUFX4 U37 ( .A(n65), .Y(n1) );
  NAND2X4 U38 ( .A(n113), .B(n135), .Y(n299) );
  NOR2BX1 U39 ( .AN(n231), .B(n20), .Y(n233) );
  INVX4 U40 ( .A(n231), .Y(n213) );
  NOR2X4 U41 ( .A(B[18]), .B(A[18]), .Y(n20) );
  XOR2X2 U42 ( .A(n134), .B(n224), .Y(SUM[1]) );
  XOR2X2 U43 ( .A(n28), .B(n85), .Y(SUM[8]) );
  NAND2X1 U44 ( .A(B[30]), .B(A[30]), .Y(n120) );
  NAND2X2 U45 ( .A(B[0]), .B(A[0]), .Y(n226) );
  AND2X2 U46 ( .A(n268), .B(n269), .Y(n266) );
  NAND2X1 U47 ( .A(A[12]), .B(B[12]), .Y(n269) );
  NAND2X2 U48 ( .A(A[16]), .B(B[16]), .Y(n218) );
  NOR2X2 U49 ( .A(A[4]), .B(B[4]), .Y(n68) );
  OR2X4 U50 ( .A(A[30]), .B(B[30]), .Y(n118) );
  NOR2BX4 U51 ( .AN(n124), .B(n130), .Y(n137) );
  INVX4 U52 ( .A(n127), .Y(n130) );
  XOR2X2 U53 ( .A(n114), .B(n131), .Y(SUM[2]) );
  NOR2BX4 U54 ( .AN(n64), .B(n26), .Y(n290) );
  NAND2X2 U55 ( .A(n64), .B(n288), .Y(n286) );
  NAND2X4 U56 ( .A(B[10]), .B(A[10]), .Y(n64) );
  NOR2X2 U57 ( .A(n298), .B(n299), .Y(n296) );
  NOR2X4 U58 ( .A(n225), .B(n226), .Y(n298) );
  CLKINVX8 U59 ( .A(n34), .Y(n25) );
  NOR2X4 U60 ( .A(B[10]), .B(A[10]), .Y(n34) );
  BUFX8 U61 ( .A(n302), .Y(SUM[4]) );
  XOR2X2 U62 ( .A(n23), .B(n106), .Y(n302) );
  CLKINVX4 U63 ( .A(n3), .Y(n180) );
  INVX1 U64 ( .A(A[17]), .Y(n5) );
  NOR2X2 U65 ( .A(n68), .B(n103), .Y(n62) );
  INVXL U66 ( .A(n22), .Y(n90) );
  INVXL U67 ( .A(n198), .Y(n17) );
  AND2X2 U68 ( .A(n235), .B(n222), .Y(n239) );
  INVX1 U69 ( .A(n268), .Y(n272) );
  NAND2X2 U70 ( .A(n82), .B(n86), .Y(n279) );
  INVX1 U71 ( .A(n13), .Y(n4) );
  NAND2X1 U72 ( .A(n25), .B(n289), .Y(n288) );
  INVX1 U73 ( .A(n115), .Y(n58) );
  NOR2X2 U74 ( .A(n129), .B(n130), .Y(n123) );
  NOR2BX1 U75 ( .AN(n157), .B(n151), .Y(n160) );
  CLKINVX3 U76 ( .A(n98), .Y(n102) );
  CLKINVX3 U77 ( .A(n95), .Y(n92) );
  NAND2X1 U78 ( .A(B[16]), .B(A[16]), .Y(n235) );
  AOI31X1 U79 ( .A0(n265), .A1(n266), .A2(n12), .B0(n267), .Y(n264) );
  NOR2BX2 U80 ( .AN(n129), .B(n138), .Y(n139) );
  XOR2X2 U81 ( .A(n99), .B(n101), .Y(SUM[5]) );
  NOR2BX1 U82 ( .AN(n100), .B(n102), .Y(n101) );
  NOR2BX1 U83 ( .AN(n82), .B(n83), .Y(n81) );
  AND2X2 U84 ( .A(n86), .B(n87), .Y(n85) );
  CLKBUFX3 U85 ( .A(n19), .Y(n28) );
  NOR2BX1 U86 ( .AN(n94), .B(n93), .Y(n96) );
  NAND2X2 U87 ( .A(B[6]), .B(A[6]), .Y(n94) );
  CLKINVX3 U88 ( .A(n154), .Y(n153) );
  NAND2X2 U89 ( .A(n74), .B(n144), .Y(n181) );
  INVX1 U90 ( .A(n18), .Y(n234) );
  OR2XL U91 ( .A(A[21]), .B(B[21]), .Y(n78) );
  OAI2BB1X2 U92 ( .A0N(n190), .A1N(n191), .B0(n78), .Y(n197) );
  CLKINVX3 U93 ( .A(n235), .Y(n238) );
  NAND2BX4 U94 ( .AN(n5), .B(B[17]), .Y(n219) );
  NAND3X2 U95 ( .A(n171), .B(n144), .C(n74), .Y(n170) );
  NAND2X4 U96 ( .A(n249), .B(n84), .Y(n6) );
  NAND2X4 U97 ( .A(n7), .B(n41), .Y(n241) );
  INVX4 U98 ( .A(n6), .Y(n7) );
  OAI21X4 U99 ( .A0(n103), .A1(n250), .B0(n251), .Y(n84) );
  BUFX3 U100 ( .A(n147), .Y(n37) );
  NAND2X4 U101 ( .A(n170), .B(n169), .Y(n168) );
  INVX1 U102 ( .A(n25), .Y(n26) );
  INVX4 U103 ( .A(n274), .Y(n248) );
  AND2X2 U104 ( .A(B[14]), .B(A[14]), .Y(n27) );
  AND2X2 U105 ( .A(n174), .B(n186), .Y(n8) );
  AND2X2 U106 ( .A(n49), .B(n150), .Y(n9) );
  AND2X2 U107 ( .A(B[22]), .B(A[22]), .Y(n10) );
  AND2X2 U108 ( .A(n126), .B(n127), .Y(n11) );
  NAND3X2 U109 ( .A(n246), .B(n274), .C(n249), .Y(n12) );
  INVX2 U110 ( .A(n75), .Y(n38) );
  AOI21X4 U111 ( .A0(n16), .A1(n39), .B0(n201), .Y(n195) );
  INVX1 U112 ( .A(n199), .Y(n13) );
  NOR2BX4 U113 ( .AN(n14), .B(B[21]), .Y(n15) );
  INVX1 U114 ( .A(A[21]), .Y(n14) );
  BUFX8 U115 ( .A(n301), .Y(SUM[6]) );
  INVX4 U116 ( .A(n43), .Y(n276) );
  NAND4BX4 U117 ( .AN(n143), .B(n171), .C(n144), .D(n46), .Y(n142) );
  XOR2X4 U118 ( .A(n289), .B(n290), .Y(SUM[10]) );
  OR2X4 U119 ( .A(A[27]), .B(B[27]), .Y(n42) );
  OAI2BB1X4 U120 ( .A0N(n17), .A1N(n74), .B0(n197), .Y(n205) );
  NOR3X4 U121 ( .A(n143), .B(n173), .C(n156), .Y(n152) );
  OAI21X4 U122 ( .A0(n103), .A1(n250), .B0(n251), .Y(n19) );
  XNOR2X4 U123 ( .A(n24), .B(n273), .Y(SUM[13]) );
  XNOR2X4 U124 ( .A(n74), .B(n21), .Y(SUM[20]) );
  NAND2XL U125 ( .A(n190), .B(n208), .Y(n21) );
  INVX1 U126 ( .A(n27), .Y(n260) );
  NOR2BX4 U127 ( .AN(n94), .B(n22), .Y(n292) );
  OAI2BB1X4 U128 ( .A0N(n98), .A1N(n99), .B0(n100), .Y(n95) );
  AND2X4 U129 ( .A(B[7]), .B(A[7]), .Y(n22) );
  INVXL U130 ( .A(n103), .Y(n23) );
  CLKBUFXL U131 ( .A(n48), .Y(n29) );
  INVX2 U132 ( .A(n171), .Y(n32) );
  NAND2X4 U133 ( .A(n11), .B(n128), .Y(n125) );
  BUFX8 U134 ( .A(B[11]), .Y(n30) );
  CLKINVX4 U135 ( .A(n157), .Y(n164) );
  OAI21X4 U136 ( .A0(n187), .A1(n10), .B0(n188), .Y(n31) );
  INVXL U137 ( .A(n35), .Y(n33) );
  NOR2X4 U138 ( .A(A[15]), .B(B[15]), .Y(n35) );
  NOR2BX1 U139 ( .AN(n191), .B(n15), .Y(n210) );
  OR2X2 U140 ( .A(A[21]), .B(B[21]), .Y(n77) );
  AOI21X4 U141 ( .A0(n30), .A1(A[11]), .B0(n281), .Y(n280) );
  INVX4 U142 ( .A(n155), .Y(n173) );
  NAND2X4 U143 ( .A(n57), .B(n31), .Y(n147) );
  NAND2X1 U144 ( .A(A[15]), .B(B[15]), .Y(n257) );
  NAND3X4 U145 ( .A(n98), .B(n97), .C(n294), .Y(n293) );
  INVX8 U146 ( .A(n151), .Y(n171) );
  INVXL U147 ( .A(B[13]), .Y(n261) );
  NAND2BX2 U148 ( .AN(A[13]), .B(n261), .Y(n259) );
  NAND2XL U149 ( .A(n202), .B(n203), .Y(n201) );
  INVXL U150 ( .A(n247), .Y(n36) );
  NAND2X2 U151 ( .A(B[8]), .B(A[8]), .Y(n86) );
  INVX8 U152 ( .A(n284), .Y(n83) );
  INVX8 U153 ( .A(n70), .Y(SUM[11]) );
  XNOR2X4 U154 ( .A(n286), .B(n71), .Y(n70) );
  NOR2BX2 U155 ( .AN(n260), .B(n264), .Y(n263) );
  NOR2X4 U156 ( .A(B[14]), .B(A[14]), .Y(n40) );
  NAND2X2 U157 ( .A(B[18]), .B(A[18]), .Y(n231) );
  AND4X4 U158 ( .A(n255), .B(n254), .C(n253), .D(n252), .Y(n41) );
  XOR2X2 U159 ( .A(n80), .B(n81), .Y(SUM[9]) );
  OAI2BB1X2 U160 ( .A0N(n29), .A1N(n28), .B0(n44), .Y(n43) );
  OR2X2 U161 ( .A(n277), .B(n248), .Y(n44) );
  NAND2X2 U162 ( .A(B[9]), .B(A[9]), .Y(n82) );
  AND2X2 U163 ( .A(n154), .B(n158), .Y(n45) );
  NAND2X1 U164 ( .A(A[23]), .B(B[23]), .Y(n174) );
  CLKINVX4 U165 ( .A(n207), .Y(n46) );
  INVX8 U166 ( .A(n74), .Y(n207) );
  NAND2X1 U167 ( .A(n47), .B(n221), .Y(n236) );
  INVX3 U168 ( .A(n116), .Y(n59) );
  NAND3BX2 U169 ( .AN(n243), .B(n84), .C(n48), .Y(n265) );
  OR2X4 U170 ( .A(A[26]), .B(B[26]), .Y(n49) );
  AND3X4 U171 ( .A(n141), .B(n142), .C(n140), .Y(n50) );
  NAND3BX4 U172 ( .AN(n123), .B(n125), .C(n124), .Y(n51) );
  NOR2X4 U173 ( .A(n152), .B(n153), .Y(n140) );
  NAND2X2 U174 ( .A(B[29]), .B(A[29]), .Y(n124) );
  INVX4 U175 ( .A(n64), .Y(n281) );
  NAND2XL U176 ( .A(A[11]), .B(n30), .Y(n287) );
  OAI2BB1X4 U177 ( .A0N(n279), .A1N(n278), .B0(n280), .Y(n52) );
  AND2X4 U178 ( .A(A[13]), .B(B[13]), .Y(n72) );
  XOR2X4 U179 ( .A(n128), .B(n139), .Y(SUM[28]) );
  NAND2X4 U180 ( .A(n49), .B(n42), .Y(n54) );
  AND2X2 U181 ( .A(n231), .B(n55), .Y(n230) );
  NOR2X4 U182 ( .A(n247), .B(n40), .Y(n245) );
  INVX4 U183 ( .A(n252), .Y(n247) );
  NAND2X4 U184 ( .A(n87), .B(n19), .Y(n291) );
  OR2X4 U185 ( .A(A[11]), .B(B[11]), .Y(n274) );
  NAND4BX4 U186 ( .AN(n243), .B(n244), .C(n52), .D(n245), .Y(n242) );
  INVX3 U187 ( .A(n249), .Y(n243) );
  NAND2X1 U188 ( .A(A[27]), .B(B[27]), .Y(n154) );
  BUFX2 U189 ( .A(n174), .Y(n57) );
  OAI2BB1X4 U190 ( .A0N(n80), .A1N(n284), .B0(n82), .Y(n289) );
  INVX8 U191 ( .A(n105), .Y(n103) );
  NAND2BX2 U192 ( .AN(n167), .B(n181), .Y(n182) );
  NAND2X1 U193 ( .A(B[3]), .B(A[3]), .Y(n109) );
  OAI2BB1X4 U194 ( .A0N(n292), .A1N(n293), .B0(n91), .Y(n251) );
  NAND2X2 U195 ( .A(n58), .B(n116), .Y(n61) );
  NOR2BX2 U196 ( .AN(n156), .B(n179), .Y(n183) );
  NAND2X4 U197 ( .A(n115), .B(n59), .Y(n60) );
  NAND2X4 U198 ( .A(n60), .B(n61), .Y(SUM[31]) );
  XNOR2X4 U199 ( .A(B[31]), .B(A[31]), .Y(n115) );
  AOI21X4 U200 ( .A0(n117), .A1(n118), .B0(n119), .Y(n116) );
  INVX8 U201 ( .A(n69), .Y(SUM[25]) );
  NAND2X4 U202 ( .A(n208), .B(n77), .Y(n198) );
  OR2X4 U203 ( .A(n62), .B(n63), .Y(n99) );
  INVXL U204 ( .A(n104), .Y(n63) );
  AOI21X4 U205 ( .A0(n146), .A1(n37), .B0(n148), .Y(n141) );
  NOR2BX1 U206 ( .AN(n113), .B(n112), .Y(n131) );
  AND2X1 U207 ( .A(n203), .B(n216), .Y(n66) );
  AND2X1 U208 ( .A(n274), .B(n287), .Y(n71) );
  OAI21X4 U209 ( .A0(n217), .A1(n218), .B0(n219), .Y(n214) );
  NOR2BX4 U210 ( .AN(n216), .B(n20), .Y(n215) );
  NOR2XL U211 ( .A(A[0]), .B(B[0]), .Y(n67) );
  NAND2X2 U212 ( .A(B[26]), .B(A[26]), .Y(n150) );
  CLKINVX3 U213 ( .A(n226), .Y(n134) );
  AND2X1 U214 ( .A(n90), .B(n91), .Y(n89) );
  NOR2X4 U215 ( .A(n35), .B(n248), .Y(n244) );
  NAND2X4 U216 ( .A(B[2]), .B(A[2]), .Y(n113) );
  NAND2X4 U217 ( .A(B[4]), .B(A[4]), .Y(n104) );
  AOI21X4 U218 ( .A0(n75), .A1(n222), .B0(n238), .Y(n228) );
  XOR2X4 U219 ( .A(n270), .B(n1), .Y(SUM[14]) );
  NAND2XL U220 ( .A(n260), .B(n254), .Y(n65) );
  XOR2X4 U221 ( .A(n227), .B(n66), .Y(SUM[19]) );
  XNOR2X4 U222 ( .A(n176), .B(n177), .Y(n69) );
  NOR2BX1 U223 ( .AN(n226), .B(n67), .Y(SUM[0]) );
  INVX1 U224 ( .A(n114), .Y(n111) );
  XOR2X1 U225 ( .A(n107), .B(n108), .Y(SUM[3]) );
  NOR2BX1 U226 ( .AN(n109), .B(n110), .Y(n108) );
  OAI21XL U227 ( .A0(n111), .A1(n112), .B0(n113), .Y(n107) );
  INVXL U228 ( .A(n295), .Y(n110) );
  NOR2BXL U229 ( .AN(n135), .B(n225), .Y(n224) );
  INVXL U230 ( .A(n132), .Y(n112) );
  NOR2BX1 U231 ( .AN(n104), .B(n68), .Y(n106) );
  OAI2BB1X1 U232 ( .A0N(n133), .A1N(n134), .B0(n135), .Y(n114) );
  NAND2XL U233 ( .A(n269), .B(n249), .Y(n275) );
  NOR2BXL U234 ( .AN(n268), .B(n247), .Y(n273) );
  NOR2BX1 U235 ( .AN(n194), .B(n189), .Y(n206) );
  NAND2XL U236 ( .A(n257), .B(n33), .Y(n262) );
  INVXL U237 ( .A(n246), .Y(n277) );
  NAND2X2 U238 ( .A(B[1]), .B(A[1]), .Y(n135) );
  INVX1 U239 ( .A(n120), .Y(n119) );
  NAND2X2 U240 ( .A(B[20]), .B(A[20]), .Y(n190) );
  AOI2BB1X4 U241 ( .A0N(n72), .A1N(n73), .B0(n40), .Y(n258) );
  AND2X4 U242 ( .A(B[12]), .B(A[12]), .Y(n73) );
  NAND2X2 U243 ( .A(B[24]), .B(A[24]), .Y(n156) );
  NAND2X2 U244 ( .A(B[25]), .B(A[25]), .Y(n149) );
  NAND2XL U245 ( .A(A[13]), .B(B[13]), .Y(n268) );
  NAND2XL U246 ( .A(B[22]), .B(A[22]), .Y(n194) );
  NAND3BX4 U247 ( .AN(n240), .B(n242), .C(n241), .Y(n200) );
  NAND2XL U248 ( .A(n252), .B(n254), .Y(n267) );
  OAI21X4 U249 ( .A0(n207), .A1(n184), .B0(n190), .Y(n209) );
  OAI21X4 U250 ( .A0(n237), .A1(n234), .B0(n47), .Y(n232) );
  XOR2X4 U251 ( .A(n88), .B(n89), .Y(SUM[7]) );
  OAI21X4 U252 ( .A0(n92), .A1(n93), .B0(n94), .Y(n88) );
  XOR2X4 U253 ( .A(n51), .B(n121), .Y(SUM[30]) );
  NOR2BX4 U254 ( .AN(n120), .B(n122), .Y(n121) );
  CLKINVX3 U255 ( .A(n118), .Y(n122) );
  XOR2X4 U256 ( .A(n136), .B(n137), .Y(SUM[29]) );
  OR2X4 U257 ( .A(A[29]), .B(B[29]), .Y(n127) );
  OAI21X4 U258 ( .A0(n50), .A1(n138), .B0(n129), .Y(n136) );
  CLKINVX3 U259 ( .A(n126), .Y(n138) );
  OR2X4 U260 ( .A(A[28]), .B(B[28]), .Y(n126) );
  NAND3X4 U261 ( .A(n142), .B(n141), .C(n140), .Y(n128) );
  OAI22X4 U262 ( .A0(n54), .A1(n149), .B0(n54), .B1(n150), .Y(n148) );
  NAND2X4 U263 ( .A(n49), .B(n158), .Y(n143) );
  XOR2X4 U264 ( .A(n159), .B(n45), .Y(SUM[27]) );
  OR2X4 U265 ( .A(B[27]), .B(A[27]), .Y(n158) );
  OAI2BB1X4 U266 ( .A0N(n160), .A1N(n161), .B0(n162), .Y(n159) );
  NOR2BX4 U267 ( .AN(n150), .B(n163), .Y(n162) );
  NOR2X4 U268 ( .A(n149), .B(n164), .Y(n163) );
  XOR2X4 U269 ( .A(n168), .B(n9), .Y(SUM[26]) );
  OR2X4 U270 ( .A(A[26]), .B(B[26]), .Y(n157) );
  AOI21X4 U271 ( .A0(n147), .A1(n171), .B0(n172), .Y(n169) );
  OAI21X4 U272 ( .A0(n173), .A1(n156), .B0(n149), .Y(n172) );
  NAND2X4 U273 ( .A(n175), .B(n155), .Y(n151) );
  NOR2BX4 U274 ( .AN(n149), .B(n173), .Y(n177) );
  OR2X4 U275 ( .A(B[25]), .B(A[25]), .Y(n155) );
  OAI21X4 U276 ( .A0(n178), .A1(n179), .B0(n156), .Y(n176) );
  NOR2X4 U277 ( .A(n180), .B(n147), .Y(n178) );
  XOR2X4 U278 ( .A(n182), .B(n183), .Y(SUM[24]) );
  OR2X4 U279 ( .A(A[24]), .B(B[24]), .Y(n175) );
  NAND4BBX4 U280 ( .AN(n15), .BN(n184), .C(n186), .D(n185), .Y(n166) );
  NAND2X4 U281 ( .A(n31), .B(n57), .Y(n167) );
  NOR2BX4 U282 ( .AN(n186), .B(n189), .Y(n188) );
  XOR2X4 U283 ( .A(n192), .B(n8), .Y(SUM[23]) );
  OR2X4 U284 ( .A(B[23]), .B(A[23]), .Y(n186) );
  OAI2BB1X4 U285 ( .A0N(n185), .A1N(n193), .B0(n194), .Y(n192) );
  OAI21X4 U286 ( .A0(n195), .A1(n196), .B0(n197), .Y(n193) );
  XOR2X4 U287 ( .A(n205), .B(n206), .Y(SUM[22]) );
  CLKINVX3 U288 ( .A(n185), .Y(n189) );
  OR2X4 U289 ( .A(A[22]), .B(B[22]), .Y(n185) );
  XOR2X4 U290 ( .A(n209), .B(n210), .Y(SUM[21]) );
  OR2X4 U291 ( .A(A[20]), .B(B[20]), .Y(n208) );
  OAI2BB1X4 U292 ( .A0N(n211), .A1N(n75), .B0(n212), .Y(n145) );
  OAI21X4 U293 ( .A0(n214), .A1(n213), .B0(n215), .Y(n202) );
  NOR2X4 U294 ( .A(n204), .B(n220), .Y(n211) );
  CLKINVX3 U295 ( .A(n199), .Y(n220) );
  NAND3X4 U296 ( .A(n221), .B(n222), .C(n223), .Y(n204) );
  OR2X4 U297 ( .A(A[19]), .B(B[19]), .Y(n216) );
  OAI21X4 U298 ( .A0(n237), .A1(n229), .B0(n230), .Y(n227) );
  XOR2X4 U299 ( .A(n232), .B(n233), .Y(n300) );
  XOR2X4 U300 ( .A(n228), .B(n236), .Y(SUM[17]) );
  AOI21X4 U301 ( .A0(n75), .A1(n222), .B0(n238), .Y(n237) );
  OR2X4 U302 ( .A(B[17]), .B(A[17]), .Y(n221) );
  XOR2X4 U303 ( .A(n39), .B(n239), .Y(SUM[16]) );
  OR2X4 U304 ( .A(A[16]), .B(B[16]), .Y(n222) );
  OAI21X4 U305 ( .A0(n256), .A1(n35), .B0(n257), .Y(n240) );
  AOI21X4 U306 ( .A0(n258), .A1(n259), .B0(n27), .Y(n256) );
  XOR2X4 U307 ( .A(n263), .B(n262), .Y(SUM[15]) );
  OR2X4 U308 ( .A(B[15]), .B(A[15]), .Y(n253) );
  AOI21X4 U309 ( .A0(n36), .A1(n271), .B0(n272), .Y(n270) );
  OR2X4 U310 ( .A(A[14]), .B(B[14]), .Y(n254) );
  OR2X4 U311 ( .A(A[13]), .B(B[13]), .Y(n252) );
  XOR2X4 U312 ( .A(n275), .B(n276), .Y(SUM[12]) );
  OAI2BB1X4 U313 ( .A0N(n279), .A1N(n278), .B0(n280), .Y(n246) );
  NOR2X4 U314 ( .A(n83), .B(n34), .Y(n278) );
  NOR2X4 U315 ( .A(n282), .B(n283), .Y(n255) );
  NAND2X4 U316 ( .A(n284), .B(n87), .Y(n283) );
  OAI21X4 U317 ( .A0(B[11]), .A1(A[11]), .B0(n285), .Y(n282) );
  OR2X4 U318 ( .A(A[12]), .B(B[12]), .Y(n249) );
  OR2X4 U319 ( .A(B[10]), .B(A[10]), .Y(n285) );
  OR2X4 U320 ( .A(A[9]), .B(B[9]), .Y(n284) );
  NAND2X4 U321 ( .A(n291), .B(n86), .Y(n80) );
  OR2X4 U322 ( .A(B[8]), .B(A[8]), .Y(n87) );
  NAND4BBX4 U323 ( .AN(n102), .BN(n68), .C(n91), .D(n97), .Y(n250) );
  OR2X4 U324 ( .A(A[7]), .B(B[7]), .Y(n91) );
  OR2X4 U325 ( .A(A[6]), .B(B[6]), .Y(n97) );
  OR2X4 U326 ( .A(B[5]), .B(A[5]), .Y(n98) );
  OAI21X4 U327 ( .A0(n296), .A1(n297), .B0(n109), .Y(n105) );
  NAND2X4 U328 ( .A(n132), .B(n295), .Y(n297) );
  OR2X4 U329 ( .A(A[3]), .B(B[3]), .Y(n295) );
  OR2X4 U330 ( .A(A[2]), .B(B[2]), .Y(n132) );
  CLKINVX3 U331 ( .A(n133), .Y(n225) );
  OR2X4 U332 ( .A(A[1]), .B(B[1]), .Y(n133) );
endmodule


module hash_core_DW01_add_29 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203;

  NAND2X2 U2 ( .A(n114), .B(n115), .Y(n91) );
  OAI21X2 U3 ( .A0(n53), .A1(n54), .B0(n55), .Y(n51) );
  NAND2X2 U4 ( .A(n87), .B(n88), .Y(n66) );
  NAND2XL U5 ( .A(B[5]), .B(A[5]), .Y(n33) );
  OAI21X2 U6 ( .A0(n66), .A1(n67), .B0(n68), .Y(n62) );
  NOR2XL U7 ( .A(A[5]), .B(B[5]), .Y(n8) );
  INVX1 U8 ( .A(n193), .Y(n163) );
  OAI21X1 U9 ( .A0(n117), .A1(n118), .B0(n119), .Y(n114) );
  INVXL U10 ( .A(n161), .Y(n197) );
  INVXL U11 ( .A(n157), .Y(n192) );
  NOR2BX1 U12 ( .AN(n77), .B(n69), .Y(n68) );
  OAI21X1 U13 ( .A0(n91), .A1(n92), .B0(n93), .Y(n87) );
  NAND3BXL U14 ( .AN(n15), .B(n130), .C(n131), .Y(n118) );
  NOR2XL U15 ( .A(n5), .B(n7), .Y(n179) );
  AOI21XL U16 ( .A0(n20), .A1(n23), .B0(n6), .Y(n180) );
  AOI21XL U17 ( .A0(n151), .A1(n152), .B0(n153), .Y(n149) );
  NAND2XL U18 ( .A(n66), .B(n75), .Y(n84) );
  NAND2XL U19 ( .A(n91), .B(n101), .Y(n112) );
  XNOR2X1 U20 ( .A(n62), .B(n1), .Y(SUM[28]) );
  NAND2X1 U21 ( .A(n65), .B(n63), .Y(n1) );
  XNOR2X1 U22 ( .A(n51), .B(n2), .Y(SUM[30]) );
  NAND2X1 U23 ( .A(n49), .B(n52), .Y(n2) );
  NOR2BXL U24 ( .AN(n150), .B(n12), .Y(n169) );
  NAND2XL U25 ( .A(n117), .B(n127), .Y(n140) );
  NAND2XL U26 ( .A(n36), .B(n37), .Y(n34) );
  NAND2XL U27 ( .A(n38), .B(n39), .Y(n36) );
  INVXL U28 ( .A(n134), .Y(n59) );
  NOR2BXL U29 ( .AN(n182), .B(n6), .Y(n190) );
  NOR2BXL U30 ( .AN(n26), .B(n3), .Y(n25) );
  NOR2BXL U31 ( .AN(n33), .B(n8), .Y(n35) );
  NOR2BXL U32 ( .AN(n20), .B(n5), .Y(n19) );
  NOR2BXL U33 ( .AN(n183), .B(n7), .Y(n187) );
  NOR2BXL U34 ( .AN(n156), .B(n4), .Y(n174) );
  NOR2BXL U35 ( .AN(n23), .B(n11), .Y(n22) );
  NOR2BXL U36 ( .AN(n44), .B(n9), .Y(n43) );
  NOR2BXL U37 ( .AN(n29), .B(n31), .Y(n30) );
  NOR2BXL U38 ( .AN(n123), .B(n124), .Y(n139) );
  NOR2BXL U39 ( .AN(n154), .B(n167), .Y(n171) );
  NOR2BXL U40 ( .AN(n128), .B(n126), .Y(n141) );
  NOR2BXL U41 ( .AN(n37), .B(n41), .Y(n40) );
  NOR2BXL U42 ( .AN(n60), .B(n133), .Y(n132) );
  AND2X1 U43 ( .A(n127), .B(n143), .Y(n144) );
  XOR2XL U44 ( .A(n61), .B(n54), .Y(SUM[29]) );
  NOR2XL U45 ( .A(A[27]), .B(B[27]), .Y(n16) );
  NAND2XL U46 ( .A(B[26]), .B(A[26]), .Y(n71) );
  NAND2XL U47 ( .A(B[24]), .B(A[24]), .Y(n75) );
  NAND2XL U48 ( .A(B[25]), .B(A[25]), .Y(n76) );
  OR2XL U49 ( .A(A[25]), .B(B[25]), .Y(n79) );
  OR2XL U50 ( .A(A[26]), .B(B[26]), .Y(n78) );
  NAND2XL U51 ( .A(B[28]), .B(A[28]), .Y(n65) );
  NAND2XL U52 ( .A(B[27]), .B(A[27]), .Y(n77) );
  OR2XL U53 ( .A(A[28]), .B(B[28]), .Y(n63) );
  OR2XL U54 ( .A(A[24]), .B(B[24]), .Y(n88) );
  INVX1 U55 ( .A(n21), .Y(n178) );
  NAND3X1 U56 ( .A(n145), .B(n146), .C(n147), .Y(n142) );
  INVX1 U57 ( .A(n148), .Y(n147) );
  AOI2BB2X1 U58 ( .B0(n162), .B1(n163), .A0N(n164), .A1N(n158), .Y(n145) );
  NAND3BX1 U59 ( .AN(n157), .B(n160), .C(n161), .Y(n146) );
  NOR2X1 U60 ( .A(n159), .B(n158), .Y(n162) );
  NOR2X1 U61 ( .A(n158), .B(n159), .Y(n160) );
  OAI21XL U62 ( .A0(n178), .A1(n159), .B0(n164), .Y(n176) );
  INVX1 U63 ( .A(n197), .Y(n38) );
  OAI2BB1X1 U64 ( .A0N(n192), .A1N(n38), .B0(n193), .Y(n21) );
  AOI21X1 U65 ( .A0(n79), .A1(n84), .B0(n85), .Y(n82) );
  INVX1 U66 ( .A(n76), .Y(n85) );
  AOI21X1 U67 ( .A0(n62), .A1(n63), .B0(n64), .Y(n54) );
  INVX1 U68 ( .A(n65), .Y(n64) );
  INVX1 U69 ( .A(n27), .Y(n31) );
  INVX1 U70 ( .A(n151), .Y(n167) );
  NAND3BX1 U71 ( .AN(n14), .B(n104), .C(n105), .Y(n92) );
  NOR2X1 U72 ( .A(n94), .B(n95), .Y(n93) );
  INVX1 U73 ( .A(n103), .Y(n94) );
  NOR2X1 U74 ( .A(n120), .B(n121), .Y(n119) );
  INVX1 U75 ( .A(n129), .Y(n120) );
  NAND3BX1 U76 ( .AN(n16), .B(n78), .C(n79), .Y(n67) );
  INVX1 U77 ( .A(n39), .Y(n41) );
  INVX1 U78 ( .A(n56), .Y(n53) );
  NAND2X1 U79 ( .A(n184), .B(n185), .Y(n159) );
  NOR2X1 U80 ( .A(n11), .B(n5), .Y(n185) );
  NOR2X1 U81 ( .A(n6), .B(n7), .Y(n184) );
  AOI21X1 U82 ( .A0(n179), .A1(n180), .B0(n181), .Y(n164) );
  OAI21XL U83 ( .A0(n182), .A1(n7), .B0(n183), .Y(n181) );
  INVX1 U84 ( .A(n58), .Y(n133) );
  AOI21X1 U85 ( .A0(n60), .A1(n134), .B0(n133), .Y(n199) );
  NAND2X1 U86 ( .A(n165), .B(n166), .Y(n158) );
  NOR2X1 U87 ( .A(n4), .B(n13), .Y(n165) );
  NOR2X1 U88 ( .A(n12), .B(n167), .Y(n166) );
  XOR2X1 U89 ( .A(n106), .B(n107), .Y(SUM[23]) );
  NOR2BX1 U90 ( .AN(n103), .B(n14), .Y(n107) );
  OAI21XL U91 ( .A0(n108), .A1(n98), .B0(n97), .Y(n106) );
  INVX1 U92 ( .A(n109), .Y(n108) );
  NAND2X1 U93 ( .A(n142), .B(n143), .Y(n117) );
  NOR2X1 U94 ( .A(n3), .B(n31), .Y(n195) );
  OAI21XL U95 ( .A0(n149), .A1(n12), .B0(n150), .Y(n148) );
  INVX1 U96 ( .A(n154), .Y(n153) );
  OAI21XL U97 ( .A0(n4), .A1(n155), .B0(n156), .Y(n152) );
  NAND2X1 U98 ( .A(n111), .B(n102), .Y(n109) );
  NAND2X1 U99 ( .A(n105), .B(n112), .Y(n111) );
  AOI21X1 U100 ( .A0(n194), .A1(n195), .B0(n196), .Y(n193) );
  AOI21X1 U101 ( .A0(n33), .A1(n37), .B0(n8), .Y(n194) );
  OAI21XL U102 ( .A0(n3), .A1(n29), .B0(n26), .Y(n196) );
  INVX1 U103 ( .A(n198), .Y(n161) );
  AOI21X1 U104 ( .A0(n199), .A1(n200), .B0(n201), .Y(n198) );
  NOR2X1 U105 ( .A(n9), .B(n10), .Y(n200) );
  OAI21XL U106 ( .A0(n9), .A1(n46), .B0(n44), .Y(n201) );
  NAND2X1 U107 ( .A(n202), .B(n203), .Y(n157) );
  NOR2X1 U108 ( .A(n3), .B(n31), .Y(n203) );
  NOR2X1 U109 ( .A(n8), .B(n41), .Y(n202) );
  XOR2X1 U110 ( .A(n80), .B(n81), .Y(SUM[27]) );
  NOR2BX1 U111 ( .AN(n77), .B(n16), .Y(n81) );
  OAI21XL U112 ( .A0(n82), .A1(n72), .B0(n71), .Y(n80) );
  OAI21XL U113 ( .A0(n11), .A1(n178), .B0(n23), .Y(n18) );
  OAI21XL U114 ( .A0(n5), .A1(n191), .B0(n20), .Y(n189) );
  INVX1 U115 ( .A(n18), .Y(n191) );
  INVX1 U116 ( .A(n104), .Y(n98) );
  INVX1 U117 ( .A(n130), .Y(n124) );
  OAI21XL U118 ( .A0(n32), .A1(n8), .B0(n33), .Y(n28) );
  INVX1 U119 ( .A(n34), .Y(n32) );
  OAI21XL U120 ( .A0(n188), .A1(n6), .B0(n182), .Y(n186) );
  INVX1 U121 ( .A(n189), .Y(n188) );
  INVX1 U122 ( .A(n79), .Y(n74) );
  INVX1 U123 ( .A(n105), .Y(n100) );
  INVX1 U124 ( .A(n131), .Y(n126) );
  OAI2BB1X1 U125 ( .A0N(n27), .A1N(n28), .B0(n29), .Y(n24) );
  AOI21X1 U126 ( .A0(n70), .A1(n71), .B0(n16), .Y(n69) );
  NAND2BX1 U127 ( .AN(n72), .B(n73), .Y(n70) );
  OAI21XL U128 ( .A0(n74), .A1(n75), .B0(n76), .Y(n73) );
  AOI21X1 U129 ( .A0(n96), .A1(n97), .B0(n14), .Y(n95) );
  NAND2BX1 U130 ( .AN(n98), .B(n99), .Y(n96) );
  OAI21XL U131 ( .A0(n100), .A1(n101), .B0(n102), .Y(n99) );
  AOI21X1 U132 ( .A0(n122), .A1(n123), .B0(n15), .Y(n121) );
  NAND2BX1 U133 ( .AN(n124), .B(n125), .Y(n122) );
  OAI21XL U134 ( .A0(n126), .A1(n127), .B0(n128), .Y(n125) );
  INVX1 U135 ( .A(n78), .Y(n72) );
  OAI2BB1X1 U136 ( .A0N(n131), .A1N(n140), .B0(n128), .Y(n138) );
  OAI21XL U137 ( .A0(n172), .A1(n4), .B0(n156), .Y(n170) );
  INVX1 U138 ( .A(n173), .Y(n172) );
  OAI21XL U139 ( .A0(n13), .A1(n175), .B0(n155), .Y(n173) );
  INVX1 U140 ( .A(n176), .Y(n175) );
  OAI21XL U141 ( .A0(n137), .A1(n124), .B0(n123), .Y(n135) );
  INVX1 U142 ( .A(n138), .Y(n137) );
  XOR2X1 U143 ( .A(n87), .B(n89), .Y(SUM[24]) );
  NOR2BX1 U144 ( .AN(n75), .B(n90), .Y(n89) );
  INVX1 U145 ( .A(n88), .Y(n90) );
  XOR2X1 U146 ( .A(n168), .B(n169), .Y(SUM[15]) );
  OAI2BB1X1 U147 ( .A0N(n151), .A1N(n170), .B0(n154), .Y(n168) );
  XOR2X1 U148 ( .A(n84), .B(n86), .Y(SUM[25]) );
  NOR2BX1 U149 ( .AN(n76), .B(n74), .Y(n86) );
  XOR2X1 U150 ( .A(n109), .B(n110), .Y(SUM[22]) );
  NOR2BX1 U151 ( .AN(n97), .B(n98), .Y(n110) );
  XOR2X1 U152 ( .A(n112), .B(n113), .Y(SUM[21]) );
  NOR2BX1 U153 ( .AN(n102), .B(n100), .Y(n113) );
  OAI21XL U154 ( .A0(n45), .A1(n10), .B0(n46), .Y(n42) );
  INVX1 U155 ( .A(n47), .Y(n45) );
  OAI2BB1X1 U156 ( .A0N(n58), .A1N(n59), .B0(n60), .Y(n47) );
  NOR2BX1 U157 ( .AN(n46), .B(n10), .Y(n57) );
  NOR2BX1 U158 ( .AN(n155), .B(n13), .Y(n177) );
  NOR2BX1 U159 ( .AN(n129), .B(n15), .Y(n136) );
  AND2X2 U160 ( .A(n101), .B(n115), .Y(n116) );
  NAND2X1 U161 ( .A(n71), .B(n78), .Y(n83) );
  NAND2X1 U162 ( .A(n55), .B(n56), .Y(n61) );
  XOR2X1 U163 ( .A(n135), .B(n136), .Y(SUM[19]) );
  XOR2X1 U164 ( .A(n138), .B(n139), .Y(SUM[18]) );
  XOR2X1 U165 ( .A(n114), .B(n116), .Y(SUM[20]) );
  XOR2X1 U166 ( .A(n83), .B(n82), .Y(SUM[26]) );
  XOR2X1 U167 ( .A(n140), .B(n141), .Y(SUM[17]) );
  XOR2X1 U168 ( .A(n142), .B(n144), .Y(SUM[16]) );
  XOR2X1 U169 ( .A(n173), .B(n174), .Y(SUM[13]) );
  XOR2X1 U170 ( .A(n176), .B(n177), .Y(SUM[12]) );
  XOR2X1 U171 ( .A(n59), .B(n132), .Y(SUM[1]) );
  XOR2X1 U172 ( .A(n170), .B(n171), .Y(SUM[14]) );
  XOR2X1 U173 ( .A(n186), .B(n187), .Y(SUM[11]) );
  XOR2X1 U174 ( .A(n189), .B(n190), .Y(SUM[10]) );
  XOR2X1 U175 ( .A(n18), .B(n19), .Y(SUM[9]) );
  XOR2X1 U176 ( .A(n21), .B(n22), .Y(SUM[8]) );
  XOR2X1 U177 ( .A(n24), .B(n25), .Y(SUM[7]) );
  XOR2X1 U178 ( .A(n28), .B(n30), .Y(SUM[6]) );
  XOR2X1 U179 ( .A(n34), .B(n35), .Y(SUM[5]) );
  XOR2X1 U180 ( .A(n42), .B(n43), .Y(SUM[3]) );
  XOR2X1 U181 ( .A(n38), .B(n40), .Y(SUM[4]) );
  NOR2BX1 U182 ( .AN(n134), .B(n17), .Y(SUM[0]) );
  XOR2X1 U183 ( .A(n47), .B(n57), .Y(SUM[2]) );
  NOR2XL U184 ( .A(A[7]), .B(B[7]), .Y(n3) );
  NOR2XL U185 ( .A(A[13]), .B(B[13]), .Y(n4) );
  NOR2XL U186 ( .A(A[9]), .B(B[9]), .Y(n5) );
  NOR2XL U187 ( .A(A[10]), .B(B[10]), .Y(n6) );
  NOR2XL U188 ( .A(A[11]), .B(B[11]), .Y(n7) );
  NOR2XL U189 ( .A(A[3]), .B(B[3]), .Y(n9) );
  NOR2XL U190 ( .A(A[2]), .B(B[2]), .Y(n10) );
  NOR2XL U191 ( .A(A[8]), .B(B[8]), .Y(n11) );
  NOR2XL U192 ( .A(A[15]), .B(B[15]), .Y(n12) );
  NOR2XL U193 ( .A(A[12]), .B(B[12]), .Y(n13) );
  NAND2XL U194 ( .A(B[12]), .B(A[12]), .Y(n155) );
  XOR3X2 U195 ( .A(B[31]), .B(A[31]), .C(n48), .Y(SUM[31]) );
  NAND2X1 U196 ( .A(n49), .B(n50), .Y(n48) );
  NAND2X1 U197 ( .A(n51), .B(n52), .Y(n50) );
  NOR2XL U198 ( .A(A[23]), .B(B[23]), .Y(n14) );
  NOR2XL U199 ( .A(A[19]), .B(B[19]), .Y(n15) );
  NAND2XL U200 ( .A(B[22]), .B(A[22]), .Y(n97) );
  NAND2XL U201 ( .A(B[16]), .B(A[16]), .Y(n127) );
  NAND2XL U202 ( .A(B[20]), .B(A[20]), .Y(n101) );
  NAND2XL U203 ( .A(B[18]), .B(A[18]), .Y(n123) );
  NAND2XL U204 ( .A(B[21]), .B(A[21]), .Y(n102) );
  NAND2XL U205 ( .A(B[13]), .B(A[13]), .Y(n156) );
  NAND2XL U206 ( .A(B[17]), .B(A[17]), .Y(n128) );
  OR2XL U207 ( .A(A[21]), .B(B[21]), .Y(n105) );
  NAND2XL U208 ( .A(B[15]), .B(A[15]), .Y(n150) );
  OR2XL U209 ( .A(A[17]), .B(B[17]), .Y(n131) );
  NAND2XL U210 ( .A(B[19]), .B(A[19]), .Y(n129) );
  OR2XL U211 ( .A(A[16]), .B(B[16]), .Y(n143) );
  OR2XL U212 ( .A(A[22]), .B(B[22]), .Y(n104) );
  OR2XL U213 ( .A(A[18]), .B(B[18]), .Y(n130) );
  NAND2XL U214 ( .A(B[23]), .B(A[23]), .Y(n103) );
  OR2XL U215 ( .A(A[20]), .B(B[20]), .Y(n115) );
  OR2X2 U216 ( .A(A[29]), .B(B[29]), .Y(n56) );
  NOR2XL U217 ( .A(A[0]), .B(B[0]), .Y(n17) );
  NAND2X1 U218 ( .A(B[30]), .B(A[30]), .Y(n49) );
  NAND2X1 U219 ( .A(B[29]), .B(A[29]), .Y(n55) );
  OR2X2 U220 ( .A(A[30]), .B(B[30]), .Y(n52) );
  NAND2XL U221 ( .A(B[0]), .B(A[0]), .Y(n134) );
  NAND2XL U222 ( .A(B[14]), .B(A[14]), .Y(n154) );
  OR2XL U223 ( .A(A[14]), .B(B[14]), .Y(n151) );
  NAND2XL U224 ( .A(B[8]), .B(A[8]), .Y(n23) );
  NAND2XL U225 ( .A(B[7]), .B(A[7]), .Y(n26) );
  OR2XL U226 ( .A(A[4]), .B(B[4]), .Y(n39) );
  NAND2XL U227 ( .A(B[4]), .B(A[4]), .Y(n37) );
  NAND2XL U228 ( .A(B[10]), .B(A[10]), .Y(n182) );
  NAND2XL U229 ( .A(B[11]), .B(A[11]), .Y(n183) );
  NAND2XL U230 ( .A(B[9]), .B(A[9]), .Y(n20) );
  NAND2XL U231 ( .A(B[2]), .B(A[2]), .Y(n46) );
  NAND2XL U232 ( .A(B[6]), .B(A[6]), .Y(n29) );
  OR2XL U233 ( .A(A[6]), .B(B[6]), .Y(n27) );
  NAND2XL U234 ( .A(B[3]), .B(A[3]), .Y(n44) );
  NAND2XL U235 ( .A(B[1]), .B(A[1]), .Y(n60) );
  OR2XL U236 ( .A(A[1]), .B(B[1]), .Y(n58) );
endmodule


module hash_core_DW01_add_28 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205;

  OAI21X1 U2 ( .A0(n118), .A1(n119), .B0(n120), .Y(n115) );
  NAND2X2 U3 ( .A(n143), .B(n144), .Y(n118) );
  NAND2X1 U4 ( .A(B[4]), .B(A[4]), .Y(n35) );
  AOI21X1 U5 ( .A0(n61), .A1(n62), .B0(n63), .Y(n53) );
  OR2X1 U6 ( .A(A[14]), .B(B[14]), .Y(n152) );
  OAI21X1 U7 ( .A0(n52), .A1(n53), .B0(n54), .Y(n48) );
  OAI21X4 U8 ( .A0(n67), .A1(n68), .B0(n69), .Y(n61) );
  NAND2X2 U9 ( .A(n88), .B(n89), .Y(n67) );
  OR2X2 U10 ( .A(A[4]), .B(B[4]), .Y(n36) );
  NOR2X1 U11 ( .A(n4), .B(n11), .Y(n188) );
  NOR2XL U12 ( .A(n6), .B(n3), .Y(n189) );
  OAI21XL U13 ( .A0(n182), .A1(n11), .B0(n183), .Y(n164) );
  NOR2BX1 U14 ( .AN(n156), .B(n9), .Y(n179) );
  OAI2BB1XL U15 ( .A0N(n196), .A1N(n162), .B0(n166), .Y(n19) );
  INVXL U16 ( .A(n158), .Y(n196) );
  INVXL U17 ( .A(n48), .Y(n50) );
  INVXL U18 ( .A(n61), .Y(n65) );
  INVXL U19 ( .A(n159), .Y(n163) );
  OAI21X1 U20 ( .A0(n92), .A1(n93), .B0(n94), .Y(n88) );
  NOR2BX1 U21 ( .AN(n78), .B(n70), .Y(n69) );
  AOI21XL U22 ( .A0(n152), .A1(n153), .B0(n154), .Y(n150) );
  NAND2XL U23 ( .A(n67), .B(n76), .Y(n85) );
  NAND2XL U24 ( .A(n92), .B(n102), .Y(n113) );
  NOR2XL U25 ( .A(n5), .B(n38), .Y(n204) );
  NOR2XL U26 ( .A(n2), .B(n29), .Y(n205) );
  NOR2BXL U27 ( .AN(n183), .B(n11), .Y(n191) );
  NAND2XL U28 ( .A(n34), .B(n35), .Y(n32) );
  NAND2XL U29 ( .A(n162), .B(n36), .Y(n34) );
  NAND2XL U30 ( .A(n118), .B(n128), .Y(n141) );
  NOR2BXL U31 ( .AN(n187), .B(n4), .Y(n194) );
  NOR2BXL U32 ( .AN(n18), .B(n3), .Y(n17) );
  NOR2BXL U33 ( .AN(n24), .B(n2), .Y(n23) );
  INVXL U34 ( .A(n135), .Y(n58) );
  NOR2BXL U35 ( .AN(n31), .B(n5), .Y(n33) );
  NOR2BXL U36 ( .AN(n157), .B(n1), .Y(n176) );
  NOR2BXL U37 ( .AN(n41), .B(n7), .Y(n40) );
  NOR2BXL U38 ( .AN(n151), .B(n8), .Y(n171) );
  NOR2BXL U39 ( .AN(n27), .B(n29), .Y(n28) );
  NOR2BXL U40 ( .AN(n155), .B(n169), .Y(n173) );
  NOR2BXL U41 ( .AN(n59), .B(n134), .Y(n133) );
  XOR2XL U42 ( .A(n60), .B(n53), .Y(SUM[29]) );
  NOR2XL U43 ( .A(A[19]), .B(B[19]), .Y(n13) );
  NAND2XL U44 ( .A(B[16]), .B(A[16]), .Y(n128) );
  NAND2XL U45 ( .A(B[20]), .B(A[20]), .Y(n102) );
  NAND2XL U46 ( .A(B[18]), .B(A[18]), .Y(n124) );
  NAND2XL U47 ( .A(B[17]), .B(A[17]), .Y(n129) );
  NAND2XL U48 ( .A(B[19]), .B(A[19]), .Y(n130) );
  OR2XL U49 ( .A(A[21]), .B(B[21]), .Y(n106) );
  OR2XL U50 ( .A(A[17]), .B(B[17]), .Y(n132) );
  OR2XL U51 ( .A(A[18]), .B(B[18]), .Y(n131) );
  OR2XL U52 ( .A(A[22]), .B(B[22]), .Y(n105) );
  OR2XL U53 ( .A(A[16]), .B(B[16]), .Y(n144) );
  NOR2XL U54 ( .A(A[23]), .B(B[23]), .Y(n12) );
  NAND2XL U55 ( .A(B[22]), .B(A[22]), .Y(n98) );
  NAND2XL U56 ( .A(B[24]), .B(A[24]), .Y(n76) );
  NAND2XL U57 ( .A(B[21]), .B(A[21]), .Y(n103) );
  NAND2XL U58 ( .A(B[25]), .B(A[25]), .Y(n77) );
  NAND2XL U59 ( .A(B[23]), .B(A[23]), .Y(n104) );
  OR2XL U60 ( .A(A[25]), .B(B[25]), .Y(n80) );
  OR2XL U61 ( .A(A[26]), .B(B[26]), .Y(n79) );
  OR2XL U62 ( .A(A[20]), .B(B[20]), .Y(n116) );
  NOR2XL U63 ( .A(A[27]), .B(B[27]), .Y(n14) );
  NAND2XL U64 ( .A(B[26]), .B(A[26]), .Y(n72) );
  NAND2XL U65 ( .A(B[27]), .B(A[27]), .Y(n78) );
  OR2XL U66 ( .A(A[24]), .B(B[24]), .Y(n89) );
  NAND2XL U67 ( .A(B[28]), .B(A[28]), .Y(n64) );
  NAND2XL U68 ( .A(B[29]), .B(A[29]), .Y(n54) );
  OR2XL U69 ( .A(A[28]), .B(B[28]), .Y(n62) );
  OR2XL U70 ( .A(A[29]), .B(B[29]), .Y(n55) );
  NAND2XL U71 ( .A(B[30]), .B(A[30]), .Y(n46) );
  OR2XL U72 ( .A(A[30]), .B(B[30]), .Y(n49) );
  INVX1 U73 ( .A(n19), .Y(n180) );
  XOR2X1 U74 ( .A(n115), .B(n117), .Y(SUM[20]) );
  XOR2X1 U75 ( .A(n178), .B(n179), .Y(SUM[12]) );
  XOR2X1 U76 ( .A(n107), .B(n108), .Y(SUM[23]) );
  XOR2X1 U77 ( .A(n26), .B(n28), .Y(SUM[6]) );
  XOR2X1 U78 ( .A(n32), .B(n33), .Y(SUM[5]) );
  XOR2X1 U79 ( .A(n58), .B(n133), .Y(SUM[1]) );
  XOR2X1 U80 ( .A(n136), .B(n137), .Y(SUM[19]) );
  XOR2X1 U81 ( .A(n172), .B(n173), .Y(SUM[14]) );
  NOR3X1 U82 ( .A(n166), .B(n160), .C(n159), .Y(n165) );
  NAND3X1 U83 ( .A(n146), .B(n147), .C(n148), .Y(n143) );
  INVX1 U84 ( .A(n149), .Y(n148) );
  NAND3BX1 U85 ( .AN(n158), .B(n161), .C(n162), .Y(n147) );
  AOI21X1 U86 ( .A0(n163), .A1(n164), .B0(n165), .Y(n146) );
  NOR2X1 U87 ( .A(n159), .B(n160), .Y(n161) );
  OAI21XL U88 ( .A0(n180), .A1(n160), .B0(n181), .Y(n178) );
  INVX1 U89 ( .A(n164), .Y(n181) );
  XOR2X1 U90 ( .A(n39), .B(n40), .Y(SUM[3]) );
  XOR2X1 U91 ( .A(n19), .B(n20), .Y(SUM[8]) );
  XOR2X1 U92 ( .A(n162), .B(n37), .Y(SUM[4]) );
  INVX1 U93 ( .A(n64), .Y(n63) );
  INVX1 U94 ( .A(n25), .Y(n29) );
  NAND3BX1 U95 ( .AN(n12), .B(n105), .C(n106), .Y(n93) );
  NOR2X1 U96 ( .A(n95), .B(n96), .Y(n94) );
  INVX1 U97 ( .A(n104), .Y(n95) );
  NAND3BX1 U98 ( .AN(n13), .B(n131), .C(n132), .Y(n119) );
  NOR2X1 U99 ( .A(n121), .B(n122), .Y(n120) );
  INVX1 U100 ( .A(n130), .Y(n121) );
  NAND3BX1 U101 ( .AN(n14), .B(n79), .C(n80), .Y(n68) );
  AOI21X1 U102 ( .A0(n184), .A1(n185), .B0(n186), .Y(n182) );
  INVX1 U103 ( .A(n187), .Y(n186) );
  NAND2X1 U104 ( .A(n18), .B(n21), .Y(n185) );
  INVX1 U105 ( .A(n55), .Y(n52) );
  AOI21X1 U106 ( .A0(n197), .A1(n198), .B0(n199), .Y(n166) );
  AOI21X1 U107 ( .A0(n31), .A1(n35), .B0(n5), .Y(n197) );
  NOR2X1 U108 ( .A(n2), .B(n29), .Y(n198) );
  OAI21XL U109 ( .A0(n2), .A1(n27), .B0(n24), .Y(n199) );
  NAND2X1 U110 ( .A(n188), .B(n189), .Y(n160) );
  NAND2X1 U111 ( .A(n167), .B(n168), .Y(n159) );
  NOR2X1 U112 ( .A(n8), .B(n169), .Y(n168) );
  NOR2X1 U113 ( .A(n1), .B(n9), .Y(n167) );
  INVX1 U114 ( .A(n152), .Y(n169) );
  INVX1 U115 ( .A(n36), .Y(n38) );
  OAI21XL U116 ( .A0(n7), .A1(n43), .B0(n41), .Y(n203) );
  INVX1 U117 ( .A(n57), .Y(n134) );
  NAND2X1 U118 ( .A(n115), .B(n116), .Y(n92) );
  OAI21XL U119 ( .A0(n150), .A1(n8), .B0(n151), .Y(n149) );
  INVX1 U120 ( .A(n155), .Y(n154) );
  OAI21XL U121 ( .A0(n1), .A1(n156), .B0(n157), .Y(n153) );
  NOR2X1 U122 ( .A(n3), .B(n4), .Y(n184) );
  INVX1 U123 ( .A(n200), .Y(n162) );
  AOI21X1 U124 ( .A0(n201), .A1(n202), .B0(n203), .Y(n200) );
  AOI21X1 U125 ( .A0(n59), .A1(n135), .B0(n134), .Y(n201) );
  NOR2X1 U126 ( .A(n7), .B(n10), .Y(n202) );
  NAND2X1 U127 ( .A(n204), .B(n205), .Y(n158) );
  AOI21X1 U128 ( .A0(n80), .A1(n85), .B0(n86), .Y(n83) );
  INVX1 U129 ( .A(n77), .Y(n86) );
  OAI21XL U130 ( .A0(n6), .A1(n180), .B0(n21), .Y(n16) );
  OAI21XL U131 ( .A0(n9), .A1(n177), .B0(n156), .Y(n175) );
  INVX1 U132 ( .A(n178), .Y(n177) );
  INVX1 U133 ( .A(n105), .Y(n99) );
  INVX1 U134 ( .A(n131), .Y(n125) );
  OAI21XL U135 ( .A0(n30), .A1(n5), .B0(n31), .Y(n26) );
  INVX1 U136 ( .A(n32), .Y(n30) );
  INVX1 U137 ( .A(n80), .Y(n75) );
  INVX1 U138 ( .A(n106), .Y(n101) );
  INVX1 U139 ( .A(n132), .Y(n127) );
  OAI21XL U140 ( .A0(n138), .A1(n125), .B0(n124), .Y(n136) );
  INVX1 U141 ( .A(n139), .Y(n138) );
  OAI21XL U142 ( .A0(n83), .A1(n73), .B0(n72), .Y(n81) );
  AOI21X1 U143 ( .A0(n97), .A1(n98), .B0(n12), .Y(n96) );
  NAND2BX1 U144 ( .AN(n99), .B(n100), .Y(n97) );
  OAI21XL U145 ( .A0(n101), .A1(n102), .B0(n103), .Y(n100) );
  AOI21X1 U146 ( .A0(n71), .A1(n72), .B0(n14), .Y(n70) );
  NAND2BX1 U147 ( .AN(n73), .B(n74), .Y(n71) );
  OAI21XL U148 ( .A0(n75), .A1(n76), .B0(n77), .Y(n74) );
  AOI21X1 U149 ( .A0(n123), .A1(n124), .B0(n13), .Y(n122) );
  NAND2BX1 U150 ( .AN(n125), .B(n126), .Y(n123) );
  OAI21XL U151 ( .A0(n127), .A1(n128), .B0(n129), .Y(n126) );
  NAND2X1 U152 ( .A(n112), .B(n103), .Y(n110) );
  NAND2X1 U153 ( .A(n106), .B(n113), .Y(n112) );
  OAI2BB1X1 U154 ( .A0N(n132), .A1N(n141), .B0(n129), .Y(n139) );
  OAI21XL U155 ( .A0(n174), .A1(n1), .B0(n157), .Y(n172) );
  INVX1 U156 ( .A(n175), .Y(n174) );
  OAI21XL U157 ( .A0(n3), .A1(n195), .B0(n18), .Y(n193) );
  INVX1 U158 ( .A(n16), .Y(n195) );
  OAI21XL U159 ( .A0(n109), .A1(n99), .B0(n98), .Y(n107) );
  INVX1 U160 ( .A(n110), .Y(n109) );
  XOR2X1 U161 ( .A(n22), .B(n23), .Y(SUM[7]) );
  OAI2BB1X1 U162 ( .A0N(n25), .A1N(n26), .B0(n27), .Y(n22) );
  XOR2X1 U163 ( .A(n88), .B(n90), .Y(SUM[24]) );
  NOR2BX1 U164 ( .AN(n76), .B(n91), .Y(n90) );
  INVX1 U165 ( .A(n89), .Y(n91) );
  XOR2X1 U166 ( .A(n193), .B(n194), .Y(SUM[10]) );
  XOR2X1 U167 ( .A(n16), .B(n17), .Y(SUM[9]) );
  XOR2X1 U168 ( .A(n190), .B(n191), .Y(SUM[11]) );
  OAI21XL U169 ( .A0(n192), .A1(n4), .B0(n187), .Y(n190) );
  INVX1 U170 ( .A(n193), .Y(n192) );
  XOR2X1 U171 ( .A(n85), .B(n87), .Y(SUM[25]) );
  NOR2BX1 U172 ( .AN(n77), .B(n75), .Y(n87) );
  XOR2X1 U173 ( .A(n110), .B(n111), .Y(SUM[22]) );
  NOR2BX1 U174 ( .AN(n98), .B(n99), .Y(n111) );
  OAI2BB1X1 U175 ( .A0N(n152), .A1N(n172), .B0(n155), .Y(n170) );
  INVX1 U176 ( .A(n79), .Y(n73) );
  NOR2BX1 U177 ( .AN(n21), .B(n6), .Y(n20) );
  XOR2X1 U178 ( .A(n44), .B(n56), .Y(SUM[2]) );
  NOR2BX1 U179 ( .AN(n43), .B(n10), .Y(n56) );
  NOR2BX1 U180 ( .AN(n124), .B(n125), .Y(n140) );
  NOR2BX1 U181 ( .AN(n78), .B(n14), .Y(n82) );
  NOR2BX1 U182 ( .AN(n104), .B(n12), .Y(n108) );
  NOR2BX1 U183 ( .AN(n130), .B(n13), .Y(n137) );
  OAI21XL U184 ( .A0(n42), .A1(n10), .B0(n43), .Y(n39) );
  INVX1 U185 ( .A(n44), .Y(n42) );
  NOR2BX1 U186 ( .AN(n103), .B(n101), .Y(n114) );
  NOR2BX1 U187 ( .AN(n129), .B(n127), .Y(n142) );
  NOR2BX1 U188 ( .AN(n35), .B(n38), .Y(n37) );
  AND2X2 U189 ( .A(n102), .B(n116), .Y(n117) );
  AND2X2 U190 ( .A(n128), .B(n144), .Y(n145) );
  OAI2BB1X1 U191 ( .A0N(n57), .A1N(n58), .B0(n59), .Y(n44) );
  NAND2X1 U192 ( .A(n64), .B(n62), .Y(n66) );
  NAND2X1 U193 ( .A(n46), .B(n49), .Y(n51) );
  NAND2X1 U194 ( .A(n72), .B(n79), .Y(n84) );
  NAND2X1 U195 ( .A(n54), .B(n55), .Y(n60) );
  XOR2X1 U196 ( .A(n139), .B(n140), .Y(SUM[18]) );
  XOR2X1 U197 ( .A(n141), .B(n142), .Y(SUM[17]) );
  XOR2X1 U198 ( .A(n113), .B(n114), .Y(SUM[21]) );
  XOR2X1 U199 ( .A(n65), .B(n66), .Y(SUM[28]) );
  XOR2X1 U200 ( .A(n81), .B(n82), .Y(SUM[27]) );
  NOR2BX1 U201 ( .AN(n135), .B(n15), .Y(SUM[0]) );
  XOR2X1 U202 ( .A(n143), .B(n145), .Y(SUM[16]) );
  XOR2X1 U203 ( .A(n170), .B(n171), .Y(SUM[15]) );
  XOR2X1 U204 ( .A(n175), .B(n176), .Y(SUM[13]) );
  XOR2X1 U205 ( .A(n84), .B(n83), .Y(SUM[26]) );
  XOR2X1 U206 ( .A(n50), .B(n51), .Y(SUM[30]) );
  NOR2XL U207 ( .A(A[13]), .B(B[13]), .Y(n1) );
  NOR2XL U208 ( .A(A[7]), .B(B[7]), .Y(n2) );
  NOR2XL U209 ( .A(A[9]), .B(B[9]), .Y(n3) );
  NOR2XL U210 ( .A(A[10]), .B(B[10]), .Y(n4) );
  NOR2XL U211 ( .A(A[5]), .B(B[5]), .Y(n5) );
  NOR2XL U212 ( .A(A[8]), .B(B[8]), .Y(n6) );
  NOR2XL U213 ( .A(A[3]), .B(B[3]), .Y(n7) );
  NOR2XL U214 ( .A(A[15]), .B(B[15]), .Y(n8) );
  NOR2XL U215 ( .A(A[12]), .B(B[12]), .Y(n9) );
  NOR2XL U216 ( .A(A[2]), .B(B[2]), .Y(n10) );
  NOR2XL U217 ( .A(A[11]), .B(B[11]), .Y(n11) );
  NAND2XL U218 ( .A(B[8]), .B(A[8]), .Y(n21) );
  XOR3X2 U219 ( .A(B[31]), .B(A[31]), .C(n45), .Y(SUM[31]) );
  NAND2X1 U220 ( .A(n46), .B(n47), .Y(n45) );
  NAND2X1 U221 ( .A(n48), .B(n49), .Y(n47) );
  OR2XL U222 ( .A(A[6]), .B(B[6]), .Y(n25) );
  OR2XL U223 ( .A(A[1]), .B(B[1]), .Y(n57) );
  NAND2XL U224 ( .A(B[12]), .B(A[12]), .Y(n156) );
  NAND2XL U225 ( .A(B[2]), .B(A[2]), .Y(n43) );
  NAND2XL U226 ( .A(B[5]), .B(A[5]), .Y(n31) );
  NAND2XL U227 ( .A(B[9]), .B(A[9]), .Y(n18) );
  NAND2XL U228 ( .A(B[13]), .B(A[13]), .Y(n157) );
  NAND2XL U229 ( .A(B[6]), .B(A[6]), .Y(n27) );
  NAND2XL U230 ( .A(B[1]), .B(A[1]), .Y(n59) );
  NAND2XL U231 ( .A(B[0]), .B(A[0]), .Y(n135) );
  NAND2XL U232 ( .A(B[10]), .B(A[10]), .Y(n187) );
  NAND2XL U233 ( .A(B[14]), .B(A[14]), .Y(n155) );
  NAND2XL U234 ( .A(B[3]), .B(A[3]), .Y(n41) );
  NAND2XL U235 ( .A(B[7]), .B(A[7]), .Y(n24) );
  NAND2XL U236 ( .A(B[15]), .B(A[15]), .Y(n151) );
  NAND2XL U237 ( .A(B[11]), .B(A[11]), .Y(n183) );
  NOR2XL U238 ( .A(A[0]), .B(B[0]), .Y(n15) );
endmodule


module hash_core_DW01_add_33 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204;

  OAI21X1 U2 ( .A0(n68), .A1(n69), .B0(n70), .Y(n62) );
  NAND2X2 U3 ( .A(n89), .B(n90), .Y(n68) );
  OAI21X2 U4 ( .A0(n92), .A1(n93), .B0(n94), .Y(n89) );
  NOR2XL U5 ( .A(A[5]), .B(B[5]), .Y(n5) );
  NOR2XL U6 ( .A(A[7]), .B(B[7]), .Y(n2) );
  NOR2XL U7 ( .A(A[3]), .B(B[3]), .Y(n7) );
  NAND2XL U8 ( .A(B[3]), .B(A[3]), .Y(n42) );
  NOR2X1 U9 ( .A(n1), .B(n8), .Y(n187) );
  NOR2BX1 U10 ( .AN(n155), .B(n11), .Y(n178) );
  INVXL U11 ( .A(n163), .Y(n180) );
  OAI2BB1XL U12 ( .A0N(n195), .A1N(n36), .B0(n165), .Y(n19) );
  INVXL U13 ( .A(n157), .Y(n195) );
  INVXL U14 ( .A(n49), .Y(n51) );
  INVXL U15 ( .A(n62), .Y(n66) );
  INVXL U16 ( .A(n158), .Y(n162) );
  NOR2BX1 U17 ( .AN(n103), .B(n95), .Y(n94) );
  OAI21X1 U18 ( .A0(n117), .A1(n118), .B0(n119), .Y(n114) );
  NOR2BX1 U19 ( .AN(n79), .B(n71), .Y(n70) );
  NOR2XL U20 ( .A(n6), .B(n4), .Y(n188) );
  AOI21XL U21 ( .A0(n151), .A1(n152), .B0(n153), .Y(n149) );
  NAND2XL U22 ( .A(n68), .B(n77), .Y(n86) );
  NAND2XL U23 ( .A(n92), .B(n101), .Y(n112) );
  NOR2XL U24 ( .A(n5), .B(n39), .Y(n203) );
  NOR2XL U25 ( .A(n2), .B(n29), .Y(n204) );
  NAND2XL U26 ( .A(n117), .B(n127), .Y(n140) );
  NAND2XL U27 ( .A(n34), .B(n35), .Y(n32) );
  NAND2XL U28 ( .A(n36), .B(n37), .Y(n34) );
  INVXL U29 ( .A(n134), .Y(n59) );
  NOR2BXL U30 ( .AN(n24), .B(n2), .Y(n23) );
  NOR2BXL U31 ( .AN(n31), .B(n5), .Y(n33) );
  NOR2BXL U32 ( .AN(n18), .B(n4), .Y(n17) );
  NOR2BXL U33 ( .AN(n186), .B(n1), .Y(n193) );
  NOR2BXL U34 ( .AN(n156), .B(n3), .Y(n175) );
  NOR2BXL U35 ( .AN(n42), .B(n7), .Y(n41) );
  NOR2BXL U36 ( .AN(n150), .B(n10), .Y(n170) );
  NOR2BXL U37 ( .AN(n182), .B(n8), .Y(n190) );
  NOR2BXL U38 ( .AN(n27), .B(n29), .Y(n28) );
  NOR2BXL U39 ( .AN(n154), .B(n168), .Y(n172) );
  NOR2BXL U40 ( .AN(n60), .B(n133), .Y(n132) );
  XOR2XL U41 ( .A(n61), .B(n54), .Y(SUM[29]) );
  NAND2XL U42 ( .A(B[24]), .B(A[24]), .Y(n77) );
  OR2XL U43 ( .A(A[24]), .B(B[24]), .Y(n90) );
  INVX1 U44 ( .A(n19), .Y(n179) );
  NOR3X1 U45 ( .A(n165), .B(n159), .C(n158), .Y(n164) );
  NAND3X1 U46 ( .A(n145), .B(n146), .C(n147), .Y(n142) );
  INVX1 U47 ( .A(n148), .Y(n147) );
  NAND3BX1 U48 ( .AN(n157), .B(n160), .C(n161), .Y(n146) );
  AOI21X1 U49 ( .A0(n162), .A1(n163), .B0(n164), .Y(n145) );
  NOR2X1 U50 ( .A(n158), .B(n159), .Y(n160) );
  OAI21XL U51 ( .A0(n179), .A1(n159), .B0(n180), .Y(n177) );
  INVX1 U52 ( .A(n199), .Y(n36) );
  INVX1 U53 ( .A(n56), .Y(n53) );
  INVX1 U54 ( .A(n151), .Y(n168) );
  NAND3BX1 U55 ( .AN(n14), .B(n104), .C(n105), .Y(n93) );
  NAND3BX1 U56 ( .AN(n12), .B(n130), .C(n131), .Y(n118) );
  NOR2X1 U57 ( .A(n120), .B(n121), .Y(n119) );
  INVX1 U58 ( .A(n129), .Y(n120) );
  NAND3BX1 U59 ( .AN(n13), .B(n80), .C(n81), .Y(n69) );
  AOI21X1 U60 ( .A0(n62), .A1(n63), .B0(n64), .Y(n54) );
  INVX1 U61 ( .A(n65), .Y(n64) );
  NAND2X1 U62 ( .A(n187), .B(n188), .Y(n159) );
  NAND2X1 U63 ( .A(n166), .B(n167), .Y(n158) );
  NOR2X1 U64 ( .A(n3), .B(n11), .Y(n166) );
  NOR2X1 U65 ( .A(n10), .B(n168), .Y(n167) );
  NAND2X1 U66 ( .A(n142), .B(n143), .Y(n117) );
  NAND2X1 U67 ( .A(n114), .B(n115), .Y(n92) );
  AOI21X1 U68 ( .A0(n81), .A1(n86), .B0(n87), .Y(n84) );
  INVX1 U69 ( .A(n78), .Y(n87) );
  INVX1 U70 ( .A(n25), .Y(n29) );
  OAI21XL U71 ( .A0(n181), .A1(n8), .B0(n182), .Y(n163) );
  AOI21X1 U72 ( .A0(n183), .A1(n184), .B0(n185), .Y(n181) );
  INVX1 U73 ( .A(n186), .Y(n185) );
  NAND2X1 U74 ( .A(n18), .B(n21), .Y(n184) );
  AOI21X1 U75 ( .A0(n196), .A1(n197), .B0(n198), .Y(n165) );
  AOI21X1 U76 ( .A0(n31), .A1(n35), .B0(n5), .Y(n196) );
  NOR2X1 U77 ( .A(n2), .B(n29), .Y(n197) );
  OAI21XL U78 ( .A0(n2), .A1(n27), .B0(n24), .Y(n198) );
  OAI21XL U79 ( .A0(n11), .A1(n176), .B0(n155), .Y(n174) );
  INVX1 U80 ( .A(n177), .Y(n176) );
  INVX1 U81 ( .A(n130), .Y(n124) );
  INVX1 U82 ( .A(n58), .Y(n133) );
  AOI21X1 U83 ( .A0(n60), .A1(n134), .B0(n133), .Y(n200) );
  INVX1 U84 ( .A(n131), .Y(n126) );
  INVX1 U85 ( .A(n37), .Y(n39) );
  OAI21XL U86 ( .A0(n84), .A1(n74), .B0(n73), .Y(n82) );
  OAI2BB1X1 U87 ( .A0N(n151), .A1N(n171), .B0(n154), .Y(n169) );
  NOR2X1 U88 ( .A(n4), .B(n1), .Y(n183) );
  OAI21XL U89 ( .A0(n149), .A1(n10), .B0(n150), .Y(n148) );
  INVX1 U90 ( .A(n154), .Y(n153) );
  OAI21XL U91 ( .A0(n3), .A1(n155), .B0(n156), .Y(n152) );
  INVX1 U92 ( .A(n199), .Y(n161) );
  AOI21X1 U93 ( .A0(n200), .A1(n201), .B0(n202), .Y(n199) );
  NOR2X1 U94 ( .A(n7), .B(n9), .Y(n201) );
  OAI21XL U95 ( .A0(n7), .A1(n44), .B0(n42), .Y(n202) );
  OAI21XL U96 ( .A0(n173), .A1(n3), .B0(n156), .Y(n171) );
  INVX1 U97 ( .A(n174), .Y(n173) );
  NAND2X1 U98 ( .A(n203), .B(n204), .Y(n157) );
  OAI21XL U99 ( .A0(n108), .A1(n98), .B0(n97), .Y(n106) );
  INVX1 U100 ( .A(n109), .Y(n108) );
  AOI21X1 U101 ( .A0(n122), .A1(n123), .B0(n12), .Y(n121) );
  NAND2BX1 U102 ( .AN(n124), .B(n125), .Y(n122) );
  OAI21XL U103 ( .A0(n126), .A1(n127), .B0(n128), .Y(n125) );
  NAND2X1 U104 ( .A(n111), .B(n102), .Y(n109) );
  NAND2X1 U105 ( .A(n105), .B(n112), .Y(n111) );
  OAI21XL U106 ( .A0(n4), .A1(n194), .B0(n18), .Y(n192) );
  INVX1 U107 ( .A(n16), .Y(n194) );
  OAI21XL U108 ( .A0(n6), .A1(n179), .B0(n21), .Y(n16) );
  INVX1 U109 ( .A(n104), .Y(n98) );
  OAI21XL U110 ( .A0(n30), .A1(n5), .B0(n31), .Y(n26) );
  INVX1 U111 ( .A(n32), .Y(n30) );
  INVX1 U112 ( .A(n81), .Y(n76) );
  INVX1 U113 ( .A(n105), .Y(n100) );
  AOI21X1 U114 ( .A0(n96), .A1(n97), .B0(n14), .Y(n95) );
  NAND2BX1 U115 ( .AN(n98), .B(n99), .Y(n96) );
  OAI21XL U116 ( .A0(n100), .A1(n101), .B0(n102), .Y(n99) );
  INVX1 U117 ( .A(n80), .Y(n74) );
  OAI2BB1X1 U118 ( .A0N(n131), .A1N(n140), .B0(n128), .Y(n138) );
  OAI21XL U119 ( .A0(n191), .A1(n1), .B0(n186), .Y(n189) );
  INVX1 U120 ( .A(n192), .Y(n191) );
  OAI21XL U121 ( .A0(n137), .A1(n124), .B0(n123), .Y(n135) );
  INVX1 U122 ( .A(n138), .Y(n137) );
  OAI2BB1X1 U123 ( .A0N(n25), .A1N(n26), .B0(n27), .Y(n22) );
  AOI21X1 U124 ( .A0(n72), .A1(n73), .B0(n13), .Y(n71) );
  NAND2BX1 U125 ( .AN(n74), .B(n75), .Y(n72) );
  OAI21XL U126 ( .A0(n76), .A1(n77), .B0(n78), .Y(n75) );
  XOR2X1 U127 ( .A(n138), .B(n139), .Y(SUM[18]) );
  NOR2BX1 U128 ( .AN(n123), .B(n124), .Y(n139) );
  OAI21XL U129 ( .A0(n43), .A1(n9), .B0(n44), .Y(n40) );
  INVX1 U130 ( .A(n45), .Y(n43) );
  OAI2BB1X1 U131 ( .A0N(n58), .A1N(n59), .B0(n60), .Y(n45) );
  NOR2BX1 U132 ( .AN(n21), .B(n6), .Y(n20) );
  NOR2BX1 U133 ( .AN(n44), .B(n9), .Y(n57) );
  NOR2BX1 U134 ( .AN(n129), .B(n12), .Y(n136) );
  NOR2BX1 U135 ( .AN(n97), .B(n98), .Y(n110) );
  NOR2BX1 U136 ( .AN(n79), .B(n13), .Y(n83) );
  NOR2BX1 U137 ( .AN(n103), .B(n14), .Y(n107) );
  NOR2BX1 U138 ( .AN(n78), .B(n76), .Y(n88) );
  NOR2BX1 U139 ( .AN(n102), .B(n100), .Y(n113) );
  NOR2BX1 U140 ( .AN(n128), .B(n126), .Y(n141) );
  NOR2BX1 U141 ( .AN(n35), .B(n39), .Y(n38) );
  NAND2X1 U142 ( .A(n65), .B(n63), .Y(n67) );
  NAND2X1 U143 ( .A(n47), .B(n50), .Y(n52) );
  NAND2X1 U144 ( .A(n73), .B(n80), .Y(n85) );
  AND2X2 U145 ( .A(n127), .B(n143), .Y(n144) );
  AND2X2 U146 ( .A(n101), .B(n115), .Y(n116) );
  AND2X2 U147 ( .A(n77), .B(n90), .Y(n91) );
  XOR2X1 U148 ( .A(n135), .B(n136), .Y(SUM[19]) );
  XOR2X1 U149 ( .A(n112), .B(n113), .Y(SUM[21]) );
  XOR2X1 U150 ( .A(n114), .B(n116), .Y(SUM[20]) );
  XOR2X1 U151 ( .A(n140), .B(n141), .Y(SUM[17]) );
  XOR2X1 U152 ( .A(n189), .B(n190), .Y(SUM[11]) );
  XOR2X1 U153 ( .A(n192), .B(n193), .Y(SUM[10]) );
  XOR2X1 U154 ( .A(n19), .B(n20), .Y(SUM[8]) );
  XOR2X1 U155 ( .A(n171), .B(n172), .Y(SUM[14]) );
  XOR2X1 U156 ( .A(n40), .B(n41), .Y(SUM[3]) );
  XOR2X1 U157 ( .A(n16), .B(n17), .Y(SUM[9]) );
  XOR2X1 U158 ( .A(n174), .B(n175), .Y(SUM[13]) );
  XOR2X1 U159 ( .A(n142), .B(n144), .Y(SUM[16]) );
  XOR2X1 U160 ( .A(n109), .B(n110), .Y(SUM[22]) );
  XOR2X1 U161 ( .A(n85), .B(n84), .Y(SUM[26]) );
  XOR2X1 U162 ( .A(n86), .B(n88), .Y(SUM[25]) );
  XOR2X1 U163 ( .A(n82), .B(n83), .Y(SUM[27]) );
  XOR2X1 U164 ( .A(n106), .B(n107), .Y(SUM[23]) );
  XOR2X1 U165 ( .A(n177), .B(n178), .Y(SUM[12]) );
  XOR2X1 U166 ( .A(n89), .B(n91), .Y(SUM[24]) );
  XOR2X1 U167 ( .A(n66), .B(n67), .Y(SUM[28]) );
  XOR2X1 U168 ( .A(n51), .B(n52), .Y(SUM[30]) );
  XOR2X1 U169 ( .A(n22), .B(n23), .Y(SUM[7]) );
  XOR2X1 U170 ( .A(n169), .B(n170), .Y(SUM[15]) );
  XOR2X1 U171 ( .A(n45), .B(n57), .Y(SUM[2]) );
  XOR2X1 U172 ( .A(n26), .B(n28), .Y(SUM[6]) );
  XOR2X1 U173 ( .A(n32), .B(n33), .Y(SUM[5]) );
  XOR2X1 U174 ( .A(n36), .B(n38), .Y(SUM[4]) );
  XOR2X1 U175 ( .A(n59), .B(n132), .Y(SUM[1]) );
  NOR2BX1 U176 ( .AN(n134), .B(n15), .Y(SUM[0]) );
  NOR2XL U177 ( .A(A[10]), .B(B[10]), .Y(n1) );
  XOR3X2 U178 ( .A(B[31]), .B(A[31]), .C(n46), .Y(SUM[31]) );
  NAND2X1 U179 ( .A(n47), .B(n48), .Y(n46) );
  NAND2X1 U180 ( .A(n49), .B(n50), .Y(n48) );
  NOR2XL U181 ( .A(A[13]), .B(B[13]), .Y(n3) );
  NOR2XL U182 ( .A(A[9]), .B(B[9]), .Y(n4) );
  NOR2XL U183 ( .A(A[8]), .B(B[8]), .Y(n6) );
  NOR2XL U184 ( .A(A[11]), .B(B[11]), .Y(n8) );
  NOR2XL U185 ( .A(A[2]), .B(B[2]), .Y(n9) );
  NOR2XL U186 ( .A(A[15]), .B(B[15]), .Y(n10) );
  NOR2XL U187 ( .A(A[12]), .B(B[12]), .Y(n11) );
  NOR2XL U188 ( .A(A[19]), .B(B[19]), .Y(n12) );
  NAND2XL U189 ( .A(B[16]), .B(A[16]), .Y(n127) );
  NAND2XL U190 ( .A(B[12]), .B(A[12]), .Y(n155) );
  NAND2XL U191 ( .A(B[17]), .B(A[17]), .Y(n128) );
  NAND2XL U192 ( .A(B[13]), .B(A[13]), .Y(n156) );
  NAND2XL U193 ( .A(B[4]), .B(A[4]), .Y(n35) );
  NAND2XL U194 ( .A(B[5]), .B(A[5]), .Y(n31) );
  NAND2XL U195 ( .A(B[6]), .B(A[6]), .Y(n27) );
  OR2XL U196 ( .A(A[17]), .B(B[17]), .Y(n131) );
  OR2XL U197 ( .A(A[4]), .B(B[4]), .Y(n37) );
  OR2XL U198 ( .A(A[18]), .B(B[18]), .Y(n130) );
  OR2XL U199 ( .A(A[6]), .B(B[6]), .Y(n25) );
  NAND2XL U200 ( .A(B[26]), .B(A[26]), .Y(n73) );
  NOR2XL U201 ( .A(A[27]), .B(B[27]), .Y(n13) );
  NOR2XL U202 ( .A(A[23]), .B(B[23]), .Y(n14) );
  NAND2XL U203 ( .A(B[22]), .B(A[22]), .Y(n97) );
  NAND2XL U204 ( .A(B[20]), .B(A[20]), .Y(n101) );
  NAND2XL U205 ( .A(B[21]), .B(A[21]), .Y(n102) );
  NAND2XL U206 ( .A(B[25]), .B(A[25]), .Y(n78) );
  NAND2XL U207 ( .A(B[18]), .B(A[18]), .Y(n123) );
  OR2XL U208 ( .A(A[25]), .B(B[25]), .Y(n81) );
  OR2XL U209 ( .A(A[21]), .B(B[21]), .Y(n105) );
  OR2XL U210 ( .A(A[26]), .B(B[26]), .Y(n80) );
  NAND2XL U211 ( .A(B[23]), .B(A[23]), .Y(n103) );
  NAND2XL U212 ( .A(B[15]), .B(A[15]), .Y(n150) );
  OR2XL U213 ( .A(A[16]), .B(B[16]), .Y(n143) );
  OR2XL U214 ( .A(A[20]), .B(B[20]), .Y(n115) );
  OR2XL U215 ( .A(A[22]), .B(B[22]), .Y(n104) );
  NAND2XL U216 ( .A(B[28]), .B(A[28]), .Y(n65) );
  NAND2XL U217 ( .A(B[27]), .B(A[27]), .Y(n79) );
  OR2XL U218 ( .A(A[28]), .B(B[28]), .Y(n63) );
  NOR2XL U219 ( .A(A[0]), .B(B[0]), .Y(n15) );
  NAND2XL U220 ( .A(B[30]), .B(A[30]), .Y(n47) );
  OR2XL U221 ( .A(A[30]), .B(B[30]), .Y(n50) );
  NAND2XL U222 ( .A(B[19]), .B(A[19]), .Y(n129) );
  NAND2XL U223 ( .A(B[8]), .B(A[8]), .Y(n21) );
  NAND2XL U224 ( .A(B[10]), .B(A[10]), .Y(n186) );
  NAND2XL U225 ( .A(B[11]), .B(A[11]), .Y(n182) );
  NAND2XL U226 ( .A(B[14]), .B(A[14]), .Y(n154) );
  OR2XL U227 ( .A(A[14]), .B(B[14]), .Y(n151) );
  NAND2XL U228 ( .A(B[9]), .B(A[9]), .Y(n18) );
  NAND2X1 U229 ( .A(B[29]), .B(A[29]), .Y(n55) );
  OR2X2 U230 ( .A(A[29]), .B(B[29]), .Y(n56) );
  OAI21XL U231 ( .A0(n53), .A1(n54), .B0(n55), .Y(n49) );
  NAND2X1 U232 ( .A(n55), .B(n56), .Y(n61) );
  NAND2XL U233 ( .A(B[7]), .B(A[7]), .Y(n24) );
  NAND2XL U234 ( .A(B[2]), .B(A[2]), .Y(n44) );
  NAND2XL U235 ( .A(B[1]), .B(A[1]), .Y(n60) );
  OR2XL U236 ( .A(A[1]), .B(B[1]), .Y(n58) );
  NAND2XL U237 ( .A(B[0]), .B(A[0]), .Y(n134) );
endmodule


module hash_core_DW01_add_32 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203;

  NAND2X2 U2 ( .A(n112), .B(n113), .Y(n90) );
  OAI21X2 U3 ( .A0(n115), .A1(n116), .B0(n117), .Y(n112) );
  OAI21XL U4 ( .A0(n66), .A1(n67), .B0(n68), .Y(n60) );
  OAI21X1 U5 ( .A0(n90), .A1(n91), .B0(n92), .Y(n87) );
  CLKINVX3 U6 ( .A(n197), .Y(n159) );
  OAI2BB1X1 U7 ( .A0N(n193), .A1N(n159), .B0(n163), .Y(n18) );
  NOR2X1 U8 ( .A(n4), .B(n10), .Y(n185) );
  NOR2BX1 U9 ( .AN(n153), .B(n9), .Y(n176) );
  INVXL U10 ( .A(n161), .Y(n178) );
  INVXL U11 ( .A(n155), .Y(n193) );
  INVXL U12 ( .A(n47), .Y(n49) );
  INVXL U13 ( .A(n60), .Y(n64) );
  INVXL U14 ( .A(n156), .Y(n160) );
  NOR2BXL U15 ( .AN(n17), .B(n3), .Y(n16) );
  NOR2BXL U16 ( .AN(n23), .B(n2), .Y(n22) );
  NOR2BXL U17 ( .AN(n26), .B(n28), .Y(n27) );
  AND2X1 U18 ( .A(n132), .B(n203), .Y(SUM[0]) );
  NOR2BX1 U19 ( .AN(n101), .B(n93), .Y(n92) );
  NOR2BX1 U20 ( .AN(n77), .B(n69), .Y(n68) );
  NOR2XL U21 ( .A(n7), .B(n3), .Y(n186) );
  AOI21XL U22 ( .A0(n149), .A1(n150), .B0(n151), .Y(n147) );
  NAND2XL U23 ( .A(n66), .B(n75), .Y(n84) );
  NAND2XL U24 ( .A(n90), .B(n99), .Y(n110) );
  NOR2XL U25 ( .A(n2), .B(n28), .Y(n202) );
  NOR2XL U26 ( .A(n5), .B(n37), .Y(n201) );
  NAND2XL U27 ( .A(n115), .B(n125), .Y(n138) );
  NOR2BXL U28 ( .AN(n184), .B(n4), .Y(n191) );
  NAND2XL U29 ( .A(n33), .B(n34), .Y(n31) );
  NAND2XL U30 ( .A(n159), .B(n35), .Y(n33) );
  NOR2BXL U31 ( .AN(n30), .B(n5), .Y(n32) );
  INVXL U32 ( .A(n132), .Y(n57) );
  NOR2BXL U33 ( .AN(n40), .B(n6), .Y(n39) );
  NOR2BXL U34 ( .AN(n154), .B(n1), .Y(n173) );
  NOR2BXL U35 ( .AN(n148), .B(n8), .Y(n168) );
  NOR2BXL U36 ( .AN(n180), .B(n10), .Y(n188) );
  NOR2BXL U37 ( .AN(n152), .B(n166), .Y(n170) );
  NOR2BXL U38 ( .AN(n58), .B(n131), .Y(n130) );
  XOR2XL U39 ( .A(n59), .B(n52), .Y(SUM[29]) );
  NOR2XL U40 ( .A(A[19]), .B(B[19]), .Y(n13) );
  NAND2XL U41 ( .A(B[16]), .B(A[16]), .Y(n125) );
  NAND2XL U42 ( .A(B[18]), .B(A[18]), .Y(n121) );
  NAND2XL U43 ( .A(B[17]), .B(A[17]), .Y(n126) );
  NAND2XL U44 ( .A(B[19]), .B(A[19]), .Y(n127) );
  OR2XL U45 ( .A(A[17]), .B(B[17]), .Y(n129) );
  OR2XL U46 ( .A(A[18]), .B(B[18]), .Y(n128) );
  OR2XL U47 ( .A(A[16]), .B(B[16]), .Y(n141) );
  NOR2XL U48 ( .A(A[23]), .B(B[23]), .Y(n12) );
  NAND2XL U49 ( .A(B[20]), .B(A[20]), .Y(n99) );
  NAND2XL U50 ( .A(B[22]), .B(A[22]), .Y(n95) );
  NAND2XL U51 ( .A(B[21]), .B(A[21]), .Y(n100) );
  NAND2XL U52 ( .A(B[23]), .B(A[23]), .Y(n101) );
  OR2XL U53 ( .A(A[25]), .B(B[25]), .Y(n79) );
  OR2XL U54 ( .A(A[21]), .B(B[21]), .Y(n103) );
  OR2XL U55 ( .A(A[22]), .B(B[22]), .Y(n102) );
  OR2XL U56 ( .A(A[20]), .B(B[20]), .Y(n113) );
  NOR2XL U57 ( .A(A[27]), .B(B[27]), .Y(n14) );
  NAND2XL U58 ( .A(B[26]), .B(A[26]), .Y(n71) );
  NAND2XL U59 ( .A(B[24]), .B(A[24]), .Y(n75) );
  NAND2XL U60 ( .A(B[25]), .B(A[25]), .Y(n76) );
  NAND2XL U61 ( .A(B[27]), .B(A[27]), .Y(n77) );
  OR2XL U62 ( .A(A[26]), .B(B[26]), .Y(n78) );
  OR2XL U63 ( .A(A[24]), .B(B[24]), .Y(n88) );
  INVX1 U64 ( .A(n18), .Y(n177) );
  NOR3X1 U65 ( .A(n163), .B(n157), .C(n156), .Y(n162) );
  NAND3X1 U66 ( .A(n143), .B(n144), .C(n145), .Y(n140) );
  NAND3BX1 U67 ( .AN(n155), .B(n158), .C(n159), .Y(n144) );
  INVX1 U68 ( .A(n146), .Y(n145) );
  AOI21X1 U69 ( .A0(n160), .A1(n161), .B0(n162), .Y(n143) );
  NOR2X1 U70 ( .A(n156), .B(n157), .Y(n158) );
  OAI21XL U71 ( .A0(n177), .A1(n157), .B0(n178), .Y(n175) );
  XOR2X1 U72 ( .A(n15), .B(n16), .Y(SUM[9]) );
  XOR2X1 U73 ( .A(n21), .B(n22), .Y(SUM[7]) );
  XOR2X1 U74 ( .A(n25), .B(n27), .Y(SUM[6]) );
  XOR2X1 U75 ( .A(n43), .B(n55), .Y(SUM[2]) );
  NOR2BX1 U76 ( .AN(n42), .B(n11), .Y(n55) );
  AOI21X1 U77 ( .A0(n60), .A1(n61), .B0(n62), .Y(n52) );
  INVX1 U78 ( .A(n63), .Y(n62) );
  INVX1 U79 ( .A(n24), .Y(n28) );
  NAND3BX1 U80 ( .AN(n12), .B(n102), .C(n103), .Y(n91) );
  NAND3BX1 U81 ( .AN(n13), .B(n128), .C(n129), .Y(n116) );
  NOR2X1 U82 ( .A(n118), .B(n119), .Y(n117) );
  INVX1 U83 ( .A(n127), .Y(n118) );
  NAND3BX1 U84 ( .AN(n14), .B(n78), .C(n79), .Y(n67) );
  OAI21XL U85 ( .A0(n179), .A1(n10), .B0(n180), .Y(n161) );
  AOI21X1 U86 ( .A0(n181), .A1(n182), .B0(n183), .Y(n179) );
  INVX1 U87 ( .A(n184), .Y(n183) );
  NAND2X1 U88 ( .A(n17), .B(n20), .Y(n182) );
  OAI21XL U89 ( .A0(n51), .A1(n52), .B0(n53), .Y(n47) );
  INVX1 U90 ( .A(n54), .Y(n51) );
  AOI21X1 U91 ( .A0(n194), .A1(n195), .B0(n196), .Y(n163) );
  NOR2X1 U92 ( .A(n2), .B(n28), .Y(n195) );
  OAI21XL U93 ( .A0(n2), .A1(n26), .B0(n23), .Y(n196) );
  AOI21X1 U94 ( .A0(n30), .A1(n34), .B0(n5), .Y(n194) );
  NAND2X1 U95 ( .A(n185), .B(n186), .Y(n157) );
  NAND2X1 U96 ( .A(n164), .B(n165), .Y(n156) );
  NOR2X1 U97 ( .A(n8), .B(n166), .Y(n165) );
  NOR2X1 U98 ( .A(n1), .B(n9), .Y(n164) );
  INVX1 U99 ( .A(n149), .Y(n166) );
  INVX1 U100 ( .A(n56), .Y(n131) );
  AOI21X1 U101 ( .A0(n58), .A1(n132), .B0(n131), .Y(n198) );
  NAND2X1 U102 ( .A(n87), .B(n88), .Y(n66) );
  NAND2X1 U103 ( .A(n140), .B(n141), .Y(n115) );
  OAI21XL U104 ( .A0(n147), .A1(n8), .B0(n148), .Y(n146) );
  INVX1 U105 ( .A(n152), .Y(n151) );
  OAI21XL U106 ( .A0(n1), .A1(n153), .B0(n154), .Y(n150) );
  NOR2X1 U107 ( .A(n3), .B(n4), .Y(n181) );
  NAND2X1 U108 ( .A(n201), .B(n202), .Y(n155) );
  AOI21X1 U109 ( .A0(n198), .A1(n199), .B0(n200), .Y(n197) );
  NOR2X1 U110 ( .A(n6), .B(n11), .Y(n199) );
  OAI21XL U111 ( .A0(n6), .A1(n42), .B0(n40), .Y(n200) );
  NAND2X1 U112 ( .A(n45), .B(n46), .Y(n44) );
  NAND2X1 U113 ( .A(n47), .B(n48), .Y(n46) );
  AOI21X1 U114 ( .A0(n79), .A1(n84), .B0(n85), .Y(n82) );
  INVX1 U115 ( .A(n76), .Y(n85) );
  OAI21XL U116 ( .A0(n7), .A1(n177), .B0(n20), .Y(n15) );
  OAI21XL U117 ( .A0(n9), .A1(n174), .B0(n153), .Y(n172) );
  INVX1 U118 ( .A(n175), .Y(n174) );
  INVX1 U119 ( .A(n102), .Y(n96) );
  INVX1 U120 ( .A(n128), .Y(n122) );
  INVX1 U121 ( .A(n103), .Y(n98) );
  INVX1 U122 ( .A(n129), .Y(n124) );
  INVX1 U123 ( .A(n35), .Y(n37) );
  OAI21XL U124 ( .A0(n106), .A1(n96), .B0(n95), .Y(n104) );
  INVX1 U125 ( .A(n107), .Y(n106) );
  OAI21XL U126 ( .A0(n82), .A1(n72), .B0(n71), .Y(n80) );
  AOI21X1 U127 ( .A0(n120), .A1(n121), .B0(n13), .Y(n119) );
  NAND2BX1 U128 ( .AN(n122), .B(n123), .Y(n120) );
  OAI21XL U129 ( .A0(n124), .A1(n125), .B0(n126), .Y(n123) );
  AOI21X1 U130 ( .A0(n94), .A1(n95), .B0(n12), .Y(n93) );
  NAND2BX1 U131 ( .AN(n96), .B(n97), .Y(n94) );
  OAI21XL U132 ( .A0(n98), .A1(n99), .B0(n100), .Y(n97) );
  OAI2BB1X1 U133 ( .A0N(n129), .A1N(n138), .B0(n126), .Y(n136) );
  OAI21XL U134 ( .A0(n189), .A1(n4), .B0(n184), .Y(n187) );
  INVX1 U135 ( .A(n190), .Y(n189) );
  OAI21XL U136 ( .A0(n171), .A1(n1), .B0(n154), .Y(n169) );
  INVX1 U137 ( .A(n172), .Y(n171) );
  OAI21XL U138 ( .A0(n3), .A1(n192), .B0(n17), .Y(n190) );
  INVX1 U139 ( .A(n15), .Y(n192) );
  OAI21XL U140 ( .A0(n135), .A1(n122), .B0(n121), .Y(n133) );
  INVX1 U141 ( .A(n136), .Y(n135) );
  OAI2BB1X1 U142 ( .A0N(n149), .A1N(n169), .B0(n152), .Y(n167) );
  XOR2X1 U143 ( .A(n190), .B(n191), .Y(SUM[10]) );
  NAND2X1 U144 ( .A(n109), .B(n100), .Y(n107) );
  NAND2X1 U145 ( .A(n103), .B(n110), .Y(n109) );
  OAI21XL U146 ( .A0(n29), .A1(n5), .B0(n30), .Y(n25) );
  INVX1 U147 ( .A(n31), .Y(n29) );
  INVX1 U148 ( .A(n79), .Y(n74) );
  AOI21X1 U149 ( .A0(n70), .A1(n71), .B0(n14), .Y(n69) );
  NAND2BX1 U150 ( .AN(n72), .B(n73), .Y(n70) );
  OAI21XL U151 ( .A0(n74), .A1(n75), .B0(n76), .Y(n73) );
  INVX1 U152 ( .A(n78), .Y(n72) );
  OAI2BB1X1 U153 ( .A0N(n56), .A1N(n57), .B0(n58), .Y(n43) );
  XOR2X1 U154 ( .A(n38), .B(n39), .Y(SUM[3]) );
  OAI21XL U155 ( .A0(n41), .A1(n11), .B0(n42), .Y(n38) );
  INVX1 U156 ( .A(n43), .Y(n41) );
  OAI2BB1X1 U157 ( .A0N(n24), .A1N(n25), .B0(n26), .Y(n21) );
  XOR2X1 U158 ( .A(n31), .B(n32), .Y(SUM[5]) );
  XOR2X1 U159 ( .A(n18), .B(n19), .Y(SUM[8]) );
  NOR2BX1 U160 ( .AN(n20), .B(n7), .Y(n19) );
  XOR2X1 U161 ( .A(n159), .B(n36), .Y(SUM[4]) );
  NOR2BX1 U162 ( .AN(n34), .B(n37), .Y(n36) );
  NOR2BX1 U163 ( .AN(n95), .B(n96), .Y(n108) );
  NOR2BX1 U164 ( .AN(n121), .B(n122), .Y(n137) );
  NOR2BX1 U165 ( .AN(n77), .B(n14), .Y(n81) );
  NOR2BX1 U166 ( .AN(n101), .B(n12), .Y(n105) );
  NOR2BX1 U167 ( .AN(n127), .B(n13), .Y(n134) );
  NOR2BX1 U168 ( .AN(n76), .B(n74), .Y(n86) );
  NOR2BX1 U169 ( .AN(n100), .B(n98), .Y(n111) );
  NOR2BX1 U170 ( .AN(n126), .B(n124), .Y(n139) );
  AND2X2 U171 ( .A(n75), .B(n88), .Y(n89) );
  AND2X2 U172 ( .A(n99), .B(n113), .Y(n114) );
  AND2X2 U173 ( .A(n125), .B(n141), .Y(n142) );
  NAND2X1 U174 ( .A(n63), .B(n61), .Y(n65) );
  NAND2X1 U175 ( .A(n45), .B(n48), .Y(n50) );
  XOR2X1 U176 ( .A(n57), .B(n130), .Y(SUM[1]) );
  NAND2X1 U177 ( .A(n71), .B(n78), .Y(n83) );
  NAND2X1 U178 ( .A(n53), .B(n54), .Y(n59) );
  XOR2X1 U179 ( .A(n87), .B(n89), .Y(SUM[24]) );
  XOR2X1 U180 ( .A(n140), .B(n142), .Y(SUM[16]) );
  XOR3X2 U181 ( .A(B[31]), .B(A[31]), .C(n44), .Y(SUM[31]) );
  XOR2X1 U182 ( .A(n83), .B(n82), .Y(SUM[26]) );
  XOR2X1 U183 ( .A(n133), .B(n134), .Y(SUM[19]) );
  XOR2X1 U184 ( .A(n136), .B(n137), .Y(SUM[18]) );
  XOR2X1 U185 ( .A(n138), .B(n139), .Y(SUM[17]) );
  XOR2X1 U186 ( .A(n107), .B(n108), .Y(SUM[22]) );
  XOR2X1 U187 ( .A(n167), .B(n168), .Y(SUM[15]) );
  XOR2X1 U188 ( .A(n169), .B(n170), .Y(SUM[14]) );
  XOR2X1 U189 ( .A(n172), .B(n173), .Y(SUM[13]) );
  XOR2X1 U190 ( .A(n175), .B(n176), .Y(SUM[12]) );
  XOR2X1 U191 ( .A(n187), .B(n188), .Y(SUM[11]) );
  XOR2X1 U192 ( .A(n84), .B(n86), .Y(SUM[25]) );
  XOR2X1 U193 ( .A(n49), .B(n50), .Y(SUM[30]) );
  XOR2X1 U194 ( .A(n104), .B(n105), .Y(SUM[23]) );
  XOR2X1 U195 ( .A(n112), .B(n114), .Y(SUM[20]) );
  XOR2X1 U196 ( .A(n80), .B(n81), .Y(SUM[27]) );
  XOR2X1 U197 ( .A(n64), .B(n65), .Y(SUM[28]) );
  XOR2X1 U198 ( .A(n110), .B(n111), .Y(SUM[21]) );
  NOR2XL U199 ( .A(A[13]), .B(B[13]), .Y(n1) );
  NOR2XL U200 ( .A(A[7]), .B(B[7]), .Y(n2) );
  NOR2XL U201 ( .A(A[9]), .B(B[9]), .Y(n3) );
  NOR2XL U202 ( .A(A[10]), .B(B[10]), .Y(n4) );
  NOR2XL U203 ( .A(A[5]), .B(B[5]), .Y(n5) );
  NOR2XL U204 ( .A(A[3]), .B(B[3]), .Y(n6) );
  NOR2XL U205 ( .A(A[8]), .B(B[8]), .Y(n7) );
  NOR2XL U206 ( .A(A[15]), .B(B[15]), .Y(n8) );
  NOR2XL U207 ( .A(A[12]), .B(B[12]), .Y(n9) );
  NOR2XL U208 ( .A(A[11]), .B(B[11]), .Y(n10) );
  OR2XL U209 ( .A(A[14]), .B(B[14]), .Y(n149) );
  OR2XL U210 ( .A(A[1]), .B(B[1]), .Y(n56) );
  OR2XL U211 ( .A(A[6]), .B(B[6]), .Y(n24) );
  NOR2XL U212 ( .A(A[2]), .B(B[2]), .Y(n11) );
  NAND2XL U213 ( .A(B[12]), .B(A[12]), .Y(n153) );
  NAND2XL U214 ( .A(B[4]), .B(A[4]), .Y(n34) );
  NAND2XL U215 ( .A(B[5]), .B(A[5]), .Y(n30) );
  NAND2XL U216 ( .A(B[13]), .B(A[13]), .Y(n154) );
  NAND2XL U217 ( .A(B[2]), .B(A[2]), .Y(n42) );
  NAND2XL U218 ( .A(B[9]), .B(A[9]), .Y(n17) );
  NAND2XL U219 ( .A(B[8]), .B(A[8]), .Y(n20) );
  NAND2XL U220 ( .A(B[1]), .B(A[1]), .Y(n58) );
  NAND2XL U221 ( .A(B[6]), .B(A[6]), .Y(n26) );
  NAND2XL U222 ( .A(B[0]), .B(A[0]), .Y(n132) );
  NAND2XL U223 ( .A(B[14]), .B(A[14]), .Y(n152) );
  NAND2XL U224 ( .A(B[10]), .B(A[10]), .Y(n184) );
  NAND2XL U225 ( .A(B[15]), .B(A[15]), .Y(n148) );
  NAND2XL U226 ( .A(B[11]), .B(A[11]), .Y(n180) );
  NAND2XL U227 ( .A(B[3]), .B(A[3]), .Y(n40) );
  NAND2XL U228 ( .A(B[7]), .B(A[7]), .Y(n23) );
  OR2XL U229 ( .A(A[4]), .B(B[4]), .Y(n35) );
  OR2X2 U230 ( .A(A[28]), .B(B[28]), .Y(n61) );
  NAND2X1 U231 ( .A(B[30]), .B(A[30]), .Y(n45) );
  NAND2X1 U232 ( .A(B[29]), .B(A[29]), .Y(n53) );
  NAND2X1 U233 ( .A(B[28]), .B(A[28]), .Y(n63) );
  OR2X2 U234 ( .A(A[30]), .B(B[30]), .Y(n48) );
  OR2X2 U235 ( .A(A[29]), .B(B[29]), .Y(n54) );
  OR2XL U236 ( .A(A[0]), .B(B[0]), .Y(n203) );
endmodule


module hash_core_DW01_add_31 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206;

  OAI21X1 U2 ( .A0(n52), .A1(n53), .B0(n54), .Y(n48) );
  OAI21X2 U3 ( .A0(n92), .A1(n93), .B0(n94), .Y(n88) );
  NOR2X1 U4 ( .A(n4), .B(n11), .Y(n189) );
  NOR2BX1 U5 ( .AN(n157), .B(n9), .Y(n180) );
  INVXL U6 ( .A(n165), .Y(n182) );
  OAI2BB1XL U7 ( .A0N(n197), .A1N(n163), .B0(n167), .Y(n19) );
  INVXL U8 ( .A(n159), .Y(n197) );
  INVXL U9 ( .A(n48), .Y(n50) );
  INVXL U10 ( .A(n61), .Y(n65) );
  INVXL U11 ( .A(n160), .Y(n164) );
  OAI21X1 U12 ( .A0(n118), .A1(n119), .B0(n120), .Y(n114) );
  NOR2BX1 U13 ( .AN(n103), .B(n95), .Y(n94) );
  NOR2BX1 U14 ( .AN(n78), .B(n70), .Y(n69) );
  NOR2XL U15 ( .A(n7), .B(n3), .Y(n190) );
  AOI21XL U16 ( .A0(n153), .A1(n154), .B0(n155), .Y(n151) );
  NAND2XL U17 ( .A(n67), .B(n76), .Y(n85) );
  NAND2XL U18 ( .A(n92), .B(n101), .Y(n112) );
  NOR2XL U19 ( .A(n5), .B(n38), .Y(n205) );
  NOR2XL U20 ( .A(n2), .B(n29), .Y(n206) );
  NOR2XL U21 ( .A(n6), .B(n10), .Y(n203) );
  NAND2XL U22 ( .A(n118), .B(n128), .Y(n141) );
  NAND2XL U23 ( .A(n34), .B(n35), .Y(n32) );
  NAND2XL U24 ( .A(n163), .B(n36), .Y(n34) );
  INVXL U25 ( .A(n135), .Y(n58) );
  NOR2BXL U26 ( .AN(n24), .B(n2), .Y(n23) );
  NOR2BXL U27 ( .AN(n31), .B(n5), .Y(n33) );
  NOR2BXL U28 ( .AN(n18), .B(n3), .Y(n17) );
  NOR2BXL U29 ( .AN(n188), .B(n4), .Y(n195) );
  NOR2BXL U30 ( .AN(n158), .B(n1), .Y(n177) );
  NOR2BXL U31 ( .AN(n41), .B(n6), .Y(n40) );
  NOR2BXL U32 ( .AN(n152), .B(n8), .Y(n172) );
  NOR2BXL U33 ( .AN(n184), .B(n11), .Y(n192) );
  NOR2BXL U34 ( .AN(n27), .B(n29), .Y(n28) );
  NOR2BXL U35 ( .AN(n156), .B(n170), .Y(n174) );
  NOR2BXL U36 ( .AN(n59), .B(n134), .Y(n133) );
  XOR2XL U37 ( .A(n60), .B(n53), .Y(SUM[29]) );
  NOR2XL U38 ( .A(A[19]), .B(B[19]), .Y(n13) );
  NAND2XL U39 ( .A(B[16]), .B(A[16]), .Y(n128) );
  NAND2XL U40 ( .A(B[18]), .B(A[18]), .Y(n124) );
  NAND2XL U41 ( .A(B[17]), .B(A[17]), .Y(n129) );
  OR2XL U42 ( .A(A[21]), .B(B[21]), .Y(n105) );
  OR2XL U43 ( .A(A[17]), .B(B[17]), .Y(n132) );
  OR2XL U44 ( .A(A[18]), .B(B[18]), .Y(n131) );
  OR2XL U45 ( .A(A[16]), .B(B[16]), .Y(n144) );
  NOR2XL U46 ( .A(A[23]), .B(B[23]), .Y(n12) );
  NAND2XL U47 ( .A(B[24]), .B(A[24]), .Y(n76) );
  NAND2XL U48 ( .A(B[25]), .B(A[25]), .Y(n77) );
  NAND2XL U49 ( .A(B[22]), .B(A[22]), .Y(n97) );
  NAND2XL U50 ( .A(B[20]), .B(A[20]), .Y(n101) );
  NAND2XL U51 ( .A(B[21]), .B(A[21]), .Y(n102) );
  NAND2XL U52 ( .A(B[23]), .B(A[23]), .Y(n103) );
  NAND2XL U53 ( .A(B[19]), .B(A[19]), .Y(n130) );
  OR2XL U54 ( .A(A[25]), .B(B[25]), .Y(n80) );
  OR2XL U55 ( .A(A[22]), .B(B[22]), .Y(n104) );
  OR2XL U56 ( .A(A[20]), .B(B[20]), .Y(n115) );
  NOR2XL U57 ( .A(A[27]), .B(B[27]), .Y(n14) );
  NAND2XL U58 ( .A(B[26]), .B(A[26]), .Y(n72) );
  NAND2XL U59 ( .A(B[27]), .B(A[27]), .Y(n78) );
  OR2XL U60 ( .A(A[26]), .B(B[26]), .Y(n79) );
  OR2XL U61 ( .A(A[24]), .B(B[24]), .Y(n89) );
  INVX1 U62 ( .A(n19), .Y(n181) );
  NOR3X1 U63 ( .A(n167), .B(n161), .C(n160), .Y(n166) );
  NAND3X1 U64 ( .A(n147), .B(n148), .C(n149), .Y(n143) );
  INVX1 U65 ( .A(n150), .Y(n149) );
  NAND3BX1 U66 ( .AN(n159), .B(n162), .C(n163), .Y(n148) );
  AOI21X1 U67 ( .A0(n164), .A1(n165), .B0(n166), .Y(n147) );
  NOR2X1 U68 ( .A(n160), .B(n161), .Y(n162) );
  OAI21XL U69 ( .A0(n181), .A1(n161), .B0(n182), .Y(n179) );
  AOI21X1 U70 ( .A0(n61), .A1(n62), .B0(n63), .Y(n53) );
  INVX1 U71 ( .A(n64), .Y(n63) );
  INVX1 U72 ( .A(n25), .Y(n29) );
  NAND3BX1 U73 ( .AN(n12), .B(n104), .C(n105), .Y(n93) );
  NAND3BX1 U74 ( .AN(n13), .B(n131), .C(n132), .Y(n119) );
  NOR2X1 U75 ( .A(n121), .B(n122), .Y(n120) );
  INVX1 U76 ( .A(n130), .Y(n121) );
  OAI21XL U77 ( .A0(n67), .A1(n68), .B0(n69), .Y(n61) );
  NAND3BX1 U78 ( .AN(n14), .B(n79), .C(n80), .Y(n68) );
  OAI21XL U79 ( .A0(n183), .A1(n11), .B0(n184), .Y(n165) );
  AOI21X1 U80 ( .A0(n185), .A1(n186), .B0(n187), .Y(n183) );
  INVX1 U81 ( .A(n188), .Y(n187) );
  NAND2X1 U82 ( .A(n18), .B(n21), .Y(n186) );
  INVX1 U83 ( .A(n55), .Y(n52) );
  AOI21X1 U84 ( .A0(n198), .A1(n199), .B0(n200), .Y(n167) );
  AOI21X1 U85 ( .A0(n31), .A1(n35), .B0(n5), .Y(n198) );
  NOR2X1 U86 ( .A(n2), .B(n29), .Y(n199) );
  OAI21XL U87 ( .A0(n2), .A1(n27), .B0(n24), .Y(n200) );
  NAND2X1 U88 ( .A(n189), .B(n190), .Y(n161) );
  NAND2X1 U89 ( .A(n168), .B(n169), .Y(n160) );
  NOR2X1 U90 ( .A(n8), .B(n170), .Y(n169) );
  NOR2X1 U91 ( .A(n1), .B(n9), .Y(n168) );
  INVX1 U92 ( .A(n153), .Y(n170) );
  INVX1 U93 ( .A(n57), .Y(n134) );
  NAND2X1 U94 ( .A(n143), .B(n144), .Y(n118) );
  NAND2X1 U95 ( .A(n88), .B(n89), .Y(n67) );
  NAND2X1 U96 ( .A(n114), .B(n115), .Y(n92) );
  OAI21XL U97 ( .A0(n151), .A1(n8), .B0(n152), .Y(n150) );
  INVX1 U98 ( .A(n156), .Y(n155) );
  OAI21XL U99 ( .A0(n1), .A1(n157), .B0(n158), .Y(n154) );
  NOR2X1 U100 ( .A(n3), .B(n4), .Y(n185) );
  INVX1 U101 ( .A(n201), .Y(n163) );
  AOI21X1 U102 ( .A0(n202), .A1(n203), .B0(n204), .Y(n201) );
  AOI21X1 U103 ( .A0(n59), .A1(n135), .B0(n134), .Y(n202) );
  OAI21XL U104 ( .A0(n6), .A1(n43), .B0(n41), .Y(n204) );
  NAND2X1 U105 ( .A(n205), .B(n206), .Y(n159) );
  AOI21X1 U106 ( .A0(n80), .A1(n85), .B0(n86), .Y(n83) );
  INVX1 U107 ( .A(n77), .Y(n86) );
  OAI21XL U108 ( .A0(n7), .A1(n181), .B0(n21), .Y(n16) );
  OAI21XL U109 ( .A0(n9), .A1(n178), .B0(n157), .Y(n176) );
  INVX1 U110 ( .A(n179), .Y(n178) );
  INVX1 U111 ( .A(n131), .Y(n125) );
  INVX1 U112 ( .A(n104), .Y(n98) );
  OAI21XL U113 ( .A0(n30), .A1(n5), .B0(n31), .Y(n26) );
  INVX1 U114 ( .A(n32), .Y(n30) );
  INVX1 U115 ( .A(n80), .Y(n75) );
  INVX1 U116 ( .A(n105), .Y(n100) );
  INVX1 U117 ( .A(n132), .Y(n127) );
  INVX1 U118 ( .A(n36), .Y(n38) );
  OAI21XL U119 ( .A0(n138), .A1(n125), .B0(n124), .Y(n136) );
  INVX1 U120 ( .A(n139), .Y(n138) );
  OAI21XL U121 ( .A0(n83), .A1(n73), .B0(n72), .Y(n81) );
  AOI21X1 U122 ( .A0(n71), .A1(n72), .B0(n14), .Y(n70) );
  NAND2BX1 U123 ( .AN(n73), .B(n74), .Y(n71) );
  OAI21XL U124 ( .A0(n75), .A1(n76), .B0(n77), .Y(n74) );
  AOI21X1 U125 ( .A0(n123), .A1(n124), .B0(n13), .Y(n122) );
  NAND2BX1 U126 ( .AN(n125), .B(n126), .Y(n123) );
  OAI21XL U127 ( .A0(n127), .A1(n128), .B0(n129), .Y(n126) );
  AOI21X1 U128 ( .A0(n96), .A1(n97), .B0(n12), .Y(n95) );
  NAND2BX1 U129 ( .AN(n98), .B(n99), .Y(n96) );
  OAI21XL U130 ( .A0(n100), .A1(n101), .B0(n102), .Y(n99) );
  NAND2X1 U131 ( .A(n111), .B(n102), .Y(n109) );
  NAND2X1 U132 ( .A(n105), .B(n112), .Y(n111) );
  OAI2BB1X1 U133 ( .A0N(n132), .A1N(n141), .B0(n129), .Y(n139) );
  OAI21XL U134 ( .A0(n193), .A1(n4), .B0(n188), .Y(n191) );
  INVX1 U135 ( .A(n194), .Y(n193) );
  OAI21XL U136 ( .A0(n175), .A1(n1), .B0(n158), .Y(n173) );
  INVX1 U137 ( .A(n176), .Y(n175) );
  OAI21XL U138 ( .A0(n3), .A1(n196), .B0(n18), .Y(n194) );
  INVX1 U139 ( .A(n16), .Y(n196) );
  OAI2BB1X1 U140 ( .A0N(n25), .A1N(n26), .B0(n27), .Y(n22) );
  OAI2BB1X1 U141 ( .A0N(n153), .A1N(n173), .B0(n156), .Y(n171) );
  XOR2X1 U142 ( .A(n88), .B(n90), .Y(SUM[24]) );
  NOR2BX1 U143 ( .AN(n76), .B(n91), .Y(n90) );
  INVX1 U144 ( .A(n89), .Y(n91) );
  XOR2X1 U145 ( .A(n85), .B(n87), .Y(SUM[25]) );
  NOR2BX1 U146 ( .AN(n77), .B(n75), .Y(n87) );
  XOR2X1 U147 ( .A(n106), .B(n107), .Y(SUM[23]) );
  NOR2BX1 U148 ( .AN(n103), .B(n12), .Y(n107) );
  OAI21XL U149 ( .A0(n108), .A1(n98), .B0(n97), .Y(n106) );
  INVX1 U150 ( .A(n109), .Y(n108) );
  OAI21XL U151 ( .A0(n42), .A1(n10), .B0(n43), .Y(n39) );
  INVX1 U152 ( .A(n44), .Y(n42) );
  INVX1 U153 ( .A(n79), .Y(n73) );
  OAI2BB1X1 U154 ( .A0N(n57), .A1N(n58), .B0(n59), .Y(n44) );
  XOR2X1 U155 ( .A(n114), .B(n116), .Y(SUM[20]) );
  NOR2BX1 U156 ( .AN(n101), .B(n117), .Y(n116) );
  INVX1 U157 ( .A(n115), .Y(n117) );
  XOR2X1 U158 ( .A(n143), .B(n145), .Y(SUM[16]) );
  NOR2BX1 U159 ( .AN(n128), .B(n146), .Y(n145) );
  INVX1 U160 ( .A(n144), .Y(n146) );
  NOR2BX1 U161 ( .AN(n21), .B(n7), .Y(n20) );
  NOR2BX1 U162 ( .AN(n43), .B(n10), .Y(n56) );
  NOR2BX1 U163 ( .AN(n97), .B(n98), .Y(n110) );
  NOR2BX1 U164 ( .AN(n124), .B(n125), .Y(n140) );
  NOR2BX1 U165 ( .AN(n78), .B(n14), .Y(n82) );
  NOR2BX1 U166 ( .AN(n130), .B(n13), .Y(n137) );
  NOR2BX1 U167 ( .AN(n102), .B(n100), .Y(n113) );
  NOR2BX1 U168 ( .AN(n129), .B(n127), .Y(n142) );
  NOR2BX1 U169 ( .AN(n35), .B(n38), .Y(n37) );
  NAND2X1 U170 ( .A(n64), .B(n62), .Y(n66) );
  NAND2X1 U171 ( .A(n46), .B(n49), .Y(n51) );
  NAND2X1 U172 ( .A(n72), .B(n79), .Y(n84) );
  NAND2X1 U173 ( .A(n54), .B(n55), .Y(n60) );
  XOR2X1 U174 ( .A(n136), .B(n137), .Y(SUM[19]) );
  XOR2X1 U175 ( .A(n19), .B(n20), .Y(SUM[8]) );
  XOR2X1 U176 ( .A(n58), .B(n133), .Y(SUM[1]) );
  XOR2X1 U177 ( .A(n173), .B(n174), .Y(SUM[14]) );
  XOR2X1 U178 ( .A(n179), .B(n180), .Y(SUM[12]) );
  XOR2X1 U179 ( .A(n26), .B(n28), .Y(SUM[6]) );
  XOR2X1 U180 ( .A(n32), .B(n33), .Y(SUM[5]) );
  XOR2X1 U181 ( .A(n163), .B(n37), .Y(SUM[4]) );
  XOR2X1 U182 ( .A(n84), .B(n83), .Y(SUM[26]) );
  XOR2X1 U183 ( .A(n139), .B(n140), .Y(SUM[18]) );
  XOR2X1 U184 ( .A(n141), .B(n142), .Y(SUM[17]) );
  XOR2X1 U185 ( .A(n112), .B(n113), .Y(SUM[21]) );
  XOR2X1 U186 ( .A(n171), .B(n172), .Y(SUM[15]) );
  XOR2X1 U187 ( .A(n176), .B(n177), .Y(SUM[13]) );
  XOR2X1 U188 ( .A(n81), .B(n82), .Y(SUM[27]) );
  XOR2X1 U189 ( .A(n65), .B(n66), .Y(SUM[28]) );
  XOR2X1 U190 ( .A(n16), .B(n17), .Y(SUM[9]) );
  XOR2X1 U191 ( .A(n109), .B(n110), .Y(SUM[22]) );
  XOR2X1 U192 ( .A(n191), .B(n192), .Y(SUM[11]) );
  XOR2X1 U193 ( .A(n194), .B(n195), .Y(SUM[10]) );
  XOR2X1 U194 ( .A(n22), .B(n23), .Y(SUM[7]) );
  XOR2X1 U195 ( .A(n39), .B(n40), .Y(SUM[3]) );
  XOR2X1 U196 ( .A(n44), .B(n56), .Y(SUM[2]) );
  NOR2BX1 U197 ( .AN(n135), .B(n15), .Y(SUM[0]) );
  XOR2X1 U198 ( .A(n50), .B(n51), .Y(SUM[30]) );
  NOR2XL U199 ( .A(A[13]), .B(B[13]), .Y(n1) );
  NOR2XL U200 ( .A(A[7]), .B(B[7]), .Y(n2) );
  NOR2XL U201 ( .A(A[9]), .B(B[9]), .Y(n3) );
  NOR2XL U202 ( .A(A[10]), .B(B[10]), .Y(n4) );
  NOR2XL U203 ( .A(A[5]), .B(B[5]), .Y(n5) );
  NOR2XL U204 ( .A(A[3]), .B(B[3]), .Y(n6) );
  NOR2XL U205 ( .A(A[8]), .B(B[8]), .Y(n7) );
  NOR2XL U206 ( .A(A[15]), .B(B[15]), .Y(n8) );
  NOR2XL U207 ( .A(A[12]), .B(B[12]), .Y(n9) );
  NOR2XL U208 ( .A(A[2]), .B(B[2]), .Y(n10) );
  NOR2XL U209 ( .A(A[11]), .B(B[11]), .Y(n11) );
  OR2XL U210 ( .A(A[14]), .B(B[14]), .Y(n153) );
  XOR3X2 U211 ( .A(B[31]), .B(A[31]), .C(n45), .Y(SUM[31]) );
  NAND2X1 U212 ( .A(n46), .B(n47), .Y(n45) );
  NAND2X1 U213 ( .A(n48), .B(n49), .Y(n47) );
  OR2XL U214 ( .A(A[1]), .B(B[1]), .Y(n57) );
  OR2XL U215 ( .A(A[6]), .B(B[6]), .Y(n25) );
  NAND2XL U216 ( .A(B[2]), .B(A[2]), .Y(n43) );
  NAND2XL U217 ( .A(B[4]), .B(A[4]), .Y(n35) );
  NAND2XL U218 ( .A(B[5]), .B(A[5]), .Y(n31) );
  NAND2XL U219 ( .A(B[12]), .B(A[12]), .Y(n157) );
  NAND2XL U220 ( .A(B[9]), .B(A[9]), .Y(n18) );
  NAND2XL U221 ( .A(B[13]), .B(A[13]), .Y(n158) );
  NAND2XL U222 ( .A(B[0]), .B(A[0]), .Y(n135) );
  NAND2XL U223 ( .A(B[8]), .B(A[8]), .Y(n21) );
  NAND2XL U224 ( .A(B[1]), .B(A[1]), .Y(n59) );
  NAND2XL U225 ( .A(B[6]), .B(A[6]), .Y(n27) );
  NAND2XL U226 ( .A(B[10]), .B(A[10]), .Y(n188) );
  NAND2XL U227 ( .A(B[14]), .B(A[14]), .Y(n156) );
  NAND2XL U228 ( .A(B[11]), .B(A[11]), .Y(n184) );
  NAND2XL U229 ( .A(B[7]), .B(A[7]), .Y(n24) );
  NAND2XL U230 ( .A(B[15]), .B(A[15]), .Y(n152) );
  NAND2XL U231 ( .A(B[3]), .B(A[3]), .Y(n41) );
  OR2XL U232 ( .A(A[4]), .B(B[4]), .Y(n36) );
  OR2X2 U233 ( .A(A[28]), .B(B[28]), .Y(n62) );
  NAND2X1 U234 ( .A(B[30]), .B(A[30]), .Y(n46) );
  NAND2X1 U235 ( .A(B[29]), .B(A[29]), .Y(n54) );
  NAND2X1 U236 ( .A(B[28]), .B(A[28]), .Y(n64) );
  OR2X2 U237 ( .A(A[30]), .B(B[30]), .Y(n49) );
  OR2X2 U238 ( .A(A[29]), .B(B[29]), .Y(n55) );
  NOR2XL U239 ( .A(A[0]), .B(B[0]), .Y(n15) );
endmodule


module hash_core_DW01_add_34 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205;

  OAI211X1 U2 ( .A0(n93), .A1(n94), .B0(n1), .C0(n103), .Y(n89) );
  INVX1 U3 ( .A(n95), .Y(n1) );
  OAI21X1 U4 ( .A0(n55), .A1(n56), .B0(n57), .Y(n51) );
  OAI21X2 U5 ( .A0(n68), .A1(n69), .B0(n70), .Y(n64) );
  NOR2X1 U6 ( .A(n6), .B(n10), .Y(n188) );
  NOR2BX1 U7 ( .AN(n156), .B(n13), .Y(n179) );
  INVXL U8 ( .A(n164), .Y(n181) );
  OAI2BB1XL U9 ( .A0N(n196), .A1N(n38), .B0(n166), .Y(n21) );
  INVXL U10 ( .A(n158), .Y(n196) );
  INVXL U11 ( .A(n51), .Y(n53) );
  INVXL U12 ( .A(n159), .Y(n163) );
  NOR2BX1 U13 ( .AN(n79), .B(n71), .Y(n70) );
  OAI21X1 U14 ( .A0(n117), .A1(n118), .B0(n119), .Y(n114) );
  NOR2XL U15 ( .A(n9), .B(n5), .Y(n189) );
  AOI21XL U16 ( .A0(n152), .A1(n153), .B0(n154), .Y(n150) );
  NAND2XL U17 ( .A(n68), .B(n77), .Y(n86) );
  NAND2XL U18 ( .A(n93), .B(n101), .Y(n112) );
  NOR2XL U19 ( .A(n7), .B(n41), .Y(n204) );
  NOR2XL U20 ( .A(n3), .B(n31), .Y(n205) );
  XNOR2X1 U21 ( .A(n64), .B(n2), .Y(SUM[28]) );
  NAND2X1 U22 ( .A(n67), .B(n65), .Y(n2) );
  NOR2BXL U23 ( .AN(n151), .B(n12), .Y(n171) );
  NAND2XL U24 ( .A(n117), .B(n127), .Y(n140) );
  NAND2XL U25 ( .A(n36), .B(n37), .Y(n34) );
  NAND2XL U26 ( .A(n38), .B(n39), .Y(n36) );
  INVXL U27 ( .A(n134), .Y(n61) );
  NOR2BXL U28 ( .AN(n26), .B(n3), .Y(n25) );
  NOR2BXL U29 ( .AN(n33), .B(n7), .Y(n35) );
  NOR2BXL U30 ( .AN(n20), .B(n5), .Y(n19) );
  NOR2BXL U31 ( .AN(n187), .B(n6), .Y(n194) );
  NOR2BXL U32 ( .AN(n157), .B(n4), .Y(n176) );
  NOR2BXL U33 ( .AN(n44), .B(n8), .Y(n43) );
  NOR2BXL U34 ( .AN(n183), .B(n10), .Y(n191) );
  NOR2BXL U35 ( .AN(n29), .B(n31), .Y(n30) );
  NOR2BXL U36 ( .AN(n155), .B(n169), .Y(n173) );
  NOR2BXL U37 ( .AN(n62), .B(n133), .Y(n132) );
  XOR2XL U38 ( .A(n63), .B(n56), .Y(SUM[29]) );
  NAND2XL U39 ( .A(B[24]), .B(A[24]), .Y(n77) );
  OR2XL U40 ( .A(A[25]), .B(B[25]), .Y(n81) );
  NOR2XL U41 ( .A(A[27]), .B(B[27]), .Y(n16) );
  NAND2XL U42 ( .A(B[26]), .B(A[26]), .Y(n73) );
  NAND2XL U43 ( .A(B[25]), .B(A[25]), .Y(n78) );
  NAND2XL U44 ( .A(B[27]), .B(A[27]), .Y(n79) );
  OR2XL U45 ( .A(A[26]), .B(B[26]), .Y(n80) );
  OR2XL U46 ( .A(A[24]), .B(B[24]), .Y(n90) );
  NAND2XL U47 ( .A(B[28]), .B(A[28]), .Y(n67) );
  OR2XL U48 ( .A(A[28]), .B(B[28]), .Y(n65) );
  INVX1 U49 ( .A(n21), .Y(n180) );
  NOR3X1 U50 ( .A(n166), .B(n160), .C(n159), .Y(n165) );
  NAND3X1 U51 ( .A(n146), .B(n147), .C(n148), .Y(n142) );
  INVX1 U52 ( .A(n149), .Y(n148) );
  NAND3BX1 U53 ( .AN(n158), .B(n161), .C(n162), .Y(n147) );
  AOI21X1 U54 ( .A0(n163), .A1(n164), .B0(n165), .Y(n146) );
  NOR2X1 U55 ( .A(n159), .B(n160), .Y(n161) );
  OAI21XL U56 ( .A0(n180), .A1(n160), .B0(n181), .Y(n178) );
  INVX1 U57 ( .A(n200), .Y(n38) );
  AOI21X1 U58 ( .A0(n81), .A1(n86), .B0(n87), .Y(n84) );
  INVX1 U59 ( .A(n78), .Y(n87) );
  AOI21X1 U60 ( .A0(n64), .A1(n65), .B0(n66), .Y(n56) );
  INVX1 U61 ( .A(n67), .Y(n66) );
  INVX1 U62 ( .A(n152), .Y(n169) );
  INVX1 U63 ( .A(n27), .Y(n31) );
  NAND3BX1 U64 ( .AN(n14), .B(n104), .C(n105), .Y(n94) );
  NAND3BX1 U65 ( .AN(n15), .B(n130), .C(n131), .Y(n118) );
  NOR2X1 U66 ( .A(n120), .B(n121), .Y(n119) );
  INVX1 U67 ( .A(n129), .Y(n120) );
  OAI21XL U68 ( .A0(n182), .A1(n10), .B0(n183), .Y(n164) );
  AOI21X1 U69 ( .A0(n184), .A1(n185), .B0(n186), .Y(n182) );
  INVX1 U70 ( .A(n187), .Y(n186) );
  NAND2X1 U71 ( .A(n20), .B(n23), .Y(n185) );
  NAND3BX1 U72 ( .AN(n16), .B(n80), .C(n81), .Y(n69) );
  INVX1 U73 ( .A(n58), .Y(n55) );
  AOI21X1 U74 ( .A0(n197), .A1(n198), .B0(n199), .Y(n166) );
  AOI21X1 U75 ( .A0(n33), .A1(n37), .B0(n7), .Y(n197) );
  NOR2X1 U76 ( .A(n3), .B(n31), .Y(n198) );
  OAI21XL U77 ( .A0(n3), .A1(n29), .B0(n26), .Y(n199) );
  NAND2X1 U78 ( .A(n188), .B(n189), .Y(n160) );
  INVX1 U79 ( .A(n60), .Y(n133) );
  AOI21X1 U80 ( .A0(n62), .A1(n134), .B0(n133), .Y(n201) );
  NAND2X1 U81 ( .A(n167), .B(n168), .Y(n159) );
  NOR2X1 U82 ( .A(n4), .B(n13), .Y(n167) );
  NOR2X1 U83 ( .A(n12), .B(n169), .Y(n168) );
  NAND2X1 U84 ( .A(n89), .B(n90), .Y(n68) );
  NAND2X1 U85 ( .A(n142), .B(n143), .Y(n117) );
  NAND2X1 U86 ( .A(n114), .B(n115), .Y(n93) );
  NOR2X1 U87 ( .A(n5), .B(n6), .Y(n184) );
  OAI21XL U88 ( .A0(n150), .A1(n12), .B0(n151), .Y(n149) );
  INVX1 U89 ( .A(n155), .Y(n154) );
  OAI21XL U90 ( .A0(n4), .A1(n156), .B0(n157), .Y(n153) );
  NAND2X1 U91 ( .A(n111), .B(n102), .Y(n109) );
  NAND2X1 U92 ( .A(n105), .B(n112), .Y(n111) );
  INVX1 U93 ( .A(n200), .Y(n162) );
  AOI21X1 U94 ( .A0(n201), .A1(n202), .B0(n203), .Y(n200) );
  NOR2X1 U95 ( .A(n8), .B(n11), .Y(n202) );
  OAI21XL U96 ( .A0(n8), .A1(n46), .B0(n44), .Y(n203) );
  NAND2X1 U97 ( .A(n204), .B(n205), .Y(n158) );
  XOR2X1 U98 ( .A(n85), .B(n84), .Y(SUM[26]) );
  NAND2X1 U99 ( .A(n73), .B(n80), .Y(n85) );
  XOR2X1 U100 ( .A(n82), .B(n83), .Y(SUM[27]) );
  NOR2BX1 U101 ( .AN(n79), .B(n16), .Y(n83) );
  OAI21XL U102 ( .A0(n84), .A1(n74), .B0(n73), .Y(n82) );
  XOR2X1 U103 ( .A(n106), .B(n107), .Y(SUM[23]) );
  NOR2BX1 U104 ( .AN(n103), .B(n14), .Y(n107) );
  OAI21XL U105 ( .A0(n108), .A1(n98), .B0(n97), .Y(n106) );
  INVX1 U106 ( .A(n109), .Y(n108) );
  NAND2X1 U107 ( .A(n49), .B(n50), .Y(n48) );
  NAND2X1 U108 ( .A(n51), .B(n52), .Y(n50) );
  OAI21XL U109 ( .A0(n5), .A1(n195), .B0(n20), .Y(n193) );
  INVX1 U110 ( .A(n18), .Y(n195) );
  OAI21XL U111 ( .A0(n9), .A1(n180), .B0(n23), .Y(n18) );
  OAI21XL U112 ( .A0(n13), .A1(n177), .B0(n156), .Y(n175) );
  INVX1 U113 ( .A(n178), .Y(n177) );
  INVX1 U114 ( .A(n130), .Y(n124) );
  INVX1 U115 ( .A(n104), .Y(n98) );
  OAI21XL U116 ( .A0(n32), .A1(n7), .B0(n33), .Y(n28) );
  INVX1 U117 ( .A(n34), .Y(n32) );
  INVX1 U118 ( .A(n105), .Y(n100) );
  INVX1 U119 ( .A(n131), .Y(n126) );
  OAI21XL U120 ( .A0(n192), .A1(n6), .B0(n187), .Y(n190) );
  INVX1 U121 ( .A(n193), .Y(n192) );
  INVX1 U122 ( .A(n39), .Y(n41) );
  OAI21XL U123 ( .A0(n137), .A1(n124), .B0(n123), .Y(n135) );
  INVX1 U124 ( .A(n138), .Y(n137) );
  AOI21X1 U125 ( .A0(n96), .A1(n97), .B0(n14), .Y(n95) );
  NAND2BX1 U126 ( .AN(n98), .B(n99), .Y(n96) );
  OAI21XL U127 ( .A0(n100), .A1(n101), .B0(n102), .Y(n99) );
  AOI21X1 U128 ( .A0(n122), .A1(n123), .B0(n15), .Y(n121) );
  NAND2BX1 U129 ( .AN(n124), .B(n125), .Y(n122) );
  OAI21XL U130 ( .A0(n126), .A1(n127), .B0(n128), .Y(n125) );
  XOR2X1 U131 ( .A(n170), .B(n171), .Y(SUM[15]) );
  OAI2BB1X1 U132 ( .A0N(n152), .A1N(n172), .B0(n155), .Y(n170) );
  OAI2BB1X1 U133 ( .A0N(n131), .A1N(n140), .B0(n128), .Y(n138) );
  OAI21XL U134 ( .A0(n174), .A1(n4), .B0(n157), .Y(n172) );
  INVX1 U135 ( .A(n175), .Y(n174) );
  OAI2BB1X1 U136 ( .A0N(n27), .A1N(n28), .B0(n29), .Y(n24) );
  XOR2X1 U137 ( .A(n89), .B(n91), .Y(SUM[24]) );
  NOR2BX1 U138 ( .AN(n77), .B(n92), .Y(n91) );
  INVX1 U139 ( .A(n90), .Y(n92) );
  XOR2X1 U140 ( .A(n86), .B(n88), .Y(SUM[25]) );
  NOR2BX1 U141 ( .AN(n78), .B(n76), .Y(n88) );
  XOR2X1 U142 ( .A(n140), .B(n141), .Y(SUM[17]) );
  NOR2BX1 U143 ( .AN(n128), .B(n126), .Y(n141) );
  OAI21XL U144 ( .A0(n45), .A1(n11), .B0(n46), .Y(n42) );
  INVX1 U145 ( .A(n47), .Y(n45) );
  OAI2BB1X1 U146 ( .A0N(n60), .A1N(n61), .B0(n62), .Y(n47) );
  INVX1 U147 ( .A(n81), .Y(n76) );
  NOR2BX1 U148 ( .AN(n46), .B(n11), .Y(n59) );
  AOI21X1 U149 ( .A0(n72), .A1(n73), .B0(n16), .Y(n71) );
  NAND2BX1 U150 ( .AN(n74), .B(n75), .Y(n72) );
  OAI21XL U151 ( .A0(n76), .A1(n77), .B0(n78), .Y(n75) );
  INVX1 U152 ( .A(n80), .Y(n74) );
  XOR2X1 U153 ( .A(n142), .B(n144), .Y(SUM[16]) );
  NOR2BX1 U154 ( .AN(n127), .B(n145), .Y(n144) );
  INVX1 U155 ( .A(n143), .Y(n145) );
  NOR2BX1 U156 ( .AN(n23), .B(n9), .Y(n22) );
  NOR2BX1 U157 ( .AN(n97), .B(n98), .Y(n110) );
  NOR2BX1 U158 ( .AN(n123), .B(n124), .Y(n139) );
  NOR2BX1 U159 ( .AN(n129), .B(n15), .Y(n136) );
  NOR2BX1 U160 ( .AN(n102), .B(n100), .Y(n113) );
  NOR2BX1 U161 ( .AN(n37), .B(n41), .Y(n40) );
  NAND2X1 U162 ( .A(n49), .B(n52), .Y(n54) );
  NAND2X1 U163 ( .A(n57), .B(n58), .Y(n63) );
  AND2X2 U164 ( .A(n101), .B(n115), .Y(n116) );
  XOR2X1 U165 ( .A(n135), .B(n136), .Y(SUM[19]) );
  XOR2X1 U166 ( .A(n53), .B(n54), .Y(SUM[30]) );
  XOR2X1 U167 ( .A(n109), .B(n110), .Y(SUM[22]) );
  XOR2X1 U168 ( .A(n112), .B(n113), .Y(SUM[21]) );
  XOR2X1 U169 ( .A(n114), .B(n116), .Y(SUM[20]) );
  XOR2X1 U170 ( .A(n138), .B(n139), .Y(SUM[18]) );
  XOR3X2 U171 ( .A(B[31]), .B(A[31]), .C(n48), .Y(SUM[31]) );
  XOR2X1 U172 ( .A(n175), .B(n176), .Y(SUM[13]) );
  XOR2X1 U173 ( .A(n28), .B(n30), .Y(SUM[6]) );
  XOR2X1 U174 ( .A(n38), .B(n40), .Y(SUM[4]) );
  XOR2X1 U175 ( .A(n24), .B(n25), .Y(SUM[7]) );
  XOR2X1 U176 ( .A(n42), .B(n43), .Y(SUM[3]) );
  XOR2X1 U177 ( .A(n172), .B(n173), .Y(SUM[14]) );
  XOR2X1 U178 ( .A(n190), .B(n191), .Y(SUM[11]) );
  XOR2X1 U179 ( .A(n21), .B(n22), .Y(SUM[8]) );
  XOR2X1 U180 ( .A(n61), .B(n132), .Y(SUM[1]) );
  NOR2BX1 U181 ( .AN(n134), .B(n17), .Y(SUM[0]) );
  XOR2X1 U182 ( .A(n193), .B(n194), .Y(SUM[10]) );
  XOR2X1 U183 ( .A(n18), .B(n19), .Y(SUM[9]) );
  XOR2X1 U184 ( .A(n47), .B(n59), .Y(SUM[2]) );
  XOR2X1 U185 ( .A(n178), .B(n179), .Y(SUM[12]) );
  XOR2X1 U186 ( .A(n34), .B(n35), .Y(SUM[5]) );
  NOR2XL U187 ( .A(A[7]), .B(B[7]), .Y(n3) );
  NOR2XL U188 ( .A(A[13]), .B(B[13]), .Y(n4) );
  NOR2XL U189 ( .A(A[9]), .B(B[9]), .Y(n5) );
  NOR2XL U190 ( .A(A[10]), .B(B[10]), .Y(n6) );
  NOR2XL U191 ( .A(A[5]), .B(B[5]), .Y(n7) );
  NOR2XL U192 ( .A(A[3]), .B(B[3]), .Y(n8) );
  NOR2XL U193 ( .A(A[8]), .B(B[8]), .Y(n9) );
  NOR2XL U194 ( .A(A[11]), .B(B[11]), .Y(n10) );
  NOR2XL U195 ( .A(A[2]), .B(B[2]), .Y(n11) );
  NOR2XL U196 ( .A(A[15]), .B(B[15]), .Y(n12) );
  NOR2XL U197 ( .A(A[12]), .B(B[12]), .Y(n13) );
  OR2XL U198 ( .A(A[6]), .B(B[6]), .Y(n27) );
  NOR2XL U199 ( .A(A[23]), .B(B[23]), .Y(n14) );
  NAND2XL U200 ( .A(B[16]), .B(A[16]), .Y(n127) );
  NAND2XL U201 ( .A(B[18]), .B(A[18]), .Y(n123) );
  NAND2XL U202 ( .A(B[4]), .B(A[4]), .Y(n37) );
  NAND2XL U203 ( .A(B[5]), .B(A[5]), .Y(n33) );
  NAND2XL U204 ( .A(B[12]), .B(A[12]), .Y(n156) );
  NAND2XL U205 ( .A(B[6]), .B(A[6]), .Y(n29) );
  NAND2XL U206 ( .A(B[17]), .B(A[17]), .Y(n128) );
  NAND2XL U207 ( .A(B[13]), .B(A[13]), .Y(n157) );
  NAND2XL U208 ( .A(B[10]), .B(A[10]), .Y(n187) );
  OR2XL U209 ( .A(A[21]), .B(B[21]), .Y(n105) );
  NAND2XL U210 ( .A(B[15]), .B(A[15]), .Y(n151) );
  OR2XL U211 ( .A(A[17]), .B(B[17]), .Y(n131) );
  OR2XL U212 ( .A(A[16]), .B(B[16]), .Y(n143) );
  OR2XL U213 ( .A(A[4]), .B(B[4]), .Y(n39) );
  OR2XL U214 ( .A(A[18]), .B(B[18]), .Y(n130) );
  OR2XL U215 ( .A(A[22]), .B(B[22]), .Y(n104) );
  NOR2XL U216 ( .A(A[19]), .B(B[19]), .Y(n15) );
  NAND2XL U217 ( .A(B[20]), .B(A[20]), .Y(n101) );
  NAND2XL U218 ( .A(B[22]), .B(A[22]), .Y(n97) );
  NAND2XL U219 ( .A(B[21]), .B(A[21]), .Y(n102) );
  NAND2XL U220 ( .A(B[23]), .B(A[23]), .Y(n103) );
  NAND2XL U221 ( .A(B[19]), .B(A[19]), .Y(n129) );
  OR2XL U222 ( .A(A[20]), .B(B[20]), .Y(n115) );
  NAND2X1 U223 ( .A(B[30]), .B(A[30]), .Y(n49) );
  NAND2X1 U224 ( .A(B[29]), .B(A[29]), .Y(n57) );
  OR2X2 U225 ( .A(A[30]), .B(B[30]), .Y(n52) );
  OR2X2 U226 ( .A(A[29]), .B(B[29]), .Y(n58) );
  NOR2XL U227 ( .A(A[0]), .B(B[0]), .Y(n17) );
  NAND2XL U228 ( .A(B[9]), .B(A[9]), .Y(n20) );
  NAND2XL U229 ( .A(B[8]), .B(A[8]), .Y(n23) );
  NAND2XL U230 ( .A(B[14]), .B(A[14]), .Y(n155) );
  OR2XL U231 ( .A(A[14]), .B(B[14]), .Y(n152) );
  NAND2XL U232 ( .A(B[3]), .B(A[3]), .Y(n44) );
  NAND2XL U233 ( .A(B[2]), .B(A[2]), .Y(n46) );
  NAND2XL U234 ( .A(B[11]), .B(A[11]), .Y(n183) );
  NAND2XL U235 ( .A(B[7]), .B(A[7]), .Y(n26) );
  NAND2XL U236 ( .A(B[1]), .B(A[1]), .Y(n62) );
  OR2XL U237 ( .A(A[1]), .B(B[1]), .Y(n60) );
  NAND2XL U238 ( .A(B[0]), .B(A[0]), .Y(n134) );
endmodule


module hash_core_DW01_add_27 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223;

  NOR2X2 U2 ( .A(n168), .B(n169), .Y(n161) );
  AOI21X1 U3 ( .A0(n161), .A1(n162), .B0(n163), .Y(n160) );
  NAND2X2 U4 ( .A(n88), .B(n84), .Y(n87) );
  NAND2BX2 U5 ( .AN(n172), .B(n173), .Y(n159) );
  OAI21X1 U6 ( .A0(n174), .A1(n170), .B0(n175), .Y(n173) );
  NAND4BBX2 U7 ( .AN(n32), .BN(n10), .C(n30), .D(n24), .Y(n179) );
  INVX1 U8 ( .A(n215), .Y(n32) );
  NAND2X2 U9 ( .A(B[6]), .B(A[6]), .Y(n27) );
  OR2X4 U10 ( .A(A[15]), .B(B[15]), .Y(n182) );
  NAND2X4 U11 ( .A(B[7]), .B(A[7]), .Y(n22) );
  OR2X4 U12 ( .A(A[7]), .B(B[7]), .Y(n24) );
  AOI21X2 U13 ( .A0(n171), .A1(n176), .B0(n177), .Y(n174) );
  INVX4 U14 ( .A(n176), .Y(n218) );
  OAI21X4 U15 ( .A0(n220), .A1(n221), .B0(n40), .Y(n176) );
  NAND2X2 U16 ( .A(n5), .B(n96), .Y(n71) );
  OAI21X2 U17 ( .A0(n99), .A1(n100), .B0(n101), .Y(n5) );
  OR2X2 U18 ( .A(A[6]), .B(B[6]), .Y(n30) );
  INVX1 U19 ( .A(n112), .Y(n111) );
  NAND2X2 U20 ( .A(n71), .B(n94), .Y(n92) );
  NAND2X2 U21 ( .A(n126), .B(n127), .Y(n122) );
  NAND3BX1 U22 ( .AN(n128), .B(n129), .C(n130), .Y(n127) );
  NAND2X1 U23 ( .A(B[4]), .B(A[4]), .Y(n36) );
  NAND2X1 U24 ( .A(n16), .B(n204), .Y(n212) );
  OR2X2 U25 ( .A(n2), .B(n3), .Y(n192) );
  NOR2X1 U26 ( .A(A[13]), .B(B[13]), .Y(n11) );
  OAI21XL U27 ( .A0(n190), .A1(n191), .B0(n165), .Y(n188) );
  INVX1 U28 ( .A(n192), .Y(n191) );
  OAI2BB1X1 U29 ( .A0N(n188), .A1N(n1), .B0(n166), .Y(n186) );
  INVX1 U30 ( .A(n11), .Y(n1) );
  INVX1 U31 ( .A(n181), .Y(n169) );
  INVX1 U32 ( .A(n149), .Y(n131) );
  OAI21XL U33 ( .A0(n153), .A1(n139), .B0(n141), .Y(n150) );
  AOI21X2 U34 ( .A0(n74), .A1(n75), .B0(n76), .Y(n73) );
  XOR2X4 U35 ( .A(n114), .B(n115), .Y(SUM[23]) );
  OAI21X2 U36 ( .A0(n116), .A1(n111), .B0(n109), .Y(n114) );
  INVX2 U37 ( .A(n117), .Y(n116) );
  NAND2X4 U38 ( .A(n122), .B(n123), .Y(n99) );
  AOI21X2 U39 ( .A0(n102), .A1(n103), .B0(n104), .Y(n101) );
  NOR2XL U40 ( .A(n194), .B(n170), .Y(n2) );
  INVXL U41 ( .A(n175), .Y(n3) );
  INVX1 U42 ( .A(n16), .Y(n194) );
  NAND4BBX2 U43 ( .AN(n19), .BN(n15), .C(n198), .D(n197), .Y(n170) );
  OAI2BB1X4 U44 ( .A0N(n195), .A1N(n196), .B0(n197), .Y(n175) );
  OR2XL U45 ( .A(n218), .B(n179), .Y(n4) );
  NAND2X4 U46 ( .A(n4), .B(n178), .Y(n16) );
  OAI2BB1X2 U47 ( .A0N(n213), .A1N(n214), .B0(n24), .Y(n178) );
  NAND2X4 U48 ( .A(n159), .B(n160), .Y(n129) );
  OAI21X4 U49 ( .A0(n58), .A1(n59), .B0(n60), .Y(n49) );
  INVX4 U50 ( .A(n69), .Y(n59) );
  NAND2XL U51 ( .A(B[18]), .B(A[18]), .Y(n142) );
  NOR2X1 U52 ( .A(A[4]), .B(B[4]), .Y(n10) );
  NOR2BX1 U53 ( .AN(n109), .B(n111), .Y(n118) );
  OR2X2 U54 ( .A(A[8]), .B(B[8]), .Y(n204) );
  NOR2BXL U55 ( .AN(n108), .B(n106), .Y(n121) );
  OR2XL U56 ( .A(A[2]), .B(B[2]), .Y(n63) );
  NAND2X1 U57 ( .A(B[8]), .B(A[8]), .Y(n18) );
  NOR2BX1 U58 ( .AN(n54), .B(n8), .Y(n48) );
  OR2X1 U59 ( .A(A[12]), .B(B[12]), .Y(n180) );
  OR2XL U60 ( .A(A[20]), .B(B[20]), .Y(n123) );
  OAI21XL U61 ( .A0(n31), .A1(n32), .B0(n33), .Y(n28) );
  NAND2X1 U62 ( .A(n91), .B(n92), .Y(n90) );
  NAND2X1 U63 ( .A(n14), .B(n18), .Y(n200) );
  NAND2X1 U64 ( .A(n33), .B(n36), .Y(n216) );
  INVX1 U65 ( .A(n182), .Y(n168) );
  NAND2X1 U66 ( .A(B[2]), .B(A[2]), .Y(n44) );
  OAI21XL U67 ( .A0(n145), .A1(n146), .B0(n66), .Y(n223) );
  INVX1 U68 ( .A(n134), .Y(n139) );
  INVX1 U69 ( .A(n119), .Y(n106) );
  OR2X2 U70 ( .A(A[11]), .B(B[11]), .Y(n197) );
  NAND2X1 U71 ( .A(B[14]), .B(A[14]), .Y(n167) );
  NAND2X4 U72 ( .A(B[0]), .B(A[0]), .Y(n146) );
  NAND2X1 U73 ( .A(B[12]), .B(A[12]), .Y(n165) );
  NOR2X1 U74 ( .A(A[30]), .B(B[30]), .Y(n51) );
  NAND2X1 U75 ( .A(A[24]), .B(B[24]), .Y(n79) );
  INVXL U76 ( .A(n219), .Y(n41) );
  OAI21X2 U77 ( .A0(n71), .A1(n72), .B0(n73), .Y(n69) );
  NAND3BXL U78 ( .AN(n78), .B(n84), .C(n83), .Y(n72) );
  INVX2 U79 ( .A(n199), .Y(n15) );
  NOR2BXL U80 ( .AN(n86), .B(n82), .Y(n89) );
  XOR2XL U81 ( .A(n70), .B(n59), .Y(SUM[28]) );
  NAND2XL U82 ( .A(n60), .B(n61), .Y(n70) );
  XNOR2X1 U83 ( .A(n6), .B(n67), .Y(SUM[29]) );
  NAND2X1 U84 ( .A(n60), .B(n68), .Y(n6) );
  XNOR2X1 U85 ( .A(n7), .B(n85), .Y(SUM[27]) );
  NAND2X1 U86 ( .A(n86), .B(n87), .Y(n7) );
  NAND2XL U87 ( .A(n69), .B(n61), .Y(n68) );
  NAND2XL U88 ( .A(B[1]), .B(A[1]), .Y(n66) );
  NAND2XL U89 ( .A(B[3]), .B(A[3]), .Y(n40) );
  NAND2XL U90 ( .A(n99), .B(n107), .Y(n120) );
  NOR2BXL U91 ( .AN(n167), .B(n169), .Y(n187) );
  NOR2BXL U92 ( .AN(n164), .B(n168), .Y(n184) );
  NAND2XL U93 ( .A(n138), .B(n143), .Y(n147) );
  INVXL U94 ( .A(n96), .Y(n98) );
  NOR2BXL U95 ( .AN(n105), .B(n110), .Y(n115) );
  NOR2BXL U96 ( .AN(n80), .B(n78), .Y(n93) );
  NAND2XL U97 ( .A(n129), .B(n133), .Y(n156) );
  NOR2BXL U98 ( .AN(n142), .B(n131), .Y(n152) );
  INVXL U99 ( .A(n198), .Y(n210) );
  NAND2XL U100 ( .A(n197), .B(n203), .Y(n205) );
  AOI21XL U101 ( .A0(n198), .A1(n207), .B0(n208), .Y(n206) );
  INVXL U102 ( .A(n201), .Y(n208) );
  NOR2BXL U103 ( .AN(n141), .B(n139), .Y(n155) );
  NAND2XL U104 ( .A(n133), .B(n134), .Y(n128) );
  NOR2BXL U105 ( .AN(n18), .B(n19), .Y(n17) );
  NOR2BXL U106 ( .AN(n165), .B(n190), .Y(n193) );
  NOR2BXL U107 ( .AN(n14), .B(n15), .Y(n13) );
  INVXL U108 ( .A(n133), .Y(n158) );
  NAND2XL U109 ( .A(B[13]), .B(A[13]), .Y(n166) );
  NAND2XL U110 ( .A(B[15]), .B(A[15]), .Y(n164) );
  NAND2XL U111 ( .A(B[27]), .B(A[27]), .Y(n77) );
  NAND2XL U112 ( .A(B[23]), .B(A[23]), .Y(n105) );
  NAND2XL U113 ( .A(B[25]), .B(A[25]), .Y(n80) );
  NAND2XL U114 ( .A(B[21]), .B(A[21]), .Y(n108) );
  NAND2XL U115 ( .A(B[17]), .B(A[17]), .Y(n141) );
  NAND2XL U116 ( .A(B[22]), .B(A[22]), .Y(n109) );
  NAND2XL U117 ( .A(B[30]), .B(A[30]), .Y(n53) );
  NOR2XL U118 ( .A(A[25]), .B(B[25]), .Y(n78) );
  NAND2XL U119 ( .A(B[26]), .B(A[26]), .Y(n81) );
  NOR2XL U120 ( .A(A[30]), .B(B[30]), .Y(n8) );
  NAND2XL U121 ( .A(B[28]), .B(A[28]), .Y(n60) );
  NAND2XL U122 ( .A(B[29]), .B(A[29]), .Y(n56) );
  NAND2XL U123 ( .A(B[24]), .B(A[24]), .Y(n94) );
  NAND2XL U124 ( .A(B[26]), .B(A[26]), .Y(n86) );
  NOR2BX1 U125 ( .AN(n146), .B(n9), .Y(SUM[0]) );
  NOR2XL U126 ( .A(A[0]), .B(B[0]), .Y(n9) );
  AOI21XL U127 ( .A0(n48), .A1(n49), .B0(n50), .Y(n47) );
  INVX1 U128 ( .A(n28), .Y(n25) );
  INVX1 U129 ( .A(n45), .Y(n42) );
  NAND2X1 U130 ( .A(n63), .B(n219), .Y(n221) );
  NOR2X1 U131 ( .A(n222), .B(n223), .Y(n220) );
  INVX1 U132 ( .A(n44), .Y(n222) );
  INVX1 U133 ( .A(n178), .Y(n177) );
  INVX1 U134 ( .A(n179), .Y(n171) );
  NOR2X1 U135 ( .A(n110), .B(n111), .Y(n102) );
  NOR2X1 U136 ( .A(n132), .B(n131), .Y(n135) );
  NOR2X1 U137 ( .A(n131), .B(n132), .Y(n130) );
  OAI21XL U138 ( .A0(n10), .A1(n218), .B0(n36), .Y(n34) );
  INVX1 U139 ( .A(n34), .Y(n31) );
  INVX1 U140 ( .A(n64), .Y(n145) );
  INVX1 U141 ( .A(n30), .Y(n26) );
  XOR2X1 U142 ( .A(n34), .B(n35), .Y(SUM[5]) );
  NOR2BX1 U143 ( .AN(n33), .B(n32), .Y(n35) );
  XOR2X1 U144 ( .A(n28), .B(n29), .Y(SUM[6]) );
  NOR2BX1 U145 ( .AN(n27), .B(n26), .Y(n29) );
  XOR2X1 U146 ( .A(n176), .B(n37), .Y(SUM[4]) );
  NOR2BX1 U147 ( .AN(n36), .B(n10), .Y(n37) );
  INVX1 U148 ( .A(n63), .Y(n43) );
  OAI2BB1X1 U149 ( .A0N(n64), .A1N(n65), .B0(n66), .Y(n45) );
  XOR2X1 U150 ( .A(n65), .B(n144), .Y(SUM[1]) );
  NOR2BX1 U151 ( .AN(n66), .B(n145), .Y(n144) );
  XOR2X1 U152 ( .A(n45), .B(n62), .Y(SUM[2]) );
  NOR2BX1 U153 ( .AN(n44), .B(n43), .Y(n62) );
  XOR2X1 U154 ( .A(n38), .B(n39), .Y(SUM[3]) );
  NOR2BX1 U155 ( .AN(n40), .B(n41), .Y(n39) );
  OAI21XL U156 ( .A0(n42), .A1(n43), .B0(n44), .Y(n38) );
  OAI211X1 U157 ( .A0(n11), .A1(n165), .B0(n166), .C0(n167), .Y(n162) );
  INVX1 U158 ( .A(n61), .Y(n58) );
  OAI21XL U159 ( .A0(n99), .A1(n100), .B0(n101), .Y(n95) );
  NAND3BX1 U160 ( .AN(n106), .B(n112), .C(n113), .Y(n100) );
  INVX1 U161 ( .A(n105), .Y(n104) );
  OAI211X1 U162 ( .A0(n78), .A1(n79), .B0(n80), .C0(n81), .Y(n75) );
  NAND2X1 U163 ( .A(n90), .B(n80), .Y(n88) );
  AOI21X1 U164 ( .A0(n135), .A1(n136), .B0(n137), .Y(n126) );
  INVX1 U165 ( .A(n138), .Y(n137) );
  NAND3X1 U166 ( .A(n198), .B(n199), .C(n200), .Y(n196) );
  NOR2BX1 U167 ( .AN(n201), .B(n202), .Y(n195) );
  NAND4BXL U168 ( .AN(n11), .B(n180), .C(n181), .D(n182), .Y(n172) );
  INVX1 U169 ( .A(n203), .Y(n202) );
  NAND2X1 U170 ( .A(n77), .B(n83), .Y(n85) );
  OAI211X1 U171 ( .A0(n139), .A1(n140), .B0(n141), .C0(n142), .Y(n136) );
  OAI211X1 U172 ( .A0(n106), .A1(n107), .B0(n108), .C0(n109), .Y(n103) );
  INVX1 U173 ( .A(n154), .Y(n153) );
  NAND2X1 U174 ( .A(B[5]), .B(A[5]), .Y(n33) );
  INVX1 U175 ( .A(n84), .Y(n82) );
  INVX1 U176 ( .A(n113), .Y(n110) );
  INVX1 U177 ( .A(n143), .Y(n132) );
  INVX1 U178 ( .A(n204), .Y(n19) );
  NAND2X1 U179 ( .A(n156), .B(n140), .Y(n154) );
  OAI2BB1X1 U180 ( .A0N(n119), .A1N(n120), .B0(n108), .Y(n117) );
  NAND3X1 U181 ( .A(n215), .B(n30), .C(n216), .Y(n214) );
  NOR2BX1 U182 ( .AN(n27), .B(n217), .Y(n213) );
  NOR2BX1 U183 ( .AN(n83), .B(n82), .Y(n74) );
  OR2X2 U184 ( .A(A[5]), .B(B[5]), .Y(n215) );
  INVX1 U185 ( .A(n22), .Y(n217) );
  INVX1 U186 ( .A(n164), .Y(n163) );
  XOR2X1 U187 ( .A(n150), .B(n152), .Y(SUM[18]) );
  XOR2X1 U188 ( .A(n95), .B(n97), .Y(SUM[24]) );
  NOR2BX1 U189 ( .AN(n94), .B(n98), .Y(n97) );
  XOR2X1 U190 ( .A(n147), .B(n148), .Y(SUM[19]) );
  AOI21X1 U191 ( .A0(n149), .A1(n150), .B0(n151), .Y(n148) );
  INVX1 U192 ( .A(n142), .Y(n151) );
  XOR2X1 U193 ( .A(n117), .B(n118), .Y(SUM[22]) );
  XOR2X1 U194 ( .A(n183), .B(n184), .Y(SUM[15]) );
  OAI21XL U195 ( .A0(n185), .A1(n169), .B0(n167), .Y(n183) );
  INVX1 U196 ( .A(n186), .Y(n185) );
  XOR2X1 U197 ( .A(n120), .B(n121), .Y(SUM[21]) );
  XOR2X1 U198 ( .A(n88), .B(n89), .Y(SUM[26]) );
  XOR2X1 U199 ( .A(n92), .B(n93), .Y(SUM[25]) );
  NAND2X1 U200 ( .A(n54), .B(n56), .Y(n67) );
  OAI21XL U201 ( .A0(n211), .A1(n15), .B0(n14), .Y(n207) );
  INVX1 U202 ( .A(n12), .Y(n211) );
  INVX1 U203 ( .A(n180), .Y(n190) );
  XOR2X1 U204 ( .A(n20), .B(n21), .Y(SUM[7]) );
  NOR2BX1 U205 ( .AN(n22), .B(n23), .Y(n21) );
  OAI21XL U206 ( .A0(n25), .A1(n26), .B0(n27), .Y(n20) );
  INVX1 U207 ( .A(n24), .Y(n23) );
  NAND2X1 U208 ( .A(n212), .B(n18), .Y(n12) );
  OR2X2 U209 ( .A(A[3]), .B(B[3]), .Y(n219) );
  INVX1 U210 ( .A(n77), .Y(n76) );
  OR2X2 U211 ( .A(A[1]), .B(B[1]), .Y(n64) );
  XOR2X1 U212 ( .A(n207), .B(n209), .Y(SUM[10]) );
  NOR2BX1 U213 ( .AN(n201), .B(n210), .Y(n209) );
  XOR2X1 U214 ( .A(n186), .B(n187), .Y(SUM[14]) );
  XOR2X1 U215 ( .A(n192), .B(n193), .Y(SUM[12]) );
  XOR2X1 U216 ( .A(n188), .B(n189), .Y(SUM[13]) );
  NOR2BX1 U217 ( .AN(n166), .B(n11), .Y(n189) );
  XOR2X1 U218 ( .A(n129), .B(n157), .Y(SUM[16]) );
  NOR2BX1 U219 ( .AN(n140), .B(n158), .Y(n157) );
  XOR2X1 U220 ( .A(n205), .B(n206), .Y(SUM[11]) );
  XOR2X1 U221 ( .A(n154), .B(n155), .Y(SUM[17]) );
  XOR2X1 U222 ( .A(n122), .B(n124), .Y(SUM[20]) );
  NOR2BX1 U223 ( .AN(n107), .B(n125), .Y(n124) );
  INVX1 U224 ( .A(n123), .Y(n125) );
  XOR2X1 U225 ( .A(n16), .B(n17), .Y(SUM[8]) );
  XOR2X1 U226 ( .A(n12), .B(n13), .Y(SUM[9]) );
  INVX1 U227 ( .A(n146), .Y(n65) );
  NAND2X1 U228 ( .A(B[11]), .B(A[11]), .Y(n203) );
  OR2X2 U229 ( .A(A[14]), .B(B[14]), .Y(n181) );
  XOR3X2 U230 ( .A(B[30]), .B(A[30]), .C(n55), .Y(SUM[30]) );
  NAND2X1 U231 ( .A(n56), .B(n57), .Y(n55) );
  NAND2X1 U232 ( .A(n54), .B(n49), .Y(n57) );
  OR2X2 U233 ( .A(A[10]), .B(B[10]), .Y(n198) );
  NAND2X1 U234 ( .A(B[9]), .B(A[9]), .Y(n14) );
  NAND2X1 U235 ( .A(B[10]), .B(A[10]), .Y(n201) );
  OR2X2 U236 ( .A(A[27]), .B(B[27]), .Y(n83) );
  OR2X2 U237 ( .A(A[26]), .B(B[26]), .Y(n84) );
  NAND2X1 U238 ( .A(B[19]), .B(A[19]), .Y(n138) );
  OR2X2 U239 ( .A(A[9]), .B(B[9]), .Y(n199) );
  OR2X2 U240 ( .A(A[18]), .B(B[18]), .Y(n149) );
  OR2X2 U241 ( .A(A[25]), .B(B[25]), .Y(n91) );
  OR2X2 U242 ( .A(A[19]), .B(B[19]), .Y(n143) );
  OR2X2 U243 ( .A(A[17]), .B(B[17]), .Y(n134) );
  OR2X2 U244 ( .A(A[23]), .B(B[23]), .Y(n113) );
  OR2X2 U245 ( .A(A[22]), .B(B[22]), .Y(n112) );
  OR2X2 U246 ( .A(A[21]), .B(B[21]), .Y(n119) );
  NAND2X1 U247 ( .A(B[20]), .B(A[20]), .Y(n107) );
  NAND2X1 U248 ( .A(B[16]), .B(A[16]), .Y(n140) );
  OR2X2 U249 ( .A(A[29]), .B(B[29]), .Y(n54) );
  OR2X2 U250 ( .A(A[16]), .B(B[16]), .Y(n133) );
  OR2X2 U251 ( .A(A[28]), .B(B[28]), .Y(n61) );
  OAI21XL U252 ( .A0(n51), .A1(n52), .B0(n53), .Y(n50) );
  NAND2X1 U253 ( .A(A[29]), .B(B[29]), .Y(n52) );
  OR2X2 U254 ( .A(A[24]), .B(B[24]), .Y(n96) );
  XOR2X1 U255 ( .A(n46), .B(n47), .Y(SUM[31]) );
  XNOR2X1 U256 ( .A(B[31]), .B(A[31]), .Y(n46) );
endmodule


module hash_core_DW01_add_35 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205;

  INVX4 U2 ( .A(n180), .Y(n179) );
  NOR2X2 U3 ( .A(A[2]), .B(B[2]), .Y(n12) );
  OR2X2 U4 ( .A(A[1]), .B(B[1]), .Y(n62) );
  NOR2X1 U5 ( .A(n163), .B(n164), .Y(n165) );
  NOR2BXL U6 ( .AN(n50), .B(n1), .Y(n61) );
  OAI21X2 U7 ( .A0(n11), .A1(n50), .B0(n48), .Y(n203) );
  NAND3X4 U8 ( .A(n150), .B(n151), .C(n152), .Y(n146) );
  XOR2X2 U9 ( .A(n175), .B(n176), .Y(SUM[14]) );
  XOR2X2 U10 ( .A(n34), .B(n36), .Y(SUM[6]) );
  XOR2X4 U11 ( .A(n139), .B(n140), .Y(SUM[19]) );
  OAI21X2 U12 ( .A0(n141), .A1(n128), .B0(n127), .Y(n139) );
  INVX2 U13 ( .A(n193), .Y(n192) );
  OAI21X2 U14 ( .A0(n15), .A1(n3), .B0(n26), .Y(n193) );
  XOR2X4 U15 ( .A(n173), .B(n174), .Y(SUM[15]) );
  XOR2X4 U16 ( .A(n30), .B(n31), .Y(SUM[7]) );
  NAND2X4 U17 ( .A(B[0]), .B(A[0]), .Y(n138) );
  NAND2X2 U18 ( .A(B[5]), .B(A[5]), .Y(n38) );
  BUFX4 U19 ( .A(n12), .Y(n1) );
  OR2X4 U20 ( .A(A[4]), .B(B[4]), .Y(n43) );
  NOR2X2 U21 ( .A(n16), .B(n17), .Y(n188) );
  OR2X2 U22 ( .A(A[18]), .B(B[18]), .Y(n134) );
  OR2X2 U23 ( .A(A[17]), .B(B[17]), .Y(n135) );
  INVXL U24 ( .A(n10), .Y(n5) );
  INVXL U25 ( .A(n14), .Y(n2) );
  NOR2X1 U26 ( .A(n19), .B(n172), .Y(n171) );
  OAI21XL U27 ( .A0(n103), .A1(n104), .B0(n105), .Y(n102) );
  NAND2BX1 U28 ( .AN(n128), .B(n129), .Y(n126) );
  OAI21XL U29 ( .A0(n130), .A1(n131), .B0(n132), .Y(n129) );
  AOI21X1 U30 ( .A0(n64), .A1(n138), .B0(n137), .Y(n201) );
  OAI21XL U31 ( .A0(n13), .A1(n35), .B0(n32), .Y(n199) );
  AOI21X1 U32 ( .A0(n38), .A1(n42), .B0(n10), .Y(n197) );
  NOR2X1 U33 ( .A(n10), .B(n45), .Y(n204) );
  NAND2X1 U34 ( .A(n108), .B(n115), .Y(n114) );
  INVX1 U35 ( .A(n62), .Y(n137) );
  NAND2X1 U36 ( .A(B[2]), .B(A[2]), .Y(n50) );
  NOR2X1 U37 ( .A(A[8]), .B(B[8]), .Y(n18) );
  NAND2X1 U38 ( .A(n6), .B(n169), .Y(n180) );
  NOR2X1 U39 ( .A(A[12]), .B(B[12]), .Y(n20) );
  NOR2X1 U40 ( .A(A[13]), .B(B[13]), .Y(n14) );
  OAI21XL U41 ( .A0(n57), .A1(n58), .B0(n59), .Y(n55) );
  NOR2BX1 U42 ( .AN(n38), .B(n10), .Y(n40) );
  XOR2X2 U43 ( .A(n190), .B(n191), .Y(SUM[11]) );
  OAI21X1 U44 ( .A0(n192), .A1(n16), .B0(n186), .Y(n190) );
  INVX1 U45 ( .A(n142), .Y(n141) );
  INVX1 U46 ( .A(n196), .Y(n168) );
  OAI2BB1X1 U47 ( .A0N(n156), .A1N(n175), .B0(n159), .Y(n173) );
  INVX1 U48 ( .A(n29), .Y(n4) );
  NAND2X1 U49 ( .A(B[8]), .B(A[8]), .Y(n29) );
  NOR2X2 U50 ( .A(A[15]), .B(B[15]), .Y(n19) );
  NOR2X1 U51 ( .A(A[10]), .B(B[10]), .Y(n16) );
  NOR2X4 U52 ( .A(n18), .B(n15), .Y(n189) );
  AOI2BB1X2 U53 ( .A0N(n18), .A1N(n182), .B0(n4), .Y(n3) );
  AOI21X2 U54 ( .A0(n26), .A1(n29), .B0(n16), .Y(n184) );
  OAI2BB1X4 U55 ( .A0N(n195), .A1N(n166), .B0(n196), .Y(n27) );
  OAI21X4 U56 ( .A0(n121), .A1(n122), .B0(n123), .Y(n117) );
  NAND2X4 U57 ( .A(n146), .B(n147), .Y(n121) );
  OAI21X1 U58 ( .A0(n95), .A1(n96), .B0(n97), .Y(n91) );
  OAI2BB1X2 U59 ( .A0N(n39), .A1N(n5), .B0(n38), .Y(n34) );
  NAND2X2 U60 ( .A(n41), .B(n42), .Y(n39) );
  INVXL U61 ( .A(n3), .Y(n24) );
  NOR2X2 U62 ( .A(A[5]), .B(B[5]), .Y(n10) );
  NAND2X1 U63 ( .A(B[3]), .B(A[3]), .Y(n48) );
  OAI2BB1X4 U64 ( .A0N(n177), .A1N(n2), .B0(n161), .Y(n175) );
  OAI21X4 U65 ( .A0(n20), .A1(n179), .B0(n160), .Y(n177) );
  NAND2X1 U66 ( .A(B[10]), .B(A[10]), .Y(n186) );
  XOR2X1 U67 ( .A(n87), .B(n86), .Y(SUM[26]) );
  XOR2X1 U68 ( .A(n180), .B(n181), .Y(SUM[12]) );
  XOR2X2 U69 ( .A(n55), .B(n9), .Y(SUM[30]) );
  XOR2X1 U70 ( .A(n65), .B(n58), .Y(SUM[29]) );
  OR2XL U71 ( .A(n182), .B(n164), .Y(n6) );
  INVX4 U72 ( .A(n27), .Y(n182) );
  NAND2X2 U73 ( .A(n188), .B(n189), .Y(n164) );
  AOI21X2 U74 ( .A0(n183), .A1(n184), .B0(n185), .Y(n169) );
  OAI21XL U75 ( .A0(n154), .A1(n19), .B0(n155), .Y(n153) );
  NAND2X2 U76 ( .A(n117), .B(n118), .Y(n95) );
  NOR2X2 U77 ( .A(A[3]), .B(B[3]), .Y(n11) );
  NAND2X1 U78 ( .A(B[17]), .B(A[17]), .Y(n132) );
  OAI2BB1X1 U79 ( .A0N(n33), .A1N(n34), .B0(n35), .Y(n30) );
  NOR2BXL U80 ( .AN(n32), .B(n13), .Y(n31) );
  NOR2X1 U81 ( .A(n13), .B(n37), .Y(n205) );
  INVX1 U82 ( .A(n43), .Y(n45) );
  INVX2 U83 ( .A(n33), .Y(n37) );
  OAI21XL U84 ( .A0(n14), .A1(n160), .B0(n161), .Y(n157) );
  NOR2X1 U85 ( .A(n124), .B(n125), .Y(n123) );
  NOR2BX1 U86 ( .AN(n106), .B(n22), .Y(n110) );
  NAND2X1 U87 ( .A(n75), .B(n82), .Y(n87) );
  XOR2X1 U88 ( .A(n112), .B(n113), .Y(SUM[22]) );
  NOR2BX1 U89 ( .AN(n100), .B(n101), .Y(n113) );
  OAI21XL U90 ( .A0(n49), .A1(n1), .B0(n50), .Y(n46) );
  XOR2X1 U91 ( .A(n46), .B(n47), .Y(SUM[3]) );
  NOR2X1 U92 ( .A(A[19]), .B(B[19]), .Y(n21) );
  NAND2XL U93 ( .A(B[18]), .B(A[18]), .Y(n127) );
  NAND2X1 U94 ( .A(B[20]), .B(A[20]), .Y(n104) );
  NAND2XL U95 ( .A(B[14]), .B(A[14]), .Y(n159) );
  NAND2X1 U96 ( .A(B[16]), .B(A[16]), .Y(n131) );
  OR2X2 U97 ( .A(A[21]), .B(B[21]), .Y(n108) );
  CLKINVX3 U98 ( .A(n162), .Y(n195) );
  NAND3BXL U99 ( .AN(n162), .B(n165), .C(n166), .Y(n151) );
  NOR2XL U100 ( .A(n164), .B(n163), .Y(n167) );
  NOR2BXL U101 ( .AN(n159), .B(n172), .Y(n176) );
  CLKINVX3 U102 ( .A(n200), .Y(n166) );
  NAND2XL U103 ( .A(n166), .B(n43), .Y(n41) );
  NOR2BX1 U104 ( .AN(n106), .B(n98), .Y(n97) );
  AOI21X2 U105 ( .A0(n83), .A1(n88), .B0(n89), .Y(n86) );
  NOR2BXL U106 ( .AN(n160), .B(n20), .Y(n181) );
  XOR2X2 U107 ( .A(n109), .B(n110), .Y(SUM[23]) );
  OAI21X1 U108 ( .A0(n111), .A1(n101), .B0(n100), .Y(n109) );
  XOR2X2 U109 ( .A(n84), .B(n85), .Y(SUM[27]) );
  OAI21X1 U110 ( .A0(n86), .A1(n76), .B0(n75), .Y(n84) );
  OAI2BB1X2 U111 ( .A0N(n135), .A1N(n144), .B0(n132), .Y(n142) );
  NAND2X2 U112 ( .A(n91), .B(n92), .Y(n70) );
  NAND2X2 U113 ( .A(n114), .B(n105), .Y(n112) );
  NOR2BX1 U114 ( .AN(n81), .B(n73), .Y(n72) );
  NOR2BXL U115 ( .AN(n127), .B(n128), .Y(n143) );
  NOR2BXL U116 ( .AN(n64), .B(n137), .Y(n136) );
  XNOR2X1 U117 ( .A(n66), .B(n7), .Y(SUM[28]) );
  NAND2X1 U118 ( .A(n69), .B(n67), .Y(n7) );
  NOR2X2 U119 ( .A(A[7]), .B(B[7]), .Y(n13) );
  NOR2X2 U120 ( .A(A[9]), .B(B[9]), .Y(n15) );
  NOR2X2 U121 ( .A(A[11]), .B(B[11]), .Y(n17) );
  NAND2XL U122 ( .A(B[7]), .B(A[7]), .Y(n32) );
  NAND2XL U123 ( .A(B[9]), .B(A[9]), .Y(n26) );
  NAND2XL U124 ( .A(B[13]), .B(A[13]), .Y(n161) );
  NAND2XL U125 ( .A(B[11]), .B(A[11]), .Y(n187) );
  OR2X4 U126 ( .A(A[14]), .B(B[14]), .Y(n156) );
  NAND2XL U127 ( .A(B[15]), .B(A[15]), .Y(n155) );
  NAND2XL U128 ( .A(n55), .B(n56), .Y(n54) );
  OR2XL U129 ( .A(A[16]), .B(B[16]), .Y(n147) );
  NAND2XL U130 ( .A(B[22]), .B(A[22]), .Y(n100) );
  NAND2XL U131 ( .A(B[19]), .B(A[19]), .Y(n133) );
  NOR2BX1 U132 ( .AN(n138), .B(n8), .Y(SUM[0]) );
  NOR2XL U133 ( .A(A[0]), .B(B[0]), .Y(n8) );
  OR2XL U134 ( .A(A[20]), .B(B[20]), .Y(n118) );
  AOI2BB2X1 U135 ( .B0(n167), .B1(n168), .A0N(n169), .A1N(n163), .Y(n150) );
  INVX1 U136 ( .A(n153), .Y(n152) );
  XOR2X1 U137 ( .A(n177), .B(n178), .Y(SUM[13]) );
  NOR2BX1 U138 ( .AN(n161), .B(n14), .Y(n178) );
  NOR2BX1 U139 ( .AN(n187), .B(n17), .Y(n191) );
  NOR2BX1 U140 ( .AN(n155), .B(n19), .Y(n174) );
  AOI21X1 U141 ( .A0(n197), .A1(n198), .B0(n199), .Y(n196) );
  NOR2X1 U142 ( .A(n13), .B(n37), .Y(n198) );
  AOI21X1 U143 ( .A0(n201), .A1(n202), .B0(n203), .Y(n200) );
  NOR2X1 U144 ( .A(n11), .B(n1), .Y(n202) );
  NAND2X1 U145 ( .A(n204), .B(n205), .Y(n162) );
  INVX1 U146 ( .A(n80), .Y(n89) );
  NAND3BX1 U147 ( .AN(n22), .B(n107), .C(n108), .Y(n96) );
  NAND3BX1 U148 ( .AN(n21), .B(n134), .C(n135), .Y(n122) );
  INVX1 U149 ( .A(n133), .Y(n124) );
  XOR2X1 U150 ( .A(n88), .B(n90), .Y(SUM[25]) );
  NOR2BX1 U151 ( .AN(n80), .B(n78), .Y(n90) );
  OAI21XL U152 ( .A0(n186), .A1(n17), .B0(n187), .Y(n185) );
  NOR2X1 U153 ( .A(n15), .B(n17), .Y(n183) );
  NAND2X1 U154 ( .A(n170), .B(n171), .Y(n163) );
  NOR2X1 U155 ( .A(n14), .B(n20), .Y(n170) );
  INVX1 U156 ( .A(n156), .Y(n172) );
  NOR2BX1 U157 ( .AN(n133), .B(n21), .Y(n140) );
  NAND2X1 U158 ( .A(n70), .B(n79), .Y(n88) );
  XOR2X1 U159 ( .A(n193), .B(n194), .Y(SUM[10]) );
  NOR2BX1 U160 ( .AN(n186), .B(n16), .Y(n194) );
  XOR2X1 U161 ( .A(n24), .B(n25), .Y(SUM[9]) );
  NOR2BX1 U162 ( .AN(n26), .B(n15), .Y(n25) );
  NOR2BX1 U163 ( .AN(n35), .B(n37), .Y(n36) );
  XOR2X1 U164 ( .A(n166), .B(n44), .Y(SUM[4]) );
  NOR2BX1 U165 ( .AN(n42), .B(n45), .Y(n44) );
  NOR2BX1 U166 ( .AN(n81), .B(n23), .Y(n85) );
  XOR2X1 U167 ( .A(n115), .B(n116), .Y(SUM[21]) );
  NOR2BX1 U168 ( .AN(n105), .B(n103), .Y(n116) );
  XOR2X1 U169 ( .A(n39), .B(n40), .Y(SUM[5]) );
  XOR2X1 U170 ( .A(n27), .B(n28), .Y(SUM[8]) );
  NOR2BX1 U171 ( .AN(n29), .B(n18), .Y(n28) );
  XOR2X1 U172 ( .A(n144), .B(n145), .Y(SUM[17]) );
  NOR2BX1 U173 ( .AN(n132), .B(n130), .Y(n145) );
  XOR2X1 U174 ( .A(n142), .B(n143), .Y(SUM[18]) );
  NAND2X1 U175 ( .A(n95), .B(n104), .Y(n115) );
  AOI21X1 U176 ( .A0(n156), .A1(n157), .B0(n158), .Y(n154) );
  INVX1 U177 ( .A(n159), .Y(n158) );
  NAND2X1 U178 ( .A(n121), .B(n131), .Y(n144) );
  INVX1 U179 ( .A(n112), .Y(n111) );
  AND2X2 U180 ( .A(n53), .B(n56), .Y(n9) );
  AOI21X1 U181 ( .A0(n66), .A1(n67), .B0(n68), .Y(n58) );
  INVX1 U182 ( .A(n69), .Y(n68) );
  OAI21XL U183 ( .A0(n70), .A1(n71), .B0(n72), .Y(n66) );
  NAND3BX1 U184 ( .AN(n23), .B(n82), .C(n83), .Y(n71) );
  INVX1 U185 ( .A(n60), .Y(n57) );
  INVX1 U186 ( .A(n134), .Y(n128) );
  INVX1 U187 ( .A(n107), .Y(n101) );
  XOR2X1 U188 ( .A(n91), .B(n93), .Y(SUM[24]) );
  NOR2BX1 U189 ( .AN(n79), .B(n94), .Y(n93) );
  INVX1 U190 ( .A(n92), .Y(n94) );
  NAND2X1 U191 ( .A(n59), .B(n60), .Y(n65) );
  INVX1 U192 ( .A(n108), .Y(n103) );
  INVX1 U193 ( .A(n135), .Y(n130) );
  XOR2X1 U194 ( .A(n117), .B(n119), .Y(SUM[20]) );
  NOR2BX1 U195 ( .AN(n104), .B(n120), .Y(n119) );
  INVX1 U196 ( .A(n118), .Y(n120) );
  XOR2X1 U197 ( .A(n146), .B(n148), .Y(SUM[16]) );
  NOR2BX1 U198 ( .AN(n131), .B(n149), .Y(n148) );
  INVX1 U199 ( .A(n147), .Y(n149) );
  NOR2BX1 U200 ( .AN(n48), .B(n11), .Y(n47) );
  INVX1 U201 ( .A(n51), .Y(n49) );
  XOR2X1 U202 ( .A(n63), .B(n136), .Y(SUM[1]) );
  XOR2X1 U203 ( .A(n51), .B(n61), .Y(SUM[2]) );
  AOI21X1 U204 ( .A0(n126), .A1(n127), .B0(n21), .Y(n125) );
  AOI21X1 U205 ( .A0(n99), .A1(n100), .B0(n22), .Y(n98) );
  NAND2BX1 U206 ( .AN(n101), .B(n102), .Y(n99) );
  OAI2BB1X1 U207 ( .A0N(n62), .A1N(n63), .B0(n64), .Y(n51) );
  INVX1 U208 ( .A(n138), .Y(n63) );
  INVX1 U209 ( .A(n83), .Y(n78) );
  AOI21X1 U210 ( .A0(n74), .A1(n75), .B0(n23), .Y(n73) );
  NAND2BX1 U211 ( .AN(n76), .B(n77), .Y(n74) );
  OAI21XL U212 ( .A0(n78), .A1(n79), .B0(n80), .Y(n77) );
  INVX1 U213 ( .A(n82), .Y(n76) );
  NAND2X1 U214 ( .A(B[1]), .B(A[1]), .Y(n64) );
  OR2X2 U215 ( .A(A[6]), .B(B[6]), .Y(n33) );
  NAND2X1 U216 ( .A(B[4]), .B(A[4]), .Y(n42) );
  NAND2X1 U217 ( .A(B[12]), .B(A[12]), .Y(n160) );
  NAND2X1 U218 ( .A(B[6]), .B(A[6]), .Y(n35) );
  NOR2X1 U219 ( .A(A[23]), .B(B[23]), .Y(n22) );
  NAND2X1 U220 ( .A(B[21]), .B(A[21]), .Y(n105) );
  XOR3X2 U221 ( .A(B[31]), .B(A[31]), .C(n52), .Y(SUM[31]) );
  NAND2X1 U222 ( .A(n53), .B(n54), .Y(n52) );
  OR2X2 U223 ( .A(A[22]), .B(B[22]), .Y(n107) );
  NOR2X1 U224 ( .A(A[27]), .B(B[27]), .Y(n23) );
  NAND2X1 U225 ( .A(B[24]), .B(A[24]), .Y(n79) );
  NAND2X1 U226 ( .A(B[25]), .B(A[25]), .Y(n80) );
  OR2X2 U227 ( .A(A[25]), .B(B[25]), .Y(n83) );
  OR2X2 U228 ( .A(A[26]), .B(B[26]), .Y(n82) );
  NAND2X1 U229 ( .A(B[23]), .B(A[23]), .Y(n106) );
  OR2X2 U230 ( .A(A[24]), .B(B[24]), .Y(n92) );
  NAND2X1 U231 ( .A(B[26]), .B(A[26]), .Y(n75) );
  NAND2X1 U232 ( .A(B[29]), .B(A[29]), .Y(n59) );
  NAND2X1 U233 ( .A(B[28]), .B(A[28]), .Y(n69) );
  OR2X2 U234 ( .A(A[28]), .B(B[28]), .Y(n67) );
  NAND2X1 U235 ( .A(B[27]), .B(A[27]), .Y(n81) );
  OR2X2 U236 ( .A(A[29]), .B(B[29]), .Y(n60) );
  NAND2X1 U237 ( .A(B[30]), .B(A[30]), .Y(n53) );
  OR2X2 U238 ( .A(A[30]), .B(B[30]), .Y(n56) );
endmodule


module hash_core_DW01_add_38 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n339, n340, n341, n342, n1, n2, n3, n4, n5, n6, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n80, n81, n82, n83,
         n84, n85, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338;

  NAND3X4 U2 ( .A(n64), .B(n75), .C(n28), .Y(n93) );
  NAND3X4 U3 ( .A(n263), .B(n262), .C(n272), .Y(n240) );
  NAND2X1 U4 ( .A(B[6]), .B(A[6]), .Y(n122) );
  NAND2X2 U5 ( .A(n107), .B(n65), .Y(n64) );
  AOI21X2 U6 ( .A0(n160), .A1(n161), .B0(n162), .Y(n159) );
  NOR2BX4 U7 ( .AN(n168), .B(n32), .Y(n160) );
  NOR2X2 U8 ( .A(n300), .B(n301), .Y(n299) );
  INVX8 U9 ( .A(n270), .Y(n119) );
  AND2X4 U10 ( .A(n304), .B(n9), .Y(n12) );
  BUFX16 U11 ( .A(n340), .Y(SUM[10]) );
  NOR2X4 U12 ( .A(B[17]), .B(A[17]), .Y(n1) );
  NAND2X4 U13 ( .A(n87), .B(n138), .Y(n90) );
  INVX3 U14 ( .A(n137), .Y(n87) );
  CLKINVX4 U15 ( .A(n274), .Y(n108) );
  BUFX12 U16 ( .A(n339), .Y(SUM[26]) );
  CLKINVX8 U17 ( .A(n181), .Y(n252) );
  NAND2X4 U18 ( .A(n131), .B(n3), .Y(n4) );
  NAND2X4 U19 ( .A(n2), .B(n132), .Y(n5) );
  NAND2X4 U20 ( .A(n4), .B(n5), .Y(SUM[5]) );
  CLKINVX2 U21 ( .A(n131), .Y(n2) );
  INVX4 U22 ( .A(n132), .Y(n3) );
  NAND2X2 U23 ( .A(n128), .B(n31), .Y(n131) );
  NAND2X2 U24 ( .A(n239), .B(n51), .Y(n238) );
  INVX3 U25 ( .A(n24), .Y(n25) );
  INVX2 U26 ( .A(n112), .Y(n325) );
  BUFX4 U27 ( .A(n311), .Y(n6) );
  NAND2X4 U28 ( .A(n242), .B(n80), .Y(n254) );
  NAND2X2 U29 ( .A(n163), .B(n168), .Y(n172) );
  NOR2X4 U30 ( .A(n285), .B(n286), .Y(n279) );
  NAND3X4 U31 ( .A(n127), .B(n128), .C(n129), .Y(n96) );
  BUFX12 U32 ( .A(n342), .Y(SUM[2]) );
  NAND2X1 U33 ( .A(n144), .B(n145), .Y(n143) );
  INVX8 U34 ( .A(n271), .Y(n332) );
  XOR2X4 U35 ( .A(n155), .B(n156), .Y(SUM[28]) );
  XOR2X4 U36 ( .A(n149), .B(n153), .Y(SUM[29]) );
  NAND3BX4 U37 ( .AN(n45), .B(n174), .C(n166), .Y(n72) );
  BUFX2 U38 ( .A(n126), .Y(n31) );
  NAND2X2 U39 ( .A(B[12]), .B(A[12]), .Y(n287) );
  NOR2BX4 U40 ( .AN(n167), .B(n32), .Y(n173) );
  NAND2X2 U41 ( .A(B[26]), .B(A[26]), .Y(n167) );
  NOR2BX4 U42 ( .AN(n152), .B(n55), .Y(n229) );
  DLY1X1 U43 ( .A(B[11]), .Y(n70) );
  XOR2X4 U44 ( .A(n144), .B(n146), .Y(SUM[30]) );
  DLY1X1 U45 ( .A(B[7]), .Y(n10) );
  NOR2BX2 U46 ( .AN(n193), .B(n218), .Y(n217) );
  XNOR3X4 U47 ( .A(B[31]), .B(n40), .C(n41), .Y(SUM[31]) );
  NAND2X2 U48 ( .A(n142), .B(n143), .Y(n41) );
  BUFX4 U49 ( .A(n241), .Y(n80) );
  NAND2X4 U50 ( .A(n84), .B(n85), .Y(SUM[4]) );
  NOR2BX4 U51 ( .AN(n140), .B(n100), .Y(n150) );
  XOR2X4 U52 ( .A(n15), .B(n229), .Y(SUM[1]) );
  BUFX8 U53 ( .A(n122), .Y(n9) );
  NOR2BX2 U54 ( .AN(n130), .B(n24), .Y(n136) );
  INVX8 U55 ( .A(n127), .Y(n24) );
  OAI2BB1X4 U56 ( .A0N(n212), .A1N(n56), .B0(n213), .Y(n210) );
  CLKINVX4 U57 ( .A(n252), .Y(n56) );
  INVX4 U58 ( .A(n54), .Y(n158) );
  INVX1 U59 ( .A(n208), .Y(n212) );
  NOR2X1 U60 ( .A(n325), .B(n326), .Y(n323) );
  CLKINVX2 U61 ( .A(n32), .Y(n170) );
  INVX1 U62 ( .A(B[18]), .Y(n61) );
  NAND3BX2 U63 ( .AN(n23), .B(n197), .C(n191), .Y(n188) );
  NOR2X1 U64 ( .A(A[21]), .B(B[21]), .Y(n23) );
  INVX1 U65 ( .A(n67), .Y(n66) );
  INVX1 U66 ( .A(n228), .Y(n67) );
  OAI2BB1X2 U67 ( .A0N(B[2]), .A1N(A[2]), .B0(n152), .Y(n335) );
  NOR2X2 U68 ( .A(n55), .B(n337), .Y(n334) );
  NOR2X2 U69 ( .A(n78), .B(n80), .Y(n247) );
  INVX1 U70 ( .A(n234), .Y(n249) );
  NOR2X1 U71 ( .A(n164), .B(n171), .Y(n169) );
  NOR2BX1 U72 ( .AN(n166), .B(n164), .Y(n179) );
  NOR2X2 U73 ( .A(n208), .B(n209), .Y(n204) );
  NOR2BX2 U74 ( .AN(n44), .B(n326), .Y(n328) );
  INVX1 U75 ( .A(n135), .Y(n82) );
  INVX2 U76 ( .A(n123), .Y(n120) );
  INVX4 U77 ( .A(n176), .Y(n171) );
  INVX1 U78 ( .A(n211), .Y(n36) );
  NOR2BX1 U79 ( .AN(n192), .B(n209), .Y(n211) );
  XOR2X2 U80 ( .A(n141), .B(n150), .Y(n342) );
  AOI21X1 U81 ( .A0(n234), .A1(n223), .B0(n235), .Y(n233) );
  CLKINVX3 U82 ( .A(n30), .Y(SUM[0]) );
  NAND2BX1 U83 ( .AN(n15), .B(n338), .Y(n30) );
  NAND2X1 U84 ( .A(n135), .B(n83), .Y(n84) );
  NAND2X1 U85 ( .A(n82), .B(n136), .Y(n85) );
  INVX1 U86 ( .A(n136), .Y(n83) );
  INVX1 U87 ( .A(n138), .Y(n88) );
  INVX1 U88 ( .A(n167), .Y(n59) );
  NOR2BX1 U89 ( .AN(n148), .B(n106), .Y(n153) );
  AND2X2 U90 ( .A(n142), .B(n145), .Y(n146) );
  INVX1 U91 ( .A(A[31]), .Y(n40) );
  INVX1 U92 ( .A(n206), .Y(n213) );
  BUFX1 U93 ( .A(n111), .Y(n19) );
  NOR2X1 U94 ( .A(A[28]), .B(B[28]), .Y(n105) );
  NOR2X2 U95 ( .A(n130), .B(n77), .Y(n125) );
  NOR2X2 U96 ( .A(B[5]), .B(A[5]), .Y(n77) );
  AND2X1 U97 ( .A(n227), .B(n237), .Y(n11) );
  AND3X4 U98 ( .A(n33), .B(n197), .C(n35), .Y(n13) );
  AND2X2 U99 ( .A(n176), .B(n175), .Y(n14) );
  AND2X2 U100 ( .A(B[0]), .B(A[0]), .Y(n15) );
  INVX1 U101 ( .A(n46), .Y(n326) );
  AND2X4 U102 ( .A(n228), .B(n237), .Y(n16) );
  AND2X2 U103 ( .A(n135), .B(n116), .Y(n17) );
  NAND2X2 U104 ( .A(B[3]), .B(A[3]), .Y(n18) );
  INVX1 U105 ( .A(n35), .Y(n201) );
  CLKINVX3 U106 ( .A(n196), .Y(n215) );
  INVX1 U107 ( .A(n277), .Y(n286) );
  AOI21X4 U108 ( .A0(n308), .A1(n257), .B0(n309), .Y(n306) );
  INVX1 U109 ( .A(n287), .Y(n309) );
  NAND2X4 U110 ( .A(n20), .B(n298), .Y(n257) );
  INVX4 U111 ( .A(n319), .Y(n20) );
  NAND2BX4 U112 ( .AN(B[6]), .B(n21), .Y(n76) );
  INVX1 U113 ( .A(A[6]), .Y(n21) );
  NOR2X4 U114 ( .A(n261), .B(n68), .Y(n263) );
  NAND2BX4 U115 ( .AN(B[6]), .B(n21), .Y(n318) );
  OAI2BB1X4 U116 ( .A0N(A[16]), .A1N(B[16]), .B0(n251), .Y(n250) );
  NAND2X4 U117 ( .A(n22), .B(n48), .Y(n265) );
  INVX4 U118 ( .A(B[14]), .Y(n22) );
  INVX1 U119 ( .A(A[14]), .Y(n48) );
  AOI2BB1X4 U120 ( .A0N(B[5]), .A1N(A[5]), .B0(n130), .Y(n331) );
  AND3X4 U121 ( .A(n185), .B(n13), .C(n215), .Y(n182) );
  OAI21X2 U122 ( .A0(n1), .A1(n226), .B0(n227), .Y(n234) );
  BUFX20 U123 ( .A(n269), .Y(n107) );
  BUFX2 U124 ( .A(n261), .Y(n73) );
  BUFX2 U125 ( .A(n158), .Y(n92) );
  NAND2X4 U126 ( .A(n197), .B(n189), .Y(n214) );
  AND2X4 U127 ( .A(n318), .B(n128), .Y(n101) );
  INVX2 U128 ( .A(n318), .Y(n121) );
  INVXL U129 ( .A(n302), .Y(n301) );
  NOR2BX2 U130 ( .AN(n9), .B(n121), .Y(n124) );
  BUFX2 U131 ( .A(n259), .Y(n26) );
  NOR2BX4 U132 ( .AN(n76), .B(n77), .Y(n333) );
  NOR2BX4 U133 ( .AN(n27), .B(n238), .Y(n231) );
  AND2X2 U134 ( .A(n242), .B(n80), .Y(n27) );
  NOR2BX4 U135 ( .AN(n298), .B(n43), .Y(n296) );
  NOR2X4 U136 ( .A(A[3]), .B(B[3]), .Y(n103) );
  XNOR2X4 U137 ( .A(n310), .B(n6), .Y(SUM[12]) );
  CLKBUFX2 U138 ( .A(n109), .Y(n28) );
  XNOR2X4 U139 ( .A(n305), .B(n29), .Y(SUM[13]) );
  NAND2X1 U140 ( .A(n108), .B(n276), .Y(n29) );
  NAND3BX4 U141 ( .AN(n125), .B(n96), .C(n31), .Y(n123) );
  INVX4 U142 ( .A(n189), .Y(n219) );
  NOR2X4 U143 ( .A(A[26]), .B(B[26]), .Y(n32) );
  OR2X4 U144 ( .A(A[21]), .B(B[21]), .Y(n33) );
  OR2X4 U145 ( .A(A[21]), .B(B[21]), .Y(n34) );
  OR2X4 U146 ( .A(A[22]), .B(B[22]), .Y(n35) );
  NAND3X1 U147 ( .A(n190), .B(n34), .C(n191), .Y(n186) );
  XNOR2X4 U148 ( .A(n210), .B(n36), .Y(SUM[21]) );
  NOR2X2 U149 ( .A(B[12]), .B(A[12]), .Y(n37) );
  CLKBUFX2 U150 ( .A(n103), .Y(n38) );
  NAND3BX4 U151 ( .AN(n45), .B(n174), .C(n166), .Y(n39) );
  NOR2X2 U152 ( .A(n165), .B(n164), .Y(n45) );
  BUFX3 U153 ( .A(n276), .Y(n49) );
  BUFX12 U154 ( .A(n115), .Y(n42) );
  OAI2BB1X2 U155 ( .A0N(A[11]), .A1N(B[11]), .B0(n297), .Y(n43) );
  NAND3X4 U156 ( .A(n313), .B(n314), .C(n289), .Y(n307) );
  NAND2X1 U157 ( .A(n226), .B(n228), .Y(n253) );
  BUFX8 U158 ( .A(n297), .Y(n44) );
  OAI2BB1X4 U159 ( .A0N(n288), .A1N(n257), .B0(n312), .Y(n310) );
  AND2X1 U160 ( .A(n111), .B(n109), .Y(n57) );
  NAND2BX4 U161 ( .AN(n119), .B(n107), .Y(n284) );
  NAND2X4 U162 ( .A(n177), .B(n14), .Y(n174) );
  NOR2BX2 U163 ( .AN(n194), .B(n200), .Y(n199) );
  NOR2BX2 U164 ( .AN(n277), .B(n26), .Y(n292) );
  AND2X2 U165 ( .A(n111), .B(n47), .Y(n53) );
  INVX4 U166 ( .A(n325), .Y(n47) );
  OR2X4 U167 ( .A(B[10]), .B(A[10]), .Y(n46) );
  NOR2X2 U168 ( .A(n242), .B(n78), .Y(n248) );
  NAND3X2 U169 ( .A(n169), .B(n170), .C(n168), .Y(n157) );
  AOI21X4 U170 ( .A0(n299), .A1(n42), .B0(n68), .Y(n294) );
  NAND2X4 U171 ( .A(n17), .B(n332), .Y(n110) );
  INVX8 U172 ( .A(n16), .Y(n78) );
  NAND3X4 U173 ( .A(n50), .B(n186), .C(n187), .Y(n184) );
  AND2X4 U174 ( .A(n194), .B(n195), .Y(n50) );
  NAND3X4 U175 ( .A(n263), .B(n262), .C(n272), .Y(n51) );
  NOR2X4 U176 ( .A(n260), .B(n259), .Y(n272) );
  AOI21X2 U177 ( .A0(n284), .A1(n42), .B0(n37), .Y(n281) );
  NAND2X1 U178 ( .A(n109), .B(n116), .Y(n113) );
  CLKINVX2 U179 ( .A(n258), .Y(n52) );
  XOR2X4 U180 ( .A(n93), .B(n53), .Y(SUM[9]) );
  NAND3X2 U181 ( .A(n64), .B(n75), .C(n57), .Y(n324) );
  NOR2X4 U182 ( .A(n71), .B(n283), .Y(n282) );
  NAND2X4 U183 ( .A(n267), .B(n268), .Y(n262) );
  OAI2BB1X4 U184 ( .A0N(n182), .A1N(n56), .B0(n183), .Y(n54) );
  NOR2X4 U185 ( .A(B[13]), .B(A[13]), .Y(n274) );
  INVX4 U186 ( .A(n314), .Y(n71) );
  NOR2X4 U187 ( .A(A[1]), .B(B[1]), .Y(n55) );
  NAND4BX2 U188 ( .AN(n1), .B(n228), .C(n223), .D(n62), .Y(n196) );
  NAND2X4 U189 ( .A(n114), .B(n42), .Y(n313) );
  XOR2X2 U190 ( .A(n123), .B(n124), .Y(n341) );
  XOR2X4 U191 ( .A(n39), .B(n173), .Y(n339) );
  OAI21X4 U192 ( .A0(A[11]), .A1(B[11]), .B0(n46), .Y(n315) );
  NAND4BX2 U193 ( .AN(n283), .B(n257), .C(n289), .D(n52), .Y(n278) );
  NAND2XL U194 ( .A(n289), .B(n287), .Y(n311) );
  NOR2X4 U195 ( .A(n258), .B(n259), .Y(n256) );
  NAND3X4 U196 ( .A(n330), .B(n110), .C(n28), .Y(n329) );
  AOI21X4 U197 ( .A0(n72), .A1(n170), .B0(n59), .Y(n58) );
  AOI2BB1X4 U198 ( .A0N(n60), .A1N(n61), .B0(n225), .Y(n220) );
  CLKINVX20 U199 ( .A(A[18]), .Y(n60) );
  NAND2X4 U200 ( .A(n107), .B(n65), .Y(n330) );
  NAND2X2 U201 ( .A(n107), .B(n74), .Y(n268) );
  NOR2X4 U202 ( .A(n261), .B(n260), .Y(n255) );
  OR2X4 U203 ( .A(B[19]), .B(A[19]), .Y(n62) );
  INVX4 U204 ( .A(n219), .Y(n63) );
  NAND4X4 U205 ( .A(n303), .B(n304), .C(n9), .D(n302), .Y(n269) );
  AND2X4 U206 ( .A(n270), .B(n116), .Y(n65) );
  NAND2BX4 U207 ( .AN(n119), .B(n107), .Y(n114) );
  NOR2X4 U208 ( .A(n258), .B(n37), .Y(n308) );
  NAND2X4 U209 ( .A(n181), .B(n66), .Y(n251) );
  NAND2X4 U210 ( .A(n108), .B(n265), .Y(n283) );
  NAND2BX4 U211 ( .AN(n315), .B(n102), .Y(n68) );
  INVX8 U212 ( .A(n264), .Y(n314) );
  OAI2BB1X4 U213 ( .A0N(n323), .A1N(n324), .B0(n44), .Y(n321) );
  NAND2X4 U214 ( .A(A[9]), .B(B[9]), .Y(n111) );
  INVX2 U215 ( .A(n130), .Y(n133) );
  NOR2X4 U216 ( .A(n260), .B(n259), .Y(n69) );
  NAND2X4 U217 ( .A(B[1]), .B(A[1]), .Y(n152) );
  INVX8 U218 ( .A(n266), .Y(n260) );
  AND2X4 U219 ( .A(n112), .B(n116), .Y(n102) );
  OAI21X2 U220 ( .A0(A[7]), .A1(B[7]), .B0(n127), .Y(n317) );
  INVX4 U221 ( .A(n141), .Y(n139) );
  NAND2X4 U222 ( .A(B[25]), .B(A[25]), .Y(n166) );
  NAND2X1 U223 ( .A(B[2]), .B(A[2]), .Y(n140) );
  XOR2X2 U224 ( .A(n177), .B(n180), .Y(SUM[24]) );
  NAND2X4 U225 ( .A(A[13]), .B(B[13]), .Y(n276) );
  NAND2X4 U226 ( .A(A[7]), .B(B[7]), .Y(n302) );
  NAND2X2 U227 ( .A(B[17]), .B(A[17]), .Y(n227) );
  OAI21X4 U228 ( .A0(n1), .A1(n226), .B0(n227), .Y(n225) );
  NAND3BX4 U229 ( .AN(n254), .B(n239), .C(n240), .Y(n181) );
  NOR2X4 U230 ( .A(A[2]), .B(B[2]), .Y(n100) );
  BUFX8 U231 ( .A(n341), .Y(SUM[6]) );
  NOR2BX2 U232 ( .AN(n165), .B(n171), .Y(n180) );
  OR2X4 U233 ( .A(A[7]), .B(B[7]), .Y(n104) );
  INVX4 U234 ( .A(n34), .Y(n209) );
  AOI21X4 U235 ( .A0(n206), .A1(n33), .B0(n207), .Y(n205) );
  NAND2BX2 U236 ( .AN(n271), .B(n129), .Y(n267) );
  NAND3X4 U237 ( .A(n104), .B(n333), .C(n25), .Y(n271) );
  CLKINVX2 U238 ( .A(n119), .Y(n74) );
  OAI21X4 U239 ( .A0(n158), .A1(n171), .B0(n165), .Y(n178) );
  INVX4 U240 ( .A(n149), .Y(n147) );
  OR2X2 U241 ( .A(n51), .B(n78), .Y(n246) );
  NAND3X4 U242 ( .A(n116), .B(n332), .C(n135), .Y(n75) );
  NAND2X4 U243 ( .A(n18), .B(n134), .Y(n135) );
  OAI2BB1X4 U244 ( .A0N(B[11]), .A1N(A[11]), .B0(n297), .Y(n319) );
  NAND2X4 U245 ( .A(A[5]), .B(B[5]), .Y(n126) );
  NAND3X4 U246 ( .A(n320), .B(n112), .C(n316), .Y(n298) );
  AOI21X4 U247 ( .A0(n12), .A1(n303), .B0(n119), .Y(n300) );
  NOR2X4 U248 ( .A(n103), .B(n100), .Y(n336) );
  NOR2BX4 U249 ( .AN(n18), .B(n38), .Y(n138) );
  OAI211X1 U250 ( .A0(n164), .A1(n165), .B0(n166), .C0(n167), .Y(n161) );
  INVX8 U251 ( .A(n175), .Y(n164) );
  OAI2BB1X2 U252 ( .A0N(n215), .A1N(n181), .B0(n219), .Y(n216) );
  NAND3BX4 U253 ( .AN(n244), .B(n246), .C(n245), .Y(n243) );
  NAND2X2 U254 ( .A(n313), .B(n314), .Y(n312) );
  AOI21X2 U255 ( .A0(n276), .A1(n287), .B0(n283), .Y(n285) );
  NAND2X4 U256 ( .A(B[16]), .B(A[16]), .Y(n226) );
  NAND2X2 U257 ( .A(B[14]), .B(A[14]), .Y(n277) );
  NAND3BX4 U258 ( .AN(n317), .B(n101), .C(n135), .Y(n115) );
  AND2X2 U259 ( .A(n129), .B(n127), .Y(n81) );
  NOR2X4 U260 ( .A(n81), .B(n133), .Y(n132) );
  NAND2X4 U261 ( .A(n18), .B(n134), .Y(n129) );
  OAI21X2 U262 ( .A0(n139), .A1(n100), .B0(n140), .Y(n137) );
  NAND2X2 U263 ( .A(B[22]), .B(A[22]), .Y(n195) );
  NAND2X4 U264 ( .A(B[28]), .B(A[28]), .Y(n154) );
  NAND2X2 U265 ( .A(B[27]), .B(A[27]), .Y(n163) );
  NAND2X2 U266 ( .A(n88), .B(n137), .Y(n89) );
  NAND2X4 U267 ( .A(n89), .B(n90), .Y(SUM[3]) );
  INVX1 U268 ( .A(n105), .Y(n91) );
  OAI2BB1X4 U269 ( .A0N(n91), .A1N(n155), .B0(n154), .Y(n149) );
  NAND2X4 U270 ( .A(B[21]), .B(A[21]), .Y(n192) );
  OAI2BB1X4 U271 ( .A0N(n151), .A1N(n15), .B0(n152), .Y(n141) );
  NAND2X2 U272 ( .A(B[24]), .B(A[24]), .Y(n165) );
  NAND2XL U273 ( .A(A[0]), .B(B[0]), .Y(n337) );
  NAND2BX4 U274 ( .AN(n126), .B(n76), .Y(n304) );
  NAND2X2 U275 ( .A(n284), .B(n42), .Y(n95) );
  AND2X1 U276 ( .A(n236), .B(n223), .Y(n94) );
  NAND2XL U277 ( .A(B[15]), .B(A[15]), .Y(n241) );
  NAND2X2 U278 ( .A(B[20]), .B(A[20]), .Y(n193) );
  XNOR2X4 U279 ( .A(n95), .B(n113), .Y(SUM[8]) );
  XOR2X4 U280 ( .A(n97), .B(n98), .Y(SUM[15]) );
  NAND3X4 U281 ( .A(n278), .B(n279), .C(n280), .Y(n97) );
  AND2X1 U282 ( .A(n241), .B(n266), .Y(n98) );
  OAI21X4 U283 ( .A0(n106), .A1(n147), .B0(n148), .Y(n144) );
  OAI21X4 U284 ( .A0(n157), .A1(n92), .B0(n159), .Y(n155) );
  XOR2X4 U285 ( .A(n178), .B(n179), .Y(SUM[25]) );
  NOR2BX2 U286 ( .AN(n195), .B(n201), .Y(n203) );
  AND2X1 U287 ( .A(n222), .B(n224), .Y(n99) );
  OR2X4 U288 ( .A(A[18]), .B(B[18]), .Y(n223) );
  OAI21X4 U289 ( .A0(n120), .A1(n121), .B0(n9), .Y(n117) );
  OR2X4 U290 ( .A(A[16]), .B(B[16]), .Y(n228) );
  INVXL U291 ( .A(n197), .Y(n218) );
  NAND2X1 U292 ( .A(n192), .B(n193), .Y(n190) );
  INVX1 U293 ( .A(n192), .Y(n207) );
  INVXL U294 ( .A(n185), .Y(n200) );
  NOR2BX1 U295 ( .AN(n154), .B(n105), .Y(n156) );
  INVX1 U296 ( .A(n236), .Y(n235) );
  NAND3XL U297 ( .A(n237), .B(n223), .C(n228), .Y(n232) );
  INVX1 U298 ( .A(n163), .Y(n162) );
  NAND2BX4 U299 ( .AN(n315), .B(n102), .Y(n264) );
  OR2XL U300 ( .A(A[0]), .B(B[0]), .Y(n338) );
  NAND2X2 U301 ( .A(B[10]), .B(A[10]), .Y(n297) );
  NAND2XL U302 ( .A(B[18]), .B(A[18]), .Y(n236) );
  NAND2X1 U303 ( .A(B[19]), .B(A[19]), .Y(n222) );
  NAND2X1 U304 ( .A(B[30]), .B(A[30]), .Y(n142) );
  OR2X2 U305 ( .A(A[30]), .B(B[30]), .Y(n145) );
  NOR2X4 U306 ( .A(A[29]), .B(B[29]), .Y(n106) );
  INVX8 U307 ( .A(n288), .Y(n258) );
  OAI21X2 U308 ( .A0(n239), .A1(n78), .B0(n249), .Y(n244) );
  OAI2BB1X4 U309 ( .A0N(n202), .A1N(n35), .B0(n195), .Y(n198) );
  AOI21X2 U310 ( .A0(n10), .A1(A[7]), .B0(n119), .Y(n118) );
  NAND2X2 U311 ( .A(B[23]), .B(A[23]), .Y(n194) );
  INVX8 U312 ( .A(n265), .Y(n259) );
  AOI21X2 U313 ( .A0(n70), .A1(A[11]), .B0(n258), .Y(n322) );
  NAND2X1 U314 ( .A(A[12]), .B(B[12]), .Y(n275) );
  OAI2BB1X4 U315 ( .A0N(n56), .A1N(n182), .B0(n183), .Y(n177) );
  XOR2X4 U316 ( .A(n117), .B(n118), .Y(SUM[7]) );
  NAND2X4 U317 ( .A(B[29]), .B(A[29]), .Y(n148) );
  XOR2X4 U318 ( .A(n58), .B(n172), .Y(SUM[27]) );
  OR2X4 U319 ( .A(A[27]), .B(B[27]), .Y(n168) );
  OR2X4 U320 ( .A(A[25]), .B(B[25]), .Y(n175) );
  OR2X4 U321 ( .A(A[24]), .B(B[24]), .Y(n176) );
  NAND2X4 U322 ( .A(n184), .B(n185), .Y(n183) );
  NAND2BX4 U323 ( .AN(n188), .B(n63), .Y(n187) );
  XOR2X4 U324 ( .A(n198), .B(n199), .Y(SUM[23]) );
  OR2X4 U325 ( .A(A[23]), .B(B[23]), .Y(n185) );
  XOR2X4 U326 ( .A(n202), .B(n203), .Y(SUM[22]) );
  OR2X4 U327 ( .A(B[22]), .B(A[22]), .Y(n191) );
  OAI2BB1X4 U328 ( .A0N(n204), .A1N(n181), .B0(n205), .Y(n202) );
  NAND2X4 U329 ( .A(n214), .B(n193), .Y(n206) );
  NAND2X4 U330 ( .A(n215), .B(n197), .Y(n208) );
  XOR2X4 U331 ( .A(n216), .B(n217), .Y(SUM[20]) );
  OR2X4 U332 ( .A(A[20]), .B(B[20]), .Y(n197) );
  OAI21X4 U333 ( .A0(n220), .A1(n221), .B0(n222), .Y(n189) );
  NAND2X4 U334 ( .A(n223), .B(n224), .Y(n221) );
  XOR2X4 U335 ( .A(n230), .B(n99), .Y(SUM[19]) );
  OR2X4 U336 ( .A(A[19]), .B(B[19]), .Y(n224) );
  OAI21X4 U337 ( .A0(n231), .A1(n232), .B0(n233), .Y(n230) );
  XOR2X4 U338 ( .A(n243), .B(n94), .Y(SUM[18]) );
  NOR2X4 U339 ( .A(n247), .B(n248), .Y(n245) );
  XOR2X4 U340 ( .A(n250), .B(n11), .Y(SUM[17]) );
  OR2X4 U341 ( .A(B[17]), .B(A[17]), .Y(n237) );
  XOR2X4 U342 ( .A(n252), .B(n253), .Y(SUM[16]) );
  NAND3X4 U343 ( .A(n255), .B(n257), .C(n256), .Y(n239) );
  NAND2X4 U344 ( .A(n69), .B(n273), .Y(n242) );
  OAI211X2 U345 ( .A0(n274), .A1(n275), .B0(n276), .C0(n277), .Y(n273) );
  OR2X4 U346 ( .A(B[15]), .B(A[15]), .Y(n266) );
  NAND2X4 U347 ( .A(n281), .B(n282), .Y(n280) );
  XOR2X4 U348 ( .A(n291), .B(n292), .Y(SUM[14]) );
  OAI21X4 U349 ( .A0(n293), .A1(n73), .B0(n49), .Y(n291) );
  NAND2X4 U350 ( .A(n290), .B(n289), .Y(n261) );
  NOR2X4 U351 ( .A(n294), .B(n295), .Y(n293) );
  OAI21X4 U352 ( .A0(n296), .A1(n258), .B0(n287), .Y(n295) );
  OR2X4 U353 ( .A(B[13]), .B(A[13]), .Y(n290) );
  NAND2X4 U354 ( .A(n307), .B(n306), .Y(n305) );
  OR2X4 U355 ( .A(B[12]), .B(A[12]), .Y(n289) );
  NAND2X4 U356 ( .A(n111), .B(n109), .Y(n320) );
  XOR2X4 U357 ( .A(n321), .B(n322), .Y(SUM[11]) );
  OR2X4 U358 ( .A(B[11]), .B(A[11]), .Y(n288) );
  XOR2X4 U359 ( .A(n327), .B(n328), .Y(n340) );
  OR2X4 U360 ( .A(A[10]), .B(B[10]), .Y(n316) );
  OAI2BB1X4 U361 ( .A0N(n47), .A1N(n329), .B0(n19), .Y(n327) );
  NAND2X4 U362 ( .A(n331), .B(n318), .Y(n303) );
  NAND2X4 U363 ( .A(B[4]), .B(A[4]), .Y(n130) );
  OR2X4 U364 ( .A(A[7]), .B(B[7]), .Y(n270) );
  NAND2X4 U365 ( .A(A[8]), .B(B[8]), .Y(n109) );
  OR2X4 U366 ( .A(A[5]), .B(B[5]), .Y(n128) );
  OR2X4 U367 ( .A(A[4]), .B(B[4]), .Y(n127) );
  OAI21X4 U368 ( .A0(n334), .A1(n335), .B0(n336), .Y(n134) );
  OR2X4 U369 ( .A(A[1]), .B(B[1]), .Y(n151) );
  OR2X4 U370 ( .A(A[8]), .B(B[8]), .Y(n116) );
  OR2X4 U371 ( .A(B[9]), .B(A[9]), .Y(n112) );
endmodule


module hash_core_DW01_add_40 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n278, n279, n280, n1, n2, n3, n5, n6, n7, n9, n10, n11, n12, n13, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277;

  NAND2X4 U2 ( .A(n61), .B(n53), .Y(n268) );
  XOR2X2 U3 ( .A(n118), .B(n119), .Y(n279) );
  OAI2BB1X4 U4 ( .A0N(n124), .A1N(n12), .B0(n126), .Y(n120) );
  NAND2X1 U5 ( .A(B[0]), .B(A[0]), .Y(n273) );
  CLKINVX4 U6 ( .A(n50), .Y(n49) );
  INVX2 U7 ( .A(n125), .Y(n11) );
  NOR2X4 U8 ( .A(n48), .B(n201), .Y(n1) );
  NOR3X4 U9 ( .A(n2), .B(n204), .C(n203), .Y(n187) );
  INVX3 U10 ( .A(n1), .Y(n2) );
  NAND4BX2 U11 ( .AN(n260), .B(n261), .C(n262), .D(n263), .Y(n259) );
  BUFX3 U12 ( .A(n92), .Y(n3) );
  AOI21X2 U13 ( .A0(n161), .A1(n162), .B0(n163), .Y(n159) );
  NOR2X2 U14 ( .A(n29), .B(n167), .Y(n161) );
  BUFX8 U15 ( .A(n278), .Y(SUM[26]) );
  NAND2X1 U16 ( .A(n42), .B(n34), .Y(n41) );
  BUFX16 U17 ( .A(n43), .Y(n34) );
  CLKINVX4 U18 ( .A(n256), .Y(n42) );
  NOR2X1 U19 ( .A(n139), .B(n138), .Y(n124) );
  NAND2X2 U20 ( .A(n140), .B(n141), .Y(n138) );
  AOI2BB1X1 U21 ( .A0N(n139), .A1N(n11), .B0(n128), .Y(n158) );
  NAND2X4 U22 ( .A(n168), .B(n169), .Y(n139) );
  CLKINVX4 U23 ( .A(n37), .Y(n5) );
  INVX4 U24 ( .A(n5), .Y(n6) );
  XOR2X4 U25 ( .A(n71), .B(n72), .Y(SUM[3]) );
  NAND3X2 U26 ( .A(A[6]), .B(B[6]), .C(n53), .Y(n266) );
  OAI21X4 U27 ( .A0(n159), .A1(n32), .B0(n160), .Y(n128) );
  OAI21X4 U28 ( .A0(n175), .A1(n29), .B0(n164), .Y(n173) );
  BUFX4 U29 ( .A(n196), .Y(n7) );
  NAND2X1 U30 ( .A(B[14]), .B(A[14]), .Y(n196) );
  NOR2BX2 U31 ( .AN(n90), .B(n24), .Y(SUM[0]) );
  NAND2X2 U32 ( .A(B[0]), .B(A[0]), .Y(n90) );
  NAND4X4 U33 ( .A(n31), .B(n210), .C(n190), .D(n200), .Y(n201) );
  OR2X2 U34 ( .A(A[14]), .B(B[14]), .Y(n31) );
  NOR2X4 U35 ( .A(n198), .B(n199), .Y(n192) );
  INVX8 U36 ( .A(n217), .Y(n198) );
  XOR2X2 U37 ( .A(n147), .B(n149), .Y(SUM[22]) );
  NAND2X4 U38 ( .A(n120), .B(n121), .Y(n98) );
  BUFX3 U39 ( .A(n279), .Y(SUM[25]) );
  NAND2X4 U40 ( .A(n98), .B(n107), .Y(n118) );
  NAND2X1 U41 ( .A(B[4]), .B(A[4]), .Y(n63) );
  NOR2BXL U42 ( .AN(n160), .B(n32), .Y(n174) );
  NOR3BX2 U43 ( .AN(n18), .B(n205), .C(n206), .Y(n203) );
  NAND2X2 U44 ( .A(B[3]), .B(A[3]), .Y(n73) );
  INVX4 U45 ( .A(n34), .Y(n47) );
  CLKINVX3 U46 ( .A(n13), .Y(n183) );
  OAI2BB1X1 U47 ( .A0N(n181), .A1N(n125), .B0(n166), .Y(n13) );
  NAND2XL U48 ( .A(n63), .B(n68), .Y(n19) );
  NAND2X1 U49 ( .A(n165), .B(n166), .Y(n162) );
  OR2X2 U50 ( .A(A[8]), .B(B[8]), .Y(n269) );
  NAND2BX2 U51 ( .AN(n75), .B(n15), .Y(n207) );
  INVX1 U52 ( .A(n73), .Y(n205) );
  NOR2X2 U53 ( .A(n276), .B(n277), .Y(n274) );
  INVX1 U54 ( .A(n164), .Y(n163) );
  NOR2X1 U55 ( .A(n167), .B(n170), .Y(n168) );
  NOR2X2 U56 ( .A(A[18]), .B(B[18]), .Y(n29) );
  OAI21X1 U57 ( .A0(n82), .A1(n83), .B0(n84), .Y(n80) );
  CLKINVX3 U58 ( .A(n11), .Y(n12) );
  NAND3X2 U59 ( .A(n219), .B(n226), .C(n236), .Y(n234) );
  NAND2BX2 U60 ( .AN(n39), .B(n258), .Y(n263) );
  NAND2X1 U61 ( .A(n58), .B(n63), .Y(n62) );
  NOR2BX1 U62 ( .AN(n73), .B(n276), .Y(n72) );
  OAI21X2 U63 ( .A0(n114), .A1(n104), .B0(n103), .Y(n112) );
  XOR2X2 U64 ( .A(n145), .B(n146), .Y(SUM[23]) );
  AOI21X2 U65 ( .A0(n133), .A1(n147), .B0(n135), .Y(n146) );
  XNOR2X2 U66 ( .A(n150), .B(n152), .Y(SUM[21]) );
  INVX1 U67 ( .A(n110), .Y(n104) );
  NAND2X1 U68 ( .A(n190), .B(n195), .Y(n211) );
  AND3X2 U69 ( .A(n212), .B(n213), .C(n214), .Y(n27) );
  NOR2X1 U70 ( .A(n224), .B(n225), .Y(n212) );
  NOR2X1 U71 ( .A(n63), .B(n60), .Y(n65) );
  NOR2BX1 U72 ( .AN(n58), .B(n60), .Y(n70) );
  NOR2BX1 U73 ( .AN(n75), .B(n277), .Y(n86) );
  XNOR2X2 U74 ( .A(n90), .B(n171), .Y(SUM[1]) );
  NOR2BX2 U75 ( .AN(n89), .B(n172), .Y(n171) );
  INVX1 U76 ( .A(n87), .Y(n172) );
  OAI2BB1X2 U77 ( .A0N(n252), .A1N(n253), .B0(n244), .Y(n250) );
  NOR2X4 U78 ( .A(n34), .B(n62), .Y(n54) );
  BUFX3 U79 ( .A(n271), .Y(n15) );
  CLKINVX3 U80 ( .A(n151), .Y(n150) );
  AND2X4 U81 ( .A(n274), .B(n275), .Y(n9) );
  NAND2X1 U82 ( .A(B[16]), .B(A[16]), .Y(n166) );
  NAND2X1 U83 ( .A(B[1]), .B(A[1]), .Y(n89) );
  NAND2X1 U84 ( .A(B[5]), .B(A[5]), .Y(n58) );
  INVX4 U85 ( .A(n258), .Y(n38) );
  NOR2X1 U86 ( .A(n32), .B(n29), .Y(n169) );
  NAND2X2 U87 ( .A(B[2]), .B(A[2]), .Y(n75) );
  NAND2X1 U88 ( .A(n42), .B(n34), .Y(n255) );
  XOR2X2 U89 ( .A(n176), .B(n177), .Y(n280) );
  NAND2X2 U90 ( .A(n209), .B(n10), .Y(n185) );
  NOR3BX1 U91 ( .AN(n217), .B(n226), .C(n223), .Y(n224) );
  NAND2X2 U92 ( .A(n210), .B(n200), .Y(n223) );
  INVX8 U93 ( .A(n49), .Y(n10) );
  NOR2X2 U94 ( .A(n204), .B(n201), .Y(n209) );
  NAND4X2 U95 ( .A(B[5]), .B(A[5]), .C(n53), .D(n61), .Y(n265) );
  NAND2X1 U96 ( .A(n208), .B(n9), .Y(n18) );
  NAND3X2 U97 ( .A(n39), .B(n40), .C(n41), .Y(n35) );
  NAND2XL U98 ( .A(n200), .B(n197), .Y(n232) );
  OAI2BB1XL U99 ( .A0N(n230), .A1N(n197), .B0(n200), .Y(n218) );
  OAI2BB1X2 U100 ( .A0N(n153), .A1N(n125), .B0(n154), .Y(n151) );
  XOR2X2 U101 ( .A(n12), .B(n184), .Y(SUM[16]) );
  NOR3BX4 U102 ( .AN(n202), .B(n201), .C(n30), .Y(n188) );
  NAND2BX4 U103 ( .AN(n30), .B(n202), .Y(n226) );
  NAND3X2 U104 ( .A(B[4]), .B(A[4]), .C(n67), .Y(n267) );
  NAND3BX4 U105 ( .AN(n65), .B(n58), .C(n66), .Y(n64) );
  INVX1 U106 ( .A(n207), .Y(n206) );
  AOI21X2 U107 ( .A0(n3), .A1(n93), .B0(n94), .Y(n83) );
  INVX2 U108 ( .A(n76), .Y(n74) );
  OR2X4 U109 ( .A(A[1]), .B(B[1]), .Y(n87) );
  NAND3BX1 U110 ( .AN(n256), .B(n258), .C(n34), .Y(n261) );
  NOR2X2 U111 ( .A(n215), .B(n216), .Y(n214) );
  NOR2X1 U112 ( .A(n219), .B(n220), .Y(n215) );
  NAND2BX4 U113 ( .AN(n204), .B(n10), .Y(n219) );
  NAND3BX4 U114 ( .AN(n205), .B(n207), .C(n270), .Y(n43) );
  XNOR2X4 U115 ( .A(n34), .B(n19), .Y(SUM[4]) );
  INVX4 U116 ( .A(n176), .Y(n175) );
  NOR3X4 U117 ( .A(n187), .B(n188), .C(n189), .Y(n186) );
  XOR2X4 U118 ( .A(n112), .B(n113), .Y(SUM[27]) );
  NAND2X2 U119 ( .A(n25), .B(n34), .Y(n236) );
  NAND2X4 U120 ( .A(n25), .B(n34), .Y(n222) );
  AND2X4 U121 ( .A(n239), .B(n240), .Y(n25) );
  NOR2X2 U122 ( .A(A[3]), .B(B[3]), .Y(n276) );
  NAND3X2 U123 ( .A(n67), .B(n68), .C(n34), .Y(n66) );
  INVX4 U124 ( .A(n48), .Y(n240) );
  OAI21X2 U125 ( .A0(n47), .A1(n48), .B0(n49), .Y(n44) );
  NAND4BX4 U126 ( .AN(n23), .B(n68), .C(n61), .D(n53), .Y(n48) );
  XOR2X4 U127 ( .A(n44), .B(n45), .Y(SUM[8]) );
  XOR2X2 U128 ( .A(n76), .B(n86), .Y(SUM[2]) );
  BUFX4 U129 ( .A(n280), .Y(SUM[18]) );
  NOR2X4 U130 ( .A(A[2]), .B(B[2]), .Y(n277) );
  NOR2X2 U131 ( .A(A[19]), .B(B[19]), .Y(n32) );
  NOR2X1 U132 ( .A(A[5]), .B(B[5]), .Y(n23) );
  INVXL U133 ( .A(n28), .Y(n16) );
  OAI21X1 U134 ( .A0(n74), .A1(n277), .B0(n75), .Y(n71) );
  NOR2BX1 U135 ( .AN(n164), .B(n29), .Y(n177) );
  INVX1 U136 ( .A(n200), .Y(n199) );
  OR2X2 U137 ( .A(A[1]), .B(B[1]), .Y(n275) );
  NAND2X1 U138 ( .A(B[22]), .B(A[22]), .Y(n148) );
  NAND2X1 U139 ( .A(B[21]), .B(A[21]), .Y(n137) );
  OR2X2 U140 ( .A(A[16]), .B(B[16]), .Y(n181) );
  OAI21XL U141 ( .A0(n130), .A1(n131), .B0(n132), .Y(n129) );
  NOR2X2 U142 ( .A(A[21]), .B(B[21]), .Y(n28) );
  NAND2X4 U143 ( .A(n151), .B(n16), .Y(n17) );
  NAND2X4 U144 ( .A(n17), .B(n137), .Y(n147) );
  NAND2X1 U145 ( .A(B[11]), .B(A[11]), .Y(n246) );
  NAND2X1 U146 ( .A(B[15]), .B(A[15]), .Y(n195) );
  NOR2X4 U147 ( .A(A[11]), .B(B[11]), .Y(n30) );
  AOI21X4 U148 ( .A0(n234), .A1(n210), .B0(n235), .Y(n233) );
  INVXL U149 ( .A(n230), .Y(n235) );
  INVXL U150 ( .A(n136), .Y(n156) );
  NAND2X1 U151 ( .A(B[9]), .B(A[9]), .Y(n37) );
  NAND2X2 U152 ( .A(B[10]), .B(A[10]), .Y(n244) );
  NOR2BXL U153 ( .AN(n108), .B(n106), .Y(n119) );
  INVX3 U154 ( .A(n231), .Y(n229) );
  NAND3BXL U155 ( .AN(n33), .B(n110), .C(n111), .Y(n99) );
  NAND2X1 U156 ( .A(B[26]), .B(A[26]), .Y(n103) );
  NAND2XL U157 ( .A(B[25]), .B(A[25]), .Y(n108) );
  NAND3X4 U158 ( .A(n219), .B(n226), .C(n222), .Y(n231) );
  NAND2XL U159 ( .A(n132), .B(n143), .Y(n145) );
  XOR2X4 U160 ( .A(n27), .B(n211), .Y(SUM[15]) );
  XOR2X4 U161 ( .A(n64), .B(n20), .Y(SUM[6]) );
  AND2X1 U162 ( .A(n56), .B(n61), .Y(n20) );
  NAND3X1 U163 ( .A(n254), .B(n39), .C(n255), .Y(n253) );
  XOR2X4 U164 ( .A(n51), .B(n21), .Y(SUM[7]) );
  AND2X1 U165 ( .A(n52), .B(n53), .Y(n21) );
  NOR2BXL U166 ( .AN(n148), .B(n142), .Y(n149) );
  AND2X1 U167 ( .A(n244), .B(n257), .Y(n22) );
  NOR2BX1 U168 ( .AN(n109), .B(n101), .Y(n100) );
  INVXL U169 ( .A(n7), .Y(n225) );
  XOR2X2 U170 ( .A(n80), .B(n26), .Y(SUM[30]) );
  NOR2BXL U171 ( .AN(n166), .B(n170), .Y(n184) );
  INVX4 U172 ( .A(n180), .Y(n167) );
  OAI21X1 U173 ( .A0(n28), .A1(n136), .B0(n137), .Y(n134) );
  INVX2 U174 ( .A(n155), .Y(n144) );
  NOR2BX1 U175 ( .AN(n61), .B(n60), .Y(n59) );
  NAND2XL U176 ( .A(n136), .B(n155), .Y(n157) );
  NOR2XL U177 ( .A(n166), .B(n167), .Y(n178) );
  NAND3X2 U178 ( .A(n180), .B(n181), .C(n125), .Y(n179) );
  NOR2BXL U179 ( .AN(n109), .B(n33), .Y(n113) );
  XOR2XL U180 ( .A(n91), .B(n83), .Y(SUM[29]) );
  NAND2XL U181 ( .A(n80), .B(n81), .Y(n79) );
  OR2XL U182 ( .A(A[3]), .B(B[3]), .Y(n271) );
  NAND2XL U183 ( .A(B[23]), .B(A[23]), .Y(n132) );
  NAND2XL U184 ( .A(B[19]), .B(A[19]), .Y(n160) );
  OR2X4 U185 ( .A(A[22]), .B(B[22]), .Y(n133) );
  NOR2XL U186 ( .A(A[0]), .B(B[0]), .Y(n24) );
  OR2X4 U187 ( .A(A[25]), .B(B[25]), .Y(n111) );
  NAND2XL U188 ( .A(B[27]), .B(A[27]), .Y(n109) );
  INVX1 U189 ( .A(n223), .Y(n221) );
  AOI21X1 U190 ( .A0(n127), .A1(n128), .B0(n129), .Y(n126) );
  INVX1 U191 ( .A(n138), .Y(n127) );
  INVX1 U192 ( .A(n95), .Y(n94) );
  OAI21XL U193 ( .A0(n98), .A1(n99), .B0(n100), .Y(n92) );
  NOR2BX1 U194 ( .AN(n246), .B(n30), .Y(n251) );
  NOR2XL U195 ( .A(n38), .B(n247), .Y(n252) );
  INVX1 U196 ( .A(n85), .Y(n82) );
  INVX1 U197 ( .A(n143), .Y(n131) );
  INVX1 U198 ( .A(n133), .Y(n142) );
  INVX1 U199 ( .A(n181), .Y(n170) );
  XOR2X2 U200 ( .A(n115), .B(n116), .Y(n278) );
  NOR2BX1 U201 ( .AN(n103), .B(n104), .Y(n116) );
  XOR2X2 U202 ( .A(n231), .B(n237), .Y(SUM[12]) );
  NOR2BX1 U203 ( .AN(n230), .B(n238), .Y(n237) );
  INVX1 U204 ( .A(n210), .Y(n238) );
  NOR2BXL U205 ( .AN(n40), .B(n46), .Y(n45) );
  INVX1 U206 ( .A(n115), .Y(n114) );
  NOR2BX1 U207 ( .AN(n7), .B(n198), .Y(n228) );
  AOI21X1 U208 ( .A0(n133), .A1(n134), .B0(n135), .Y(n130) );
  NAND2X1 U209 ( .A(n180), .B(n165), .Y(n182) );
  XOR2X2 U210 ( .A(n157), .B(n158), .Y(SUM[20]) );
  XOR2X1 U211 ( .A(n120), .B(n122), .Y(SUM[24]) );
  NOR2BX1 U212 ( .AN(n107), .B(n123), .Y(n122) );
  INVX1 U213 ( .A(n121), .Y(n123) );
  NOR2BXL U214 ( .AN(n6), .B(n38), .Y(n36) );
  NOR2BX1 U215 ( .AN(n137), .B(n28), .Y(n152) );
  AND2X2 U216 ( .A(n78), .B(n81), .Y(n26) );
  NAND3BXL U217 ( .AN(n222), .B(n217), .C(n221), .Y(n213) );
  OAI2BB1X2 U218 ( .A0N(n87), .A1N(n88), .B0(n89), .Y(n76) );
  CLKINVX3 U219 ( .A(n90), .Y(n88) );
  NOR2X2 U220 ( .A(n139), .B(n144), .Y(n153) );
  AOI21X2 U221 ( .A0(n128), .A1(n155), .B0(n156), .Y(n154) );
  NOR2X1 U222 ( .A(n131), .B(n142), .Y(n141) );
  NOR2X1 U223 ( .A(n28), .B(n144), .Y(n140) );
  NOR2BX1 U224 ( .AN(n244), .B(n245), .Y(n243) );
  NAND2X1 U225 ( .A(n6), .B(n40), .Y(n242) );
  NOR2X2 U226 ( .A(n38), .B(n247), .Y(n241) );
  NOR2BX1 U227 ( .AN(n217), .B(n218), .Y(n216) );
  NAND2XL U228 ( .A(n221), .B(n217), .Y(n220) );
  NAND2X2 U229 ( .A(n240), .B(n269), .Y(n256) );
  NAND2BXL U230 ( .AN(n40), .B(n258), .Y(n262) );
  OAI2BB1X1 U231 ( .A0N(n57), .A1N(n58), .B0(n59), .Y(n55) );
  INVX1 U232 ( .A(n246), .Y(n245) );
  INVX1 U233 ( .A(n6), .Y(n260) );
  INVX1 U234 ( .A(n111), .Y(n106) );
  INVX1 U235 ( .A(n148), .Y(n135) );
  XOR2X1 U236 ( .A(n3), .B(n96), .Y(SUM[28]) );
  NOR2BX1 U237 ( .AN(n95), .B(n97), .Y(n96) );
  INVX1 U238 ( .A(n93), .Y(n97) );
  NAND2X1 U239 ( .A(n84), .B(n85), .Y(n91) );
  AOI21X1 U240 ( .A0(n102), .A1(n103), .B0(n33), .Y(n101) );
  NAND2BX1 U241 ( .AN(n104), .B(n105), .Y(n102) );
  OAI21XL U242 ( .A0(n106), .A1(n107), .B0(n108), .Y(n105) );
  NOR2X2 U243 ( .A(n267), .B(n268), .Y(n264) );
  NAND2X2 U244 ( .A(B[8]), .B(A[8]), .Y(n40) );
  NAND2XL U245 ( .A(B[13]), .B(A[13]), .Y(n197) );
  NAND2X1 U246 ( .A(B[18]), .B(A[18]), .Y(n164) );
  OR2X2 U247 ( .A(A[20]), .B(B[20]), .Y(n155) );
  NAND2XL U248 ( .A(B[7]), .B(A[7]), .Y(n52) );
  NAND2XL U249 ( .A(B[6]), .B(A[6]), .Y(n56) );
  NAND2XL U250 ( .A(B[12]), .B(A[12]), .Y(n230) );
  AOI21X2 U251 ( .A0(n192), .A1(n193), .B0(n194), .Y(n191) );
  OAI2BB1X1 U252 ( .A0N(B[12]), .A1N(A[12]), .B0(n197), .Y(n193) );
  NAND2X2 U253 ( .A(n195), .B(n7), .Y(n194) );
  OR2X2 U254 ( .A(A[23]), .B(B[23]), .Y(n143) );
  OAI2BB1X1 U255 ( .A0N(B[1]), .A1N(A[1]), .B0(n273), .Y(n272) );
  OAI2BB1X1 U256 ( .A0N(B[1]), .A1N(A[1]), .B0(n90), .Y(n208) );
  NAND2X1 U257 ( .A(B[20]), .B(A[20]), .Y(n136) );
  NAND2X1 U258 ( .A(B[24]), .B(A[24]), .Y(n107) );
  OR2X2 U259 ( .A(A[24]), .B(B[24]), .Y(n121) );
  OR2X2 U260 ( .A(A[26]), .B(B[26]), .Y(n110) );
  XOR3X2 U261 ( .A(B[31]), .B(A[31]), .C(n77), .Y(SUM[31]) );
  NAND2X1 U262 ( .A(n78), .B(n79), .Y(n77) );
  OR2X2 U263 ( .A(A[28]), .B(B[28]), .Y(n93) );
  NOR2X1 U264 ( .A(A[27]), .B(B[27]), .Y(n33) );
  NAND2X1 U265 ( .A(B[30]), .B(A[30]), .Y(n78) );
  NAND2X1 U266 ( .A(B[29]), .B(A[29]), .Y(n84) );
  OR2X2 U267 ( .A(A[30]), .B(B[30]), .Y(n81) );
  NAND2X1 U268 ( .A(B[28]), .B(A[28]), .Y(n95) );
  OR2X2 U269 ( .A(A[29]), .B(B[29]), .Y(n85) );
  OR2X2 U270 ( .A(A[17]), .B(B[17]), .Y(n180) );
  NAND2X1 U271 ( .A(B[17]), .B(A[17]), .Y(n165) );
  XOR2X4 U272 ( .A(n35), .B(n36), .Y(SUM[9]) );
  OAI21X4 U273 ( .A0(n54), .A1(n55), .B0(n56), .Y(n51) );
  XOR2X4 U274 ( .A(n69), .B(n70), .Y(SUM[5]) );
  CLKINVX3 U275 ( .A(n67), .Y(n60) );
  OAI21X4 U276 ( .A0(n47), .A1(n57), .B0(n63), .Y(n69) );
  CLKINVX3 U277 ( .A(n68), .Y(n57) );
  OAI21X4 U278 ( .A0(n117), .A1(n106), .B0(n108), .Y(n115) );
  CLKINVX3 U279 ( .A(n118), .Y(n117) );
  XOR2X4 U280 ( .A(n173), .B(n174), .Y(SUM[19]) );
  NAND3BX4 U281 ( .AN(n178), .B(n165), .C(n179), .Y(n176) );
  XOR2X4 U282 ( .A(n182), .B(n183), .Y(SUM[17]) );
  NAND2X4 U283 ( .A(n185), .B(n186), .Y(n125) );
  NOR2BX4 U284 ( .AN(n190), .B(n191), .Y(n189) );
  OR2X4 U285 ( .A(A[15]), .B(B[15]), .Y(n190) );
  XOR2X4 U286 ( .A(n227), .B(n228), .Y(SUM[14]) );
  OR2X4 U287 ( .A(A[14]), .B(B[14]), .Y(n217) );
  OAI21X4 U288 ( .A0(n229), .A1(n223), .B0(n218), .Y(n227) );
  XOR2X4 U289 ( .A(n232), .B(n233), .Y(SUM[13]) );
  OR2X4 U290 ( .A(A[13]), .B(B[13]), .Y(n200) );
  OR2X4 U291 ( .A(A[12]), .B(B[12]), .Y(n210) );
  CLKINVX3 U292 ( .A(n204), .Y(n239) );
  OAI2BB1X4 U293 ( .A0N(n241), .A1N(n242), .B0(n243), .Y(n202) );
  NAND2X4 U294 ( .A(n248), .B(n249), .Y(n204) );
  NOR2X4 U295 ( .A(n46), .B(n38), .Y(n249) );
  NOR2X4 U296 ( .A(n247), .B(n30), .Y(n248) );
  XOR2X4 U297 ( .A(n250), .B(n251), .Y(SUM[11]) );
  AND2X2 U298 ( .A(n6), .B(n40), .Y(n254) );
  CLKINVX3 U299 ( .A(n257), .Y(n247) );
  XOR2X4 U300 ( .A(n259), .B(n22), .Y(SUM[10]) );
  OR2X4 U301 ( .A(A[10]), .B(B[10]), .Y(n257) );
  NAND2BX4 U302 ( .AN(n46), .B(n50), .Y(n39) );
  NAND4BX4 U303 ( .AN(n264), .B(n265), .C(n52), .D(n266), .Y(n50) );
  OR2X4 U304 ( .A(A[5]), .B(B[5]), .Y(n67) );
  CLKINVX3 U305 ( .A(n269), .Y(n46) );
  NAND2X4 U306 ( .A(n9), .B(n272), .Y(n270) );
  OR2X4 U307 ( .A(A[9]), .B(B[9]), .Y(n258) );
  OR2X4 U308 ( .A(A[7]), .B(B[7]), .Y(n53) );
  OR2X4 U309 ( .A(A[6]), .B(B[6]), .Y(n61) );
  OR2X4 U310 ( .A(A[4]), .B(B[4]), .Y(n68) );
endmodule


module hash_core_DW01_add_43 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n290, n291, n292, n293, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n45, n47, n48, n49, n50, n52, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289;

  NAND2X1 U2 ( .A(B[14]), .B(A[14]), .Y(n223) );
  NAND2X4 U3 ( .A(n112), .B(n280), .Y(n1) );
  NAND2X1 U4 ( .A(n22), .B(n202), .Y(n230) );
  NOR2X4 U5 ( .A(B[9]), .B(A[9]), .Y(n26) );
  NAND2X4 U6 ( .A(n132), .B(n141), .Y(n151) );
  OAI21X4 U7 ( .A0(n216), .A1(n217), .B0(n218), .Y(n215) );
  NAND2X4 U8 ( .A(B[18]), .B(A[18]), .Y(n195) );
  NOR3X1 U9 ( .A(n225), .B(n236), .C(n246), .Y(n242) );
  NOR2X2 U10 ( .A(n29), .B(n289), .Y(n100) );
  NAND2X2 U11 ( .A(B[3]), .B(A[3]), .Y(n102) );
  NAND3X4 U12 ( .A(n271), .B(n3), .C(n16), .Y(n268) );
  NAND2X2 U13 ( .A(n78), .B(n77), .Y(n75) );
  NAND2X4 U14 ( .A(n223), .B(n224), .Y(n222) );
  NAND2X1 U15 ( .A(n110), .B(n19), .Y(n123) );
  OAI21X1 U16 ( .A0(n31), .A1(n94), .B0(n95), .Y(n93) );
  BUFX16 U17 ( .A(n73), .Y(n65) );
  NAND2X4 U18 ( .A(A[1]), .B(B[1]), .Y(n125) );
  BUFX16 U19 ( .A(n241), .Y(n45) );
  NOR2X4 U20 ( .A(n235), .B(n60), .Y(n256) );
  NOR2X4 U21 ( .A(n289), .B(n36), .Y(n288) );
  INVX8 U22 ( .A(n23), .Y(n76) );
  NAND2X4 U23 ( .A(n18), .B(n23), .Y(n101) );
  BUFX8 U24 ( .A(n102), .Y(n23) );
  BUFX8 U25 ( .A(n226), .Y(n2) );
  NOR3X4 U26 ( .A(n76), .B(n65), .C(n75), .Y(n69) );
  OR2X4 U27 ( .A(A[3]), .B(B[3]), .Y(n28) );
  OAI21X1 U28 ( .A0(n119), .A1(n120), .B0(n121), .Y(n117) );
  AOI21X4 U29 ( .A0(n127), .A1(n128), .B0(n129), .Y(n120) );
  OR2X4 U30 ( .A(B[3]), .B(A[3]), .Y(n280) );
  NAND2X2 U31 ( .A(B[17]), .B(A[17]), .Y(n196) );
  NAND2X2 U32 ( .A(n164), .B(n165), .Y(n161) );
  NAND3X2 U33 ( .A(n166), .B(n167), .C(n168), .Y(n164) );
  NOR2X2 U34 ( .A(n173), .B(n62), .Y(n172) );
  OAI21XL U35 ( .A0(n225), .A1(n2), .B0(n224), .Y(n50) );
  OAI21XL U36 ( .A0(n225), .A1(n2), .B0(n224), .Y(n245) );
  INVX1 U37 ( .A(n219), .Y(n236) );
  BUFX8 U38 ( .A(n293), .Y(SUM[1]) );
  NOR2BX2 U39 ( .AN(n2), .B(n246), .Y(n253) );
  INVX1 U40 ( .A(n152), .Y(n20) );
  NOR2BXL U41 ( .AN(n142), .B(n140), .Y(n152) );
  NAND2X1 U42 ( .A(n219), .B(n220), .Y(n217) );
  BUFX4 U43 ( .A(n26), .Y(n24) );
  NAND2X1 U44 ( .A(n169), .B(n170), .Y(n168) );
  AND2X2 U45 ( .A(n188), .B(n187), .Y(n194) );
  NOR2X1 U46 ( .A(n197), .B(n198), .Y(n192) );
  CLKINVX4 U47 ( .A(n74), .Y(n81) );
  INVX4 U48 ( .A(n267), .Y(n262) );
  OR2X2 U49 ( .A(A[25]), .B(B[25]), .Y(n145) );
  NAND2X2 U50 ( .A(B[20]), .B(A[20]), .Y(n170) );
  OR2X2 U51 ( .A(A[19]), .B(B[19]), .Y(n188) );
  OR2X2 U52 ( .A(n198), .B(n197), .Y(n37) );
  NOR2BX1 U53 ( .AN(n196), .B(n197), .Y(n208) );
  INVX1 U54 ( .A(n67), .Y(n282) );
  CLKBUFX8 U55 ( .A(n125), .Y(n22) );
  INVX1 U56 ( .A(A[7]), .Y(n32) );
  NAND2X1 U57 ( .A(B[24]), .B(A[24]), .Y(n141) );
  NAND2X1 U58 ( .A(n171), .B(n172), .Y(n157) );
  INVX1 U59 ( .A(n159), .Y(n49) );
  INVX1 U60 ( .A(n144), .Y(n138) );
  NOR2BX1 U61 ( .AN(n198), .B(n210), .Y(n209) );
  CLKINVX3 U62 ( .A(n40), .Y(n41) );
  INVX1 U63 ( .A(n179), .Y(n4) );
  BUFX3 U64 ( .A(n272), .Y(n16) );
  NOR2X1 U65 ( .A(n246), .B(n225), .Y(n249) );
  NAND2X1 U66 ( .A(n90), .B(n43), .Y(n98) );
  NAND2X1 U67 ( .A(n220), .B(n218), .Y(n239) );
  NAND2X1 U68 ( .A(n244), .B(n15), .Y(n243) );
  AOI21X4 U69 ( .A0(n65), .A1(n273), .B0(n282), .Y(n3) );
  AOI21X2 U70 ( .A0(n65), .A1(n273), .B0(n282), .Y(n270) );
  NOR2X2 U71 ( .A(n36), .B(n38), .Y(n276) );
  XOR2X2 U72 ( .A(n127), .B(n131), .Y(SUM[28]) );
  XNOR2X4 U73 ( .A(n178), .B(n4), .Y(SUM[22]) );
  NAND2XL U74 ( .A(B[25]), .B(A[25]), .Y(n142) );
  NOR2X4 U75 ( .A(n83), .B(n275), .Y(n274) );
  INVX4 U76 ( .A(n83), .Y(n72) );
  NAND2X1 U77 ( .A(n19), .B(n111), .Y(n109) );
  INVX8 U78 ( .A(n91), .Y(n82) );
  AND3X2 U79 ( .A(n188), .B(n9), .C(n187), .Y(n5) );
  INVX1 U80 ( .A(n166), .Y(n173) );
  OR2X2 U81 ( .A(A[21]), .B(B[21]), .Y(n166) );
  AND2X2 U82 ( .A(n196), .B(n37), .Y(n6) );
  AND2X2 U83 ( .A(n67), .B(n68), .Y(n7) );
  AND2X2 U84 ( .A(n191), .B(n190), .Y(n8) );
  AND2X2 U85 ( .A(n190), .B(n191), .Y(n9) );
  NOR2BX1 U86 ( .AN(n165), .B(n174), .Y(n179) );
  INVX1 U87 ( .A(n167), .Y(n174) );
  OR2X2 U88 ( .A(A[22]), .B(B[22]), .Y(n167) );
  INVX2 U89 ( .A(n65), .Y(n84) );
  OR2X4 U90 ( .A(B[9]), .B(A[9]), .Y(n68) );
  INVX1 U91 ( .A(n289), .Y(n11) );
  CLKINVX8 U92 ( .A(n36), .Y(n43) );
  CLKINVX3 U93 ( .A(n48), .Y(n153) );
  INVX4 U94 ( .A(n38), .Y(n90) );
  NOR2X4 U95 ( .A(n1), .B(n201), .Y(n10) );
  OAI21X4 U96 ( .A0(n158), .A1(n62), .B0(n170), .Y(n180) );
  NAND2BX1 U97 ( .AN(n31), .B(n11), .Y(n12) );
  CLKINVX3 U98 ( .A(n12), .Y(n92) );
  INVX4 U99 ( .A(n89), .Y(n31) );
  AND2X1 U100 ( .A(B[15]), .B(A[15]), .Y(n13) );
  CLKINVX3 U101 ( .A(n13), .Y(n218) );
  NOR2X4 U102 ( .A(n14), .B(n25), .Y(n104) );
  CLKINVX4 U103 ( .A(n78), .Y(n14) );
  NOR2BX4 U104 ( .AN(n22), .B(n201), .Y(n200) );
  NAND2X2 U105 ( .A(B[10]), .B(A[10]), .Y(n260) );
  NAND2X4 U106 ( .A(n21), .B(n8), .Y(n54) );
  INVX4 U107 ( .A(n77), .Y(n47) );
  INVX2 U108 ( .A(n201), .Y(n52) );
  BUFX3 U109 ( .A(n223), .Y(n15) );
  BUFX8 U110 ( .A(n86), .Y(n17) );
  OAI2BB1X4 U111 ( .A0N(n22), .A1N(n202), .B0(n10), .Y(n18) );
  NAND2X1 U112 ( .A(A[5]), .B(B[5]), .Y(n94) );
  NAND2X4 U113 ( .A(A[6]), .B(B[6]), .Y(n95) );
  OR2X2 U114 ( .A(B[2]), .B(A[2]), .Y(n19) );
  XOR2X2 U115 ( .A(n126), .B(n120), .Y(SUM[29]) );
  AND2X1 U116 ( .A(n195), .B(n187), .Y(n206) );
  XNOR2X4 U117 ( .A(n151), .B(n20), .Y(SUM[25]) );
  OAI2BB1X4 U118 ( .A0N(n178), .A1N(n167), .B0(n165), .Y(n176) );
  NAND2X4 U119 ( .A(n211), .B(n212), .Y(n21) );
  NOR2BX1 U120 ( .AN(n71), .B(n81), .Y(n80) );
  INVX4 U121 ( .A(n22), .Y(n113) );
  INVX1 U122 ( .A(n189), .Y(n40) );
  AND2X2 U123 ( .A(B[5]), .B(A[5]), .Y(n286) );
  NAND2BX4 U124 ( .AN(n110), .B(n28), .Y(n77) );
  NAND2X2 U125 ( .A(n23), .B(n77), .Y(n25) );
  AND2X1 U126 ( .A(n85), .B(n17), .Y(n35) );
  NAND2X4 U127 ( .A(n67), .B(n71), .Y(n258) );
  NAND2X4 U128 ( .A(n27), .B(n72), .Y(n254) );
  AND2X4 U129 ( .A(n263), .B(n264), .Y(n27) );
  INVX4 U130 ( .A(n43), .Y(n29) );
  OR2X4 U131 ( .A(B[1]), .B(A[1]), .Y(n111) );
  NOR2BXL U132 ( .AN(n261), .B(n60), .Y(n266) );
  NAND3X2 U133 ( .A(n271), .B(n270), .C(n16), .Y(n30) );
  NAND2X1 U134 ( .A(A[7]), .B(B[7]), .Y(n85) );
  BUFX12 U135 ( .A(n291), .Y(SUM[20]) );
  XOR2X4 U136 ( .A(n42), .B(n183), .Y(n291) );
  INVX4 U137 ( .A(n149), .Y(n148) );
  OAI2BB1X4 U138 ( .A0N(n145), .A1N(n151), .B0(n142), .Y(n149) );
  NAND4X4 U139 ( .A(n219), .B(n220), .C(n237), .D(n238), .Y(n231) );
  NAND2XL U140 ( .A(n219), .B(n15), .Y(n247) );
  AOI21X2 U141 ( .A0(n43), .A1(n92), .B0(n93), .Y(n87) );
  NAND2X4 U142 ( .A(n68), .B(n74), .Y(n275) );
  NAND2X2 U143 ( .A(B[12]), .B(A[12]), .Y(n226) );
  OAI2BB1X4 U144 ( .A0N(n190), .A1N(n21), .B0(n198), .Y(n207) );
  INVX8 U145 ( .A(n86), .Y(n278) );
  INVX4 U146 ( .A(n191), .Y(n197) );
  NAND2X4 U147 ( .A(A[4]), .B(B[4]), .Y(n289) );
  NAND2X2 U148 ( .A(B[11]), .B(A[11]), .Y(n261) );
  NAND2X4 U149 ( .A(n88), .B(n87), .Y(n34) );
  NAND2X2 U150 ( .A(B[9]), .B(A[9]), .Y(n67) );
  NAND2X2 U151 ( .A(n260), .B(n261), .Y(n259) );
  NOR2BX2 U152 ( .AN(n94), .B(n100), .Y(n99) );
  OR2X4 U153 ( .A(A[6]), .B(B[6]), .Y(n89) );
  NAND2BX4 U154 ( .AN(B[7]), .B(n32), .Y(n86) );
  XOR2X4 U155 ( .A(n82), .B(n33), .Y(SUM[4]) );
  NAND2XL U156 ( .A(n289), .B(n90), .Y(n33) );
  NOR2X4 U157 ( .A(n101), .B(n47), .Y(n97) );
  NOR2X4 U158 ( .A(n225), .B(n2), .Y(n221) );
  NAND2X2 U159 ( .A(n229), .B(n230), .Y(n228) );
  INVX4 U160 ( .A(n237), .Y(n246) );
  NAND2X4 U161 ( .A(A[2]), .B(B[2]), .Y(n110) );
  XOR2X4 U162 ( .A(n34), .B(n35), .Y(SUM[7]) );
  NOR2X4 U163 ( .A(B[5]), .B(A[5]), .Y(n36) );
  NAND2X2 U164 ( .A(B[13]), .B(A[13]), .Y(n224) );
  NAND2X4 U165 ( .A(n6), .B(n54), .Y(n205) );
  NOR2X4 U166 ( .A(B[4]), .B(A[4]), .Y(n38) );
  INVX8 U167 ( .A(n111), .Y(n201) );
  OAI2BB1X4 U168 ( .A0N(n205), .A1N(n187), .B0(n195), .Y(n203) );
  OAI21X4 U169 ( .A0(n254), .A1(n82), .B0(n255), .Y(n241) );
  INVX8 U170 ( .A(n182), .Y(n158) );
  NOR2X4 U171 ( .A(n231), .B(n232), .Y(n233) );
  OAI21X4 U172 ( .A0(n75), .A1(n76), .B0(n274), .Y(n271) );
  AOI21X4 U173 ( .A0(n52), .A1(n61), .B0(n113), .Y(n124) );
  NOR2X4 U174 ( .A(B[6]), .B(A[6]), .Y(n39) );
  XOR2X4 U175 ( .A(n41), .B(n209), .Y(SUM[16]) );
  INVX2 U176 ( .A(n158), .Y(n42) );
  NOR2X4 U177 ( .A(n278), .B(n39), .Y(n277) );
  NOR2X4 U178 ( .A(n232), .B(n231), .Y(n213) );
  NAND2X4 U179 ( .A(n5), .B(n189), .Y(n186) );
  XOR2X2 U180 ( .A(n180), .B(n181), .Y(n290) );
  NOR2X4 U181 ( .A(n221), .B(n222), .Y(n216) );
  OAI21X4 U182 ( .A0(n278), .A1(n95), .B0(n85), .Y(n283) );
  XOR2X4 U183 ( .A(n205), .B(n206), .Y(n292) );
  NOR2X4 U184 ( .A(n278), .B(n39), .Y(n287) );
  XNOR2X2 U185 ( .A(n202), .B(n200), .Y(n293) );
  AND2X4 U186 ( .A(n202), .B(n281), .Y(SUM[0]) );
  NAND2X4 U187 ( .A(B[0]), .B(A[0]), .Y(n202) );
  INVXL U188 ( .A(n28), .Y(n107) );
  AOI21X4 U189 ( .A0(n65), .A1(n27), .B0(n256), .Y(n255) );
  NAND4X2 U190 ( .A(n91), .B(n89), .C(n43), .D(n90), .Y(n88) );
  INVX8 U191 ( .A(n275), .Y(n273) );
  NAND2BX1 U192 ( .AN(n71), .B(n273), .Y(n272) );
  OAI21X4 U193 ( .A0(n72), .A1(n65), .B0(n74), .Y(n70) );
  AOI2BB1X2 U194 ( .A0N(n157), .A1N(n158), .B0(n49), .Y(n48) );
  OAI21X4 U195 ( .A0(n82), .A1(n83), .B0(n84), .Y(n79) );
  OR2X1 U196 ( .A(A[24]), .B(B[24]), .Y(n154) );
  CLKINVX2 U197 ( .A(n199), .Y(n184) );
  NOR2BX1 U198 ( .AN(n169), .B(n173), .Y(n181) );
  BUFX12 U199 ( .A(n290), .Y(SUM[21]) );
  NOR2BXL U200 ( .AN(n143), .B(n63), .Y(n147) );
  XOR2X4 U201 ( .A(n149), .B(n150), .Y(SUM[26]) );
  BUFX8 U202 ( .A(n292), .Y(SUM[18]) );
  NAND2X1 U203 ( .A(B[29]), .B(A[29]), .Y(n121) );
  CLKINVX4 U204 ( .A(n55), .Y(n127) );
  OAI21X4 U205 ( .A0(n69), .A1(n70), .B0(n71), .Y(n66) );
  NOR2BX1 U206 ( .AN(n163), .B(n175), .Y(n177) );
  AND2X2 U207 ( .A(n130), .B(n128), .Y(n131) );
  NOR2X2 U208 ( .A(A[20]), .B(B[20]), .Y(n62) );
  NAND2X1 U209 ( .A(B[26]), .B(A[26]), .Y(n137) );
  NOR2X2 U210 ( .A(n113), .B(n61), .Y(n108) );
  AND2X4 U211 ( .A(B[0]), .B(A[0]), .Y(n61) );
  NAND3BX4 U212 ( .AN(n76), .B(n18), .C(n77), .Y(n91) );
  NOR2X4 U213 ( .A(n174), .B(n175), .Y(n171) );
  NAND2X4 U214 ( .A(n153), .B(n154), .Y(n132) );
  OAI21X4 U215 ( .A0(n108), .A1(n109), .B0(n110), .Y(n105) );
  AOI2BB1X1 U216 ( .A0N(n132), .A1N(n133), .B0(n56), .Y(n55) );
  OR2X4 U217 ( .A(n134), .B(n135), .Y(n56) );
  INVXL U218 ( .A(n122), .Y(n119) );
  INVXL U219 ( .A(n190), .Y(n210) );
  NOR2X4 U220 ( .A(n24), .B(n262), .Y(n257) );
  XOR2X4 U221 ( .A(n103), .B(n57), .Y(SUM[5]) );
  AND2X1 U222 ( .A(n43), .B(n94), .Y(n57) );
  AND2X1 U223 ( .A(n89), .B(n95), .Y(n58) );
  INVX8 U224 ( .A(n238), .Y(n225) );
  XOR2X2 U225 ( .A(n117), .B(n59), .Y(SUM[30]) );
  AND2X1 U226 ( .A(n199), .B(n188), .Y(n204) );
  NAND2XL U227 ( .A(n117), .B(n118), .Y(n116) );
  NAND2X1 U228 ( .A(B[22]), .B(A[22]), .Y(n165) );
  NAND2X4 U229 ( .A(B[21]), .B(A[21]), .Y(n169) );
  NAND2XL U230 ( .A(B[27]), .B(A[27]), .Y(n143) );
  NAND2XL U231 ( .A(B[28]), .B(A[28]), .Y(n130) );
  NOR2BX1 U232 ( .AN(n170), .B(n62), .Y(n183) );
  NAND2XL U233 ( .A(n238), .B(n224), .Y(n250) );
  INVX1 U234 ( .A(n2), .Y(n252) );
  OAI2BB1X4 U235 ( .A0N(n166), .A1N(n180), .B0(n169), .Y(n178) );
  NOR2BXL U236 ( .AN(n260), .B(n262), .Y(n269) );
  NOR2BX1 U237 ( .AN(n137), .B(n138), .Y(n150) );
  AOI21XL U238 ( .A0(n160), .A1(n161), .B0(n162), .Y(n159) );
  INVX1 U239 ( .A(n130), .Y(n129) );
  NAND3BX1 U240 ( .AN(n63), .B(n144), .C(n145), .Y(n133) );
  INVX1 U241 ( .A(n143), .Y(n134) );
  INVX1 U242 ( .A(n145), .Y(n140) );
  NAND2X1 U243 ( .A(n121), .B(n122), .Y(n126) );
  XOR2X1 U244 ( .A(n153), .B(n155), .Y(SUM[24]) );
  NOR2BX1 U245 ( .AN(n141), .B(n156), .Y(n155) );
  INVX1 U246 ( .A(n154), .Y(n156) );
  NAND2XL U247 ( .A(n245), .B(n219), .Y(n244) );
  NAND2X1 U248 ( .A(n195), .B(n196), .Y(n193) );
  NAND2X1 U249 ( .A(n115), .B(n116), .Y(n114) );
  INVX1 U250 ( .A(n163), .Y(n162) );
  AND2X2 U251 ( .A(n115), .B(n118), .Y(n59) );
  AOI21X1 U252 ( .A0(n136), .A1(n137), .B0(n63), .Y(n135) );
  NAND2BX1 U253 ( .AN(n138), .B(n139), .Y(n136) );
  OAI21XL U254 ( .A0(n140), .A1(n141), .B0(n142), .Y(n139) );
  NOR2X4 U255 ( .A(A[11]), .B(B[11]), .Y(n60) );
  NAND2X2 U256 ( .A(B[8]), .B(A[8]), .Y(n71) );
  OR2XL U257 ( .A(A[0]), .B(B[0]), .Y(n281) );
  NAND2X2 U258 ( .A(B[16]), .B(A[16]), .Y(n198) );
  XOR3X2 U259 ( .A(B[31]), .B(A[31]), .C(n114), .Y(SUM[31]) );
  NAND2XL U260 ( .A(B[19]), .B(A[19]), .Y(n199) );
  NAND2XL U261 ( .A(B[23]), .B(A[23]), .Y(n163) );
  OR2X2 U262 ( .A(A[26]), .B(B[26]), .Y(n144) );
  OR2X2 U263 ( .A(A[28]), .B(B[28]), .Y(n128) );
  NOR2X1 U264 ( .A(A[27]), .B(B[27]), .Y(n63) );
  NAND2X1 U265 ( .A(B[30]), .B(A[30]), .Y(n115) );
  OR2X2 U266 ( .A(A[30]), .B(B[30]), .Y(n118) );
  NAND2X4 U267 ( .A(n211), .B(n212), .Y(n189) );
  OR2X2 U268 ( .A(A[29]), .B(B[29]), .Y(n122) );
  AOI21X4 U269 ( .A0(n65), .A1(n233), .B0(n234), .Y(n211) );
  XOR2X4 U270 ( .A(n66), .B(n7), .Y(SUM[9]) );
  XOR2X4 U271 ( .A(n79), .B(n80), .Y(SUM[8]) );
  XOR2X4 U272 ( .A(n96), .B(n58), .Y(SUM[6]) );
  OAI21X4 U273 ( .A0(n97), .A1(n98), .B0(n99), .Y(n96) );
  OAI21X4 U274 ( .A0(n104), .A1(n38), .B0(n289), .Y(n103) );
  XOR2X4 U275 ( .A(n105), .B(n106), .Y(SUM[3]) );
  NOR2BX4 U276 ( .AN(n23), .B(n107), .Y(n106) );
  XOR2X4 U277 ( .A(n123), .B(n124), .Y(SUM[2]) );
  XOR2X4 U278 ( .A(n146), .B(n147), .Y(SUM[27]) );
  OAI21X4 U279 ( .A0(n148), .A1(n138), .B0(n137), .Y(n146) );
  XOR2X4 U280 ( .A(n176), .B(n177), .Y(SUM[23]) );
  CLKINVX3 U281 ( .A(n160), .Y(n175) );
  OR2X4 U282 ( .A(A[23]), .B(B[23]), .Y(n160) );
  NAND3BX4 U283 ( .AN(n184), .B(n186), .C(n185), .Y(n182) );
  OAI21X4 U284 ( .A0(n192), .A1(n193), .B0(n194), .Y(n185) );
  XOR2X4 U285 ( .A(n203), .B(n204), .Y(SUM[19]) );
  OR2X4 U286 ( .A(A[18]), .B(B[18]), .Y(n187) );
  XOR2X4 U287 ( .A(n207), .B(n208), .Y(SUM[17]) );
  OR2X4 U288 ( .A(A[17]), .B(B[17]), .Y(n191) );
  OR2X4 U289 ( .A(A[16]), .B(B[16]), .Y(n190) );
  AOI21X4 U290 ( .A0(n213), .A1(n214), .B0(n215), .Y(n212) );
  AOI21X4 U291 ( .A0(n228), .A1(n227), .B0(n83), .Y(n214) );
  NOR2X4 U292 ( .A(n76), .B(n47), .Y(n227) );
  NOR3X4 U293 ( .A(n231), .B(n235), .C(n60), .Y(n234) );
  XOR2X4 U294 ( .A(n239), .B(n240), .Y(SUM[15]) );
  AOI21X4 U295 ( .A0(n45), .A1(n242), .B0(n243), .Y(n240) );
  OR2X4 U296 ( .A(A[15]), .B(B[15]), .Y(n220) );
  XOR2X4 U297 ( .A(n248), .B(n247), .Y(SUM[14]) );
  AOI21X4 U298 ( .A0(n45), .A1(n249), .B0(n50), .Y(n248) );
  OR2X4 U299 ( .A(B[14]), .B(A[14]), .Y(n219) );
  XOR2X4 U300 ( .A(n251), .B(n250), .Y(SUM[13]) );
  AOI21X4 U301 ( .A0(n45), .A1(n237), .B0(n252), .Y(n251) );
  OR2X4 U302 ( .A(B[13]), .B(A[13]), .Y(n238) );
  XOR2X4 U303 ( .A(n45), .B(n253), .Y(SUM[12]) );
  OR2X4 U304 ( .A(B[12]), .B(A[12]), .Y(n237) );
  AOI21X4 U305 ( .A0(n257), .A1(n258), .B0(n259), .Y(n235) );
  NAND2X4 U306 ( .A(n263), .B(n264), .Y(n232) );
  NOR2X4 U307 ( .A(n81), .B(n24), .Y(n264) );
  NOR2X4 U308 ( .A(n262), .B(n60), .Y(n263) );
  XOR2X4 U309 ( .A(n265), .B(n266), .Y(SUM[11]) );
  OAI2BB1X4 U310 ( .A0N(n267), .A1N(n268), .B0(n260), .Y(n265) );
  XOR2X4 U311 ( .A(n30), .B(n269), .Y(SUM[10]) );
  OR2X4 U312 ( .A(B[10]), .B(A[10]), .Y(n267) );
  NAND2X4 U313 ( .A(n276), .B(n277), .Y(n83) );
  OAI2BB1X4 U314 ( .A0N(n22), .A1N(n202), .B0(n229), .Y(n78) );
  NOR2X4 U315 ( .A(n279), .B(n201), .Y(n229) );
  NAND2X4 U316 ( .A(n112), .B(n280), .Y(n279) );
  OR2X4 U317 ( .A(B[2]), .B(A[2]), .Y(n112) );
  NAND3BX4 U318 ( .AN(n283), .B(n284), .C(n285), .Y(n73) );
  NAND3BX4 U319 ( .AN(n39), .B(n17), .C(n286), .Y(n285) );
  NAND2X4 U320 ( .A(n288), .B(n287), .Y(n284) );
  OR2X4 U321 ( .A(B[8]), .B(A[8]), .Y(n74) );
endmodule


module hash_core_DW01_add_49 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331;

  NOR2BXL U2 ( .AN(n226), .B(n63), .Y(n270) );
  NAND2X4 U3 ( .A(n198), .B(n199), .Y(n1) );
  XOR2X4 U4 ( .A(n181), .B(n2), .Y(SUM[27]) );
  CLKINVX20 U5 ( .A(n15), .Y(n2) );
  INVX2 U6 ( .A(n231), .Y(n25) );
  NOR2BX4 U7 ( .AN(n3), .B(A[18]), .Y(n265) );
  CLKINVX20 U8 ( .A(B[18]), .Y(n3) );
  OAI21X4 U9 ( .A0(n301), .A1(n287), .B0(n71), .Y(n299) );
  CLKINVX3 U10 ( .A(n302), .Y(n301) );
  NOR2X4 U11 ( .A(n53), .B(n287), .Y(n286) );
  NAND2X2 U12 ( .A(B[21]), .B(A[21]), .Y(n218) );
  INVX2 U13 ( .A(n242), .Y(n253) );
  INVX2 U14 ( .A(n230), .Y(n31) );
  BUFX12 U15 ( .A(n21), .Y(n63) );
  NAND2BXL U16 ( .AN(n146), .B(n142), .Y(n196) );
  CLKINVX3 U17 ( .A(n21), .Y(n45) );
  INVX4 U18 ( .A(n257), .Y(n61) );
  NOR2X4 U19 ( .A(n47), .B(n204), .Y(n208) );
  INVX4 U20 ( .A(n201), .Y(n209) );
  CLKINVX4 U21 ( .A(n101), .Y(n89) );
  NAND2X2 U22 ( .A(n295), .B(n244), .Y(n282) );
  NAND2X1 U23 ( .A(n118), .B(n122), .Y(n325) );
  NAND2X2 U24 ( .A(B[5]), .B(A[5]), .Y(n118) );
  NOR2X2 U25 ( .A(n100), .B(n14), .Y(n84) );
  CLKINVX3 U26 ( .A(n314), .Y(n100) );
  XNOR2X2 U27 ( .A(n192), .B(n193), .Y(SUM[25]) );
  NOR2BXL U28 ( .AN(n205), .B(n47), .Y(n213) );
  CLKINVX4 U29 ( .A(n291), .Y(n289) );
  NOR2X4 U30 ( .A(n121), .B(n291), .Y(n76) );
  NAND2X4 U31 ( .A(n205), .B(n206), .Y(n202) );
  OR2X4 U32 ( .A(A[14]), .B(B[14]), .Y(n293) );
  NAND2X1 U33 ( .A(B[8]), .B(A[8]), .Y(n103) );
  OR2X2 U34 ( .A(A[8]), .B(B[8]), .Y(n315) );
  NOR2X2 U35 ( .A(n40), .B(B[25]), .Y(n189) );
  INVX4 U36 ( .A(n39), .Y(n40) );
  INVX2 U37 ( .A(n173), .Y(n171) );
  INVX4 U38 ( .A(n107), .Y(n326) );
  NAND2X2 U39 ( .A(B[7]), .B(A[7]), .Y(n107) );
  OAI2BB1X2 U40 ( .A0N(n97), .A1N(n314), .B0(n99), .Y(n320) );
  NAND2X4 U41 ( .A(n322), .B(n103), .Y(n97) );
  CLKINVX8 U42 ( .A(n9), .Y(n238) );
  INVX8 U43 ( .A(n8), .Y(n9) );
  NOR2BX1 U44 ( .AN(n244), .B(n42), .Y(n300) );
  INVX4 U45 ( .A(n244), .Y(n243) );
  INVX1 U46 ( .A(n307), .Y(n30) );
  XNOR2X2 U47 ( .A(n279), .B(n82), .Y(SUM[17]) );
  INVX1 U48 ( .A(n213), .Y(n36) );
  INVX2 U49 ( .A(n42), .Y(n296) );
  INVX1 U50 ( .A(B[25]), .Y(n69) );
  INVX1 U51 ( .A(B[30]), .Y(n54) );
  INVXL U52 ( .A(n171), .Y(n60) );
  NOR2BXL U53 ( .AN(n71), .B(n287), .Y(n303) );
  INVXL U54 ( .A(n29), .Y(n305) );
  INVX1 U55 ( .A(n313), .Y(n312) );
  BUFX3 U56 ( .A(n254), .Y(n37) );
  NOR2BX2 U57 ( .AN(n112), .B(n326), .Y(n323) );
  CLKINVX3 U58 ( .A(n123), .Y(n121) );
  NAND4BBX2 U59 ( .AN(n120), .BN(n93), .C(n115), .D(n109), .Y(n291) );
  OAI2BB1X2 U60 ( .A0N(n116), .A1N(n11), .B0(n118), .Y(n113) );
  BUFX3 U61 ( .A(n206), .Y(n24) );
  INVX1 U62 ( .A(n151), .Y(n81) );
  INVX1 U63 ( .A(n35), .Y(n70) );
  CLKINVX3 U64 ( .A(n43), .Y(n44) );
  NOR2X1 U65 ( .A(n188), .B(n189), .Y(n66) );
  AOI2BB1X1 U66 ( .A0N(n35), .A1N(n184), .B0(n185), .Y(n182) );
  INVX1 U67 ( .A(n116), .Y(n120) );
  NAND2X1 U68 ( .A(A[15]), .B(B[15]), .Y(n244) );
  BUFX3 U69 ( .A(n240), .Y(n71) );
  INVX4 U70 ( .A(n293), .Y(n287) );
  BUFX1 U71 ( .A(A[13]), .Y(n26) );
  NAND2X2 U72 ( .A(n259), .B(n254), .Y(n310) );
  INVX1 U73 ( .A(n315), .Y(n104) );
  NAND2X1 U74 ( .A(B[2]), .B(A[2]), .Y(n131) );
  XNOR2X2 U75 ( .A(n316), .B(n317), .Y(SUM[11]) );
  NAND2X1 U76 ( .A(n313), .B(n319), .Y(n316) );
  NOR2BX2 U77 ( .AN(n151), .B(n161), .Y(n165) );
  NOR2X4 U78 ( .A(n29), .B(n288), .Y(n74) );
  XNOR2X4 U79 ( .A(n190), .B(n94), .Y(SUM[26]) );
  INVX2 U80 ( .A(n273), .Y(n245) );
  AOI21X1 U81 ( .A0(n28), .A1(n242), .B0(n280), .Y(n279) );
  NAND2X2 U82 ( .A(n278), .B(n242), .Y(n277) );
  INVXL U83 ( .A(n248), .Y(n4) );
  AND2X2 U84 ( .A(n177), .B(n178), .Y(n162) );
  INVX4 U85 ( .A(n147), .Y(n178) );
  NOR2X4 U86 ( .A(n209), .B(n210), .Y(n207) );
  XOR2X4 U87 ( .A(n160), .B(n5), .Y(SUM[29]) );
  AND2X2 U88 ( .A(n152), .B(n153), .Y(n5) );
  NAND2X2 U89 ( .A(n194), .B(n180), .Y(n6) );
  NAND2X4 U90 ( .A(n1), .B(n7), .Y(n186) );
  CLKINVX3 U91 ( .A(n6), .Y(n7) );
  OR2X2 U92 ( .A(A[23]), .B(B[23]), .Y(n194) );
  CLKINVX3 U93 ( .A(n186), .Y(n43) );
  NAND3X4 U94 ( .A(n260), .B(n13), .C(n61), .Y(n221) );
  CLKINVX8 U95 ( .A(n249), .Y(n248) );
  INVX8 U96 ( .A(n252), .Y(n8) );
  INVX8 U97 ( .A(n8), .Y(n10) );
  CLKINVX2 U98 ( .A(n227), .Y(n223) );
  BUFX3 U99 ( .A(n117), .Y(n11) );
  AND2X1 U100 ( .A(B[20]), .B(A[20]), .Y(n12) );
  INVX1 U101 ( .A(n200), .Y(n41) );
  AND2X2 U102 ( .A(n242), .B(n79), .Y(n13) );
  NOR2X2 U103 ( .A(A[10]), .B(B[10]), .Y(n14) );
  NAND2X1 U104 ( .A(n60), .B(n144), .Y(n15) );
  AND2X2 U105 ( .A(n211), .B(n201), .Y(n16) );
  INVX1 U106 ( .A(B[29]), .Y(n55) );
  NOR2X2 U107 ( .A(A[12]), .B(B[12]), .Y(n91) );
  NAND3X2 U108 ( .A(n12), .B(n201), .C(n200), .Y(n199) );
  NAND2X1 U109 ( .A(B[14]), .B(A[14]), .Y(n240) );
  INVX8 U110 ( .A(n261), .Y(n255) );
  NOR2X4 U111 ( .A(n218), .B(n204), .Y(n203) );
  NOR2BX2 U112 ( .AN(n145), .B(n167), .Y(n166) );
  NAND2BX2 U113 ( .AN(n42), .B(n10), .Y(n17) );
  NAND2X4 U114 ( .A(B[24]), .B(A[24]), .Y(n175) );
  NAND2X4 U115 ( .A(n45), .B(n20), .Y(n257) );
  NAND2BX4 U116 ( .AN(A[18]), .B(n18), .Y(n92) );
  CLKINVX20 U117 ( .A(B[18]), .Y(n18) );
  NAND3X4 U118 ( .A(n255), .B(n259), .C(n37), .Y(n284) );
  OAI21X4 U119 ( .A0(n168), .A1(n169), .B0(n170), .Y(n19) );
  OR2X2 U120 ( .A(A[20]), .B(B[20]), .Y(n211) );
  NAND2X4 U121 ( .A(B[18]), .B(A[18]), .Y(n273) );
  OR2X4 U122 ( .A(B[18]), .B(A[18]), .Y(n20) );
  NOR2X4 U123 ( .A(A[19]), .B(B[19]), .Y(n21) );
  NAND2X4 U124 ( .A(n49), .B(B[19]), .Y(n226) );
  OAI2BB1X1 U125 ( .A0N(n68), .A1N(n69), .B0(n183), .Y(n193) );
  INVX2 U126 ( .A(n51), .Y(n52) );
  NAND3X4 U127 ( .A(n145), .B(n144), .C(n143), .Y(n163) );
  NAND3X2 U128 ( .A(n145), .B(n144), .C(n19), .Y(n22) );
  CLKINVX3 U129 ( .A(n290), .Y(n77) );
  NOR2BX1 U130 ( .AN(n206), .B(n41), .Y(n216) );
  NAND2X2 U131 ( .A(n19), .B(n144), .Y(n167) );
  AOI2BB1X2 U132 ( .A0N(A[25]), .A1N(B[25]), .B0(n175), .Y(n168) );
  XNOR2X4 U133 ( .A(n23), .B(n195), .Y(SUM[24]) );
  NAND2X2 U134 ( .A(n196), .B(n197), .Y(n23) );
  INVX4 U135 ( .A(n142), .Y(n231) );
  NAND2BX2 U136 ( .AN(n224), .B(n222), .Y(n32) );
  OAI2BB1X4 U137 ( .A0N(n211), .A1N(n142), .B0(n46), .Y(n229) );
  CLKINVX4 U138 ( .A(n278), .Y(n27) );
  INVX4 U139 ( .A(n27), .Y(n28) );
  AOI21X4 U140 ( .A0(n78), .A1(n308), .B0(n30), .Y(n29) );
  AND2X4 U141 ( .A(n48), .B(n142), .Y(n38) );
  OAI2BB1X4 U142 ( .A0N(n48), .A1N(n25), .B0(n166), .Y(n164) );
  XNOR2X4 U143 ( .A(n229), .B(n31), .Y(SUM[21]) );
  NOR2X4 U144 ( .A(n22), .B(n38), .Y(n149) );
  NOR2X4 U145 ( .A(n223), .B(n32), .Y(n72) );
  NAND2X1 U146 ( .A(n174), .B(n95), .Y(n94) );
  INVX1 U147 ( .A(n174), .Y(n185) );
  BUFX1 U148 ( .A(A[19]), .Y(n49) );
  NAND4X2 U149 ( .A(n260), .B(n79), .C(n61), .D(n242), .Y(n33) );
  NAND2XL U150 ( .A(n243), .B(n96), .Y(n34) );
  NAND2X4 U151 ( .A(n219), .B(n16), .Y(n217) );
  OAI21X4 U152 ( .A0(n149), .A1(n50), .B0(n150), .Y(n148) );
  XNOR2X4 U153 ( .A(n214), .B(n216), .Y(SUM[22]) );
  CLKINVX4 U154 ( .A(n215), .Y(n214) );
  NAND2XL U155 ( .A(B[25]), .B(n59), .Y(n35) );
  XOR2X4 U156 ( .A(n231), .B(n232), .Y(SUM[20]) );
  XNOR2X4 U157 ( .A(n212), .B(n36), .Y(SUM[23]) );
  INVX2 U158 ( .A(n59), .Y(n39) );
  INVXL U159 ( .A(A[27]), .Y(n51) );
  NAND4X4 U160 ( .A(n228), .B(n34), .C(n72), .D(n33), .Y(n219) );
  NOR2X4 U161 ( .A(n171), .B(n172), .Y(n170) );
  OR2X4 U162 ( .A(B[22]), .B(A[22]), .Y(n200) );
  NOR2X4 U163 ( .A(A[15]), .B(B[15]), .Y(n42) );
  NOR2X2 U164 ( .A(A[15]), .B(B[15]), .Y(n53) );
  NAND3X4 U165 ( .A(n293), .B(n292), .C(n297), .Y(n239) );
  NAND2X4 U166 ( .A(n92), .B(n242), .Y(n241) );
  OAI21X4 U167 ( .A0(n238), .A1(n250), .B0(n251), .Y(n246) );
  CLKBUFX8 U168 ( .A(n225), .Y(n46) );
  NAND3X2 U169 ( .A(n187), .B(n175), .C(n44), .Y(n67) );
  NAND2X4 U170 ( .A(B[23]), .B(A[23]), .Y(n205) );
  AOI21X4 U171 ( .A0(n142), .A1(n162), .B0(n163), .Y(n134) );
  AND2XL U172 ( .A(n10), .B(n251), .Y(n82) );
  NOR2X4 U173 ( .A(A[23]), .B(B[23]), .Y(n47) );
  NAND2X4 U174 ( .A(n52), .B(B[27]), .Y(n144) );
  NAND2X4 U175 ( .A(n46), .B(n226), .Y(n224) );
  NAND2BX1 U176 ( .AN(n55), .B(A[29]), .Y(n152) );
  NAND2X1 U177 ( .A(B[20]), .B(A[20]), .Y(n225) );
  INVX2 U178 ( .A(n211), .Y(n210) );
  BUFX3 U179 ( .A(n141), .Y(n50) );
  AND2X4 U180 ( .A(n177), .B(n178), .Y(n48) );
  NOR2X1 U181 ( .A(A[4]), .B(B[4]), .Y(n93) );
  NAND2XL U182 ( .A(n194), .B(n1), .Y(n197) );
  NAND2X2 U183 ( .A(n101), .B(n315), .Y(n322) );
  NAND2X4 U184 ( .A(n227), .B(n226), .Y(n234) );
  NAND2X4 U185 ( .A(B[9]), .B(A[9]), .Y(n99) );
  XOR2X2 U186 ( .A(n302), .B(n303), .Y(SUM[14]) );
  OAI2BB1X4 U187 ( .A0N(n200), .A1N(n215), .B0(n24), .Y(n212) );
  INVX4 U188 ( .A(n253), .Y(n62) );
  NAND3X1 U189 ( .A(n116), .B(n115), .C(n325), .Y(n324) );
  NAND3BX4 U190 ( .AN(n262), .B(n263), .C(n255), .Y(n283) );
  NAND2BX4 U191 ( .AN(A[30]), .B(n54), .Y(n138) );
  OAI2BB1X2 U192 ( .A0N(n71), .A1N(n239), .B0(n296), .Y(n295) );
  NAND2BX4 U193 ( .AN(A[29]), .B(n55), .Y(n153) );
  OAI2BB1X4 U194 ( .A0N(B[25]), .A1N(n59), .B0(n174), .Y(n169) );
  XNOR2X4 U195 ( .A(n148), .B(n56), .Y(SUM[30]) );
  NAND2X2 U196 ( .A(n138), .B(n140), .Y(n56) );
  OR2X4 U197 ( .A(n76), .B(n77), .Y(n101) );
  XNOR2X4 U198 ( .A(n133), .B(n57), .Y(SUM[31]) );
  XNOR2X4 U199 ( .A(A[31]), .B(B[31]), .Y(n57) );
  CLKINVX8 U200 ( .A(n58), .Y(n204) );
  NOR2BX1 U201 ( .AN(n99), .B(n100), .Y(n98) );
  INVX2 U202 ( .A(n137), .Y(n150) );
  NOR2X2 U203 ( .A(A[26]), .B(B[26]), .Y(n172) );
  XOR2X4 U204 ( .A(n275), .B(n83), .Y(SUM[18]) );
  OAI21X4 U205 ( .A0(n262), .A1(n89), .B0(n310), .Y(n308) );
  OR2X4 U206 ( .A(A[22]), .B(B[22]), .Y(n58) );
  INVX8 U207 ( .A(n68), .Y(n59) );
  CLKINVX8 U208 ( .A(A[25]), .Y(n68) );
  AND2X1 U209 ( .A(n273), .B(n4), .Y(n83) );
  NAND2XL U210 ( .A(n10), .B(n20), .Y(n272) );
  NAND2X4 U211 ( .A(n220), .B(n222), .Y(n235) );
  NOR2X4 U212 ( .A(n21), .B(n265), .Y(n264) );
  CLKINVX8 U213 ( .A(n146), .Y(n177) );
  NAND2X2 U214 ( .A(n73), .B(n320), .Y(n319) );
  NAND4X4 U215 ( .A(n256), .B(n255), .C(n37), .D(n62), .Y(n228) );
  NOR2X4 U216 ( .A(n17), .B(n63), .Y(n237) );
  NAND2X4 U217 ( .A(n187), .B(n64), .Y(n192) );
  AND2X4 U218 ( .A(n186), .B(n175), .Y(n64) );
  INVX2 U219 ( .A(n140), .Y(n139) );
  NOR2BX4 U220 ( .AN(n251), .B(n274), .Y(n271) );
  OAI21X4 U221 ( .A0(n271), .A1(n272), .B0(n273), .Y(n269) );
  AOI21X4 U222 ( .A0(n137), .A1(n138), .B0(n139), .Y(n136) );
  OAI21X4 U223 ( .A0(n135), .A1(n134), .B0(n136), .Y(n133) );
  BUFX8 U224 ( .A(A[28]), .Y(n65) );
  OAI2BB1X4 U225 ( .A0N(n66), .A1N(n67), .B0(n182), .Y(n181) );
  NOR2X4 U226 ( .A(n257), .B(n258), .Y(n256) );
  INVX4 U227 ( .A(n154), .Y(n161) );
  NAND2X4 U228 ( .A(n80), .B(n176), .Y(n145) );
  OAI2BB1X4 U229 ( .A0N(n39), .A1N(n69), .B0(n192), .Y(n191) );
  NAND2BX4 U230 ( .AN(n70), .B(n191), .Y(n190) );
  XOR2X4 U231 ( .A(n164), .B(n165), .Y(SUM[28]) );
  AOI21X4 U232 ( .A0(n71), .A1(n239), .B0(n241), .Y(n236) );
  AND2X4 U233 ( .A(n263), .B(n9), .Y(n79) );
  NAND2X4 U234 ( .A(B[10]), .B(A[10]), .Y(n313) );
  NAND2BX4 U235 ( .AN(n141), .B(n138), .Y(n135) );
  NAND2X4 U236 ( .A(n153), .B(n154), .Y(n141) );
  OAI2BB1X4 U237 ( .A0N(n81), .A1N(n153), .B0(n152), .Y(n137) );
  XOR2X4 U238 ( .A(n269), .B(n270), .Y(SUM[19]) );
  INVX8 U239 ( .A(n87), .Y(n142) );
  NAND2X4 U240 ( .A(n142), .B(n88), .Y(n187) );
  OR2X4 U241 ( .A(A[10]), .B(B[10]), .Y(n73) );
  NAND2X4 U242 ( .A(B[4]), .B(A[4]), .Y(n122) );
  NAND2XL U243 ( .A(B[1]), .B(A[1]), .Y(n159) );
  OR2XL U244 ( .A(A[2]), .B(B[2]), .Y(n156) );
  NOR2X4 U245 ( .A(n261), .B(n262), .Y(n260) );
  AND2X4 U246 ( .A(n177), .B(n180), .Y(n88) );
  NOR2X4 U247 ( .A(n147), .B(n47), .Y(n80) );
  NOR2X4 U248 ( .A(n63), .B(n248), .Y(n247) );
  XOR2X1 U249 ( .A(n101), .B(n102), .Y(SUM[8]) );
  NAND2X4 U250 ( .A(B[28]), .B(A[28]), .Y(n151) );
  INVXL U251 ( .A(n304), .Y(n75) );
  OR2X4 U252 ( .A(n74), .B(n75), .Y(n302) );
  INVX8 U253 ( .A(n292), .Y(n288) );
  OAI21X4 U254 ( .A0(n245), .A1(n246), .B0(n247), .Y(n227) );
  OAI21X4 U255 ( .A0(n134), .A1(n161), .B0(n151), .Y(n160) );
  INVXL U256 ( .A(n91), .Y(n78) );
  AND3X4 U257 ( .A(n264), .B(n10), .C(n242), .Y(n96) );
  NOR2BX1 U258 ( .AN(n112), .B(n111), .Y(n114) );
  INVX1 U259 ( .A(n157), .Y(n267) );
  OAI2BB1X2 U260 ( .A0N(B[13]), .A1N(A[13]), .B0(n298), .Y(n297) );
  NAND2X2 U261 ( .A(B[6]), .B(A[6]), .Y(n112) );
  NAND2X1 U262 ( .A(B[0]), .B(A[0]), .Y(n268) );
  OAI21X4 U263 ( .A0(n328), .A1(n329), .B0(n127), .Y(n123) );
  NAND2X2 U264 ( .A(n156), .B(n327), .Y(n329) );
  OAI2BB1X4 U265 ( .A0N(n323), .A1N(n324), .B0(n109), .Y(n290) );
  OAI21X1 U266 ( .A0(n110), .A1(n111), .B0(n112), .Y(n105) );
  NOR2BXL U267 ( .AN(n307), .B(n91), .Y(n309) );
  INVXL U268 ( .A(n327), .Y(n128) );
  NOR2BXL U269 ( .AN(n159), .B(n267), .Y(n266) );
  NAND2X4 U270 ( .A(B[16]), .B(A[16]), .Y(n250) );
  NAND2XL U271 ( .A(B[3]), .B(A[3]), .Y(n127) );
  OAI2BB1X4 U272 ( .A0N(n84), .A1N(n85), .B0(n311), .Y(n254) );
  NAND2X2 U273 ( .A(n99), .B(n103), .Y(n85) );
  NOR2BX1 U274 ( .AN(n268), .B(n86), .Y(SUM[0]) );
  NOR2XL U275 ( .A(A[0]), .B(B[0]), .Y(n86) );
  INVX1 U276 ( .A(n132), .Y(n129) );
  INVX1 U277 ( .A(n250), .Y(n280) );
  AND3X4 U278 ( .A(n233), .B(n228), .C(n221), .Y(n87) );
  NAND2XL U279 ( .A(n175), .B(n180), .Y(n195) );
  NOR2X1 U280 ( .A(n330), .B(n331), .Y(n328) );
  NAND2X1 U281 ( .A(n131), .B(n159), .Y(n331) );
  OAI21XL U282 ( .A0(n93), .A1(n121), .B0(n122), .Y(n117) );
  NOR2BXL U283 ( .AN(n218), .B(n209), .Y(n230) );
  NOR2BXL U284 ( .AN(n250), .B(n253), .Y(n281) );
  NOR2X1 U285 ( .A(n267), .B(n268), .Y(n330) );
  NAND2XL U286 ( .A(n46), .B(n211), .Y(n232) );
  NOR2BXL U287 ( .AN(n103), .B(n104), .Y(n102) );
  XOR2X1 U288 ( .A(n320), .B(n321), .Y(SUM[10]) );
  NOR2BX1 U289 ( .AN(n313), .B(n14), .Y(n321) );
  XOR2X1 U290 ( .A(n305), .B(n306), .Y(SUM[13]) );
  NOR2BXL U291 ( .AN(n304), .B(n288), .Y(n306) );
  INVXL U292 ( .A(n109), .Y(n108) );
  XOR2X1 U293 ( .A(n97), .B(n98), .Y(SUM[9]) );
  XOR2X1 U294 ( .A(n308), .B(n309), .Y(SUM[12]) );
  XOR2X1 U295 ( .A(n105), .B(n106), .Y(SUM[7]) );
  NOR2BX1 U296 ( .AN(n107), .B(n108), .Y(n106) );
  INVX1 U297 ( .A(n113), .Y(n110) );
  INVXL U298 ( .A(n115), .Y(n111) );
  XOR2X1 U299 ( .A(n113), .B(n114), .Y(SUM[6]) );
  XOR2X1 U300 ( .A(n123), .B(n124), .Y(SUM[4]) );
  NOR2BX1 U301 ( .AN(n122), .B(n93), .Y(n124) );
  XOR2X1 U302 ( .A(n11), .B(n119), .Y(SUM[5]) );
  NOR2BXL U303 ( .AN(n118), .B(n120), .Y(n119) );
  INVX1 U304 ( .A(n156), .Y(n130) );
  XOR2X1 U305 ( .A(n158), .B(n266), .Y(SUM[1]) );
  OAI2BB1X1 U306 ( .A0N(n157), .A1N(n158), .B0(n159), .Y(n132) );
  INVX1 U307 ( .A(n268), .Y(n158) );
  XOR2X1 U308 ( .A(n132), .B(n155), .Y(SUM[2]) );
  NOR2BX1 U309 ( .AN(n131), .B(n130), .Y(n155) );
  XOR2X1 U310 ( .A(n125), .B(n126), .Y(SUM[3]) );
  NOR2BX1 U311 ( .AN(n127), .B(n128), .Y(n126) );
  OAI21XL U312 ( .A0(n129), .A1(n130), .B0(n131), .Y(n125) );
  NAND4BX4 U313 ( .AN(n179), .B(n90), .C(n173), .D(n180), .Y(n147) );
  OR2X4 U314 ( .A(A[26]), .B(B[26]), .Y(n90) );
  NAND2X2 U315 ( .A(A[22]), .B(B[22]), .Y(n206) );
  NAND2X2 U316 ( .A(A[30]), .B(B[30]), .Y(n140) );
  NAND2X2 U317 ( .A(A[17]), .B(B[17]), .Y(n251) );
  NAND2XL U318 ( .A(B[12]), .B(A[12]), .Y(n307) );
  NAND2XL U319 ( .A(B[13]), .B(n26), .Y(n304) );
  OR2X2 U320 ( .A(A[3]), .B(B[3]), .Y(n327) );
  NAND2XL U321 ( .A(n259), .B(n318), .Y(n317) );
  NAND2XL U322 ( .A(A[11]), .B(B[11]), .Y(n318) );
  OR2X2 U323 ( .A(A[1]), .B(B[1]), .Y(n157) );
  XOR2X1 U324 ( .A(n28), .B(n281), .Y(SUM[16]) );
  OR2XL U325 ( .A(A[26]), .B(B[26]), .Y(n95) );
  NAND2X2 U326 ( .A(n259), .B(n10), .Y(n258) );
  NAND2X2 U327 ( .A(n274), .B(n10), .Y(n276) );
  NOR2XL U328 ( .A(A[26]), .B(B[26]), .Y(n188) );
  NOR2XL U329 ( .A(B[26]), .B(A[26]), .Y(n184) );
  NAND2X2 U330 ( .A(B[26]), .B(A[26]), .Y(n174) );
  NAND2XL U331 ( .A(B[25]), .B(n59), .Y(n183) );
  OR2X4 U332 ( .A(n65), .B(B[28]), .Y(n154) );
  OAI21X4 U333 ( .A0(n168), .A1(n169), .B0(n170), .Y(n143) );
  NOR2X4 U334 ( .A(A[25]), .B(B[25]), .Y(n179) );
  OR2X4 U335 ( .A(A[27]), .B(B[27]), .Y(n173) );
  OR2X4 U336 ( .A(A[24]), .B(B[24]), .Y(n180) );
  NAND2X4 U337 ( .A(n199), .B(n198), .Y(n176) );
  NOR2X4 U338 ( .A(n203), .B(n202), .Y(n198) );
  NAND2X4 U339 ( .A(n207), .B(n208), .Y(n146) );
  NAND2X4 U340 ( .A(n217), .B(n218), .Y(n215) );
  OR2X4 U341 ( .A(A[21]), .B(B[21]), .Y(n201) );
  NOR2X4 U342 ( .A(n235), .B(n234), .Y(n233) );
  NAND2X4 U343 ( .A(n237), .B(n236), .Y(n222) );
  NAND2X4 U344 ( .A(n96), .B(n243), .Y(n220) );
  OR2X4 U345 ( .A(A[18]), .B(B[18]), .Y(n249) );
  NAND2X4 U346 ( .A(n251), .B(n276), .Y(n275) );
  NAND2X4 U347 ( .A(n277), .B(n250), .Y(n274) );
  OR2X4 U348 ( .A(A[17]), .B(B[17]), .Y(n252) );
  OR2X4 U349 ( .A(A[16]), .B(B[16]), .Y(n242) );
  NAND3BX4 U350 ( .AN(n282), .B(n283), .C(n284), .Y(n278) );
  NAND2X4 U351 ( .A(n286), .B(n285), .Y(n261) );
  NOR2X4 U352 ( .A(n288), .B(n91), .Y(n285) );
  OAI2BB1X4 U353 ( .A0N(n289), .A1N(n123), .B0(n290), .Y(n263) );
  NAND2X4 U354 ( .A(B[12]), .B(A[12]), .Y(n298) );
  XOR2X4 U355 ( .A(n299), .B(n300), .Y(SUM[15]) );
  OR2X4 U356 ( .A(A[13]), .B(B[13]), .Y(n292) );
  AOI21X4 U357 ( .A0(B[11]), .A1(A[11]), .B0(n312), .Y(n311) );
  NAND4BX4 U358 ( .AN(n104), .B(n314), .C(n73), .D(n294), .Y(n262) );
  OR2X4 U359 ( .A(A[11]), .B(B[11]), .Y(n294) );
  OR2X4 U360 ( .A(A[11]), .B(B[11]), .Y(n259) );
  OR2X4 U361 ( .A(A[9]), .B(B[9]), .Y(n314) );
  OR2X4 U362 ( .A(A[7]), .B(B[7]), .Y(n109) );
  OR2X4 U363 ( .A(A[6]), .B(B[6]), .Y(n115) );
  OR2X4 U364 ( .A(A[5]), .B(B[5]), .Y(n116) );
endmodule


module hash_core ( clk, reset, Wt, inner_busy, first_block_core, output_enable, 
        digest, output_valid );
  input [31:0] Wt;
  output [3:0] digest;
  input clk, reset, inner_busy, first_block_core, output_enable;
  output output_valid;
  wire   mux_control_0_, N152, N153, N154, N155, N156, N157, N158, N841, N842,
         N843, N844, N845, N846, N847, N848, N849, N850, N851, N852, N853,
         N854, N855, N856, N857, N858, N859, N860, N861, N862, N863, N864,
         N865, N866, N867, N868, N869, N870, N871, N872, N873, N874, N875,
         N876, N877, N878, N879, N880, N881, N882, N883, N884, N885, N886,
         N887, N888, N889, N890, N891, N892, N893, N894, N895, N896, N897,
         N898, N899, N900, N901, N902, N903, N904, N905, N906, N907, N908,
         N909, N910, N911, N912, N913, N914, N915, N916, N917, N918, N919,
         N920, N921, N922, N923, N924, N925, N926, N927, N928, N929, N930,
         N931, N932, N933, N934, N935, N936, N937, N938, N939, N940, N941,
         N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952,
         N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963,
         N964, N965, N966, N967, N968, N969, N970, N971, N972, N973, N974,
         N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985,
         N986, N987, N988, N989, N990, N991, N992, N993, N994, N995, N996,
         N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006,
         N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016,
         N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026,
         N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036,
         N1037, N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046,
         N1047, N1048, N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056,
         N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066,
         N1067, N1068, N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076,
         N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086,
         N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096,
         N3133, N3134, N3135, N3136, N3137, N3138, N3139, N3140, N3141, N3142,
         N3143, N3144, N3145, N3146, N3147, N3148, N3149, N3150, N3151, N3152,
         N3153, N3154, N3155, N3156, N3157, N3158, N3159, N3160, N3161, N3162,
         N3163, N3164, N3564, N3565, N3566, N3575, N3576, N3577, N3578, N3579,
         N3580, N3581, N3582, N3583, N3584, n2878, n2906, n2925, n2938, n2943,
         n2946, n2947, n3114, n3115, n3116, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3377, n3378, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3564, n3574, n3576, n3577,
         n3578, n3579, n3580, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3881, n3882, n3883, n3885,
         n3886, n3887, n3888, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3943, n3944, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3975, n3976, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N118,
         N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107,
         N106, N105, N104, N103, N102, N101, N100, N150, N149, N148, N147,
         N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136,
         N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125,
         N124, N123, N122, N121, N120, N119, T2_32_9_, T2_32_8_, T2_32_7_,
         T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_, T2_32_31_, T2_32_30_,
         T2_32_2_, T2_32_29_, T2_32_28_, T2_32_27_, T2_32_26_, T2_32_25_,
         T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_, T2_32_20_, T2_32_1_,
         T2_32_19_, T2_32_18_, T2_32_17_, T2_32_16_, T2_32_15_, T2_32_14_,
         T2_32_13_, T2_32_12_, T2_32_11_, T2_32_10_, T2_32_0_, n11, n12, n14,
         n15, n16, n17, n18, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n217, n218, n219, n220, n221, n222, n226, n229, n230, n231, n232,
         n233, n234, n235, n237, n238, n239, n243, n244, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n264, n265, n266, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431;
  wire   [31:0] f1_EFG_32;
  wire   [31:0] f2_ABC_32;
  wire   [31:0] f3_A_32;
  wire   [31:0] f4_E_32;
  wire   [31:0] mux2;
  wire   [31:0] mux1;
  wire   [31:0] Kt;
  wire   [31:0] M_w;
  wire   [31:0] M;
  wire   [31:0] T1_32;
  wire   [31:0] next_E;
  wire   [31:0] L;
  wire   [31:0] next_A;
  wire   [255:0] SHA256_result;
  wire   [6:0] round;
  wire   [31:0] H0;
  wire   [31:0] H1;
  wire   [31:0] H2;
  wire   [31:0] H3;
  wire   [31:0] H4;
  wire   [31:0] H5;
  wire   [31:0] H6;
  wire   [31:0] H7;
  wire   [5:0] read_counter;

  DFFTRX4 M_reg_7_ ( .D(M_w[7]), .RN(n402), .CK(clk), .Q(M[7]) );
  DFFHQX4 A_reg_0_ ( .D(n4764), .CK(clk), .Q(SHA256_result[224]) );
  DFFHQX4 A_reg_1_ ( .D(n4763), .CK(clk), .Q(SHA256_result[225]) );
  DFFHQX4 A_reg_2_ ( .D(n4762), .CK(clk), .Q(SHA256_result[226]) );
  DFFHQX4 A_reg_4_ ( .D(n4760), .CK(clk), .Q(SHA256_result[228]) );
  DFFHQX4 A_reg_5_ ( .D(n4759), .CK(clk), .Q(SHA256_result[229]) );
  DFFHQX4 A_reg_6_ ( .D(n4758), .CK(clk), .Q(SHA256_result[230]) );
  DFFHQX4 A_reg_8_ ( .D(n4756), .CK(clk), .Q(SHA256_result[232]) );
  DFFHQX4 A_reg_9_ ( .D(n4755), .CK(clk), .Q(SHA256_result[233]) );
  DFFHQX4 A_reg_11_ ( .D(n4753), .CK(clk), .Q(SHA256_result[235]) );
  DFFHQX4 A_reg_12_ ( .D(n4752), .CK(clk), .Q(SHA256_result[236]) );
  DFFHQX4 A_reg_13_ ( .D(n4751), .CK(clk), .Q(SHA256_result[237]) );
  DFFHQX4 A_reg_15_ ( .D(n4749), .CK(clk), .Q(SHA256_result[239]) );
  DFFHQX4 B_reg_1_ ( .D(n4697), .CK(clk), .Q(SHA256_result[193]) );
  DFFHQX4 B_reg_4_ ( .D(n4694), .CK(clk), .Q(SHA256_result[196]) );
  DFFHQX4 B_reg_5_ ( .D(n4693), .CK(clk), .Q(SHA256_result[197]) );
  DFFHQX4 B_reg_6_ ( .D(n4692), .CK(clk), .Q(SHA256_result[198]) );
  DFFHQX4 B_reg_7_ ( .D(n4691), .CK(clk), .Q(SHA256_result[199]) );
  DFFHQX4 B_reg_8_ ( .D(n4690), .CK(clk), .Q(SHA256_result[200]) );
  DFFHQX4 B_reg_9_ ( .D(n4689), .CK(clk), .Q(SHA256_result[201]) );
  DFFHQX4 B_reg_10_ ( .D(n4688), .CK(clk), .Q(SHA256_result[202]) );
  DFFHQX4 B_reg_11_ ( .D(n4687), .CK(clk), .Q(SHA256_result[203]) );
  DFFHQX4 B_reg_12_ ( .D(n4686), .CK(clk), .Q(SHA256_result[204]) );
  DFFHQX4 B_reg_13_ ( .D(n4685), .CK(clk), .Q(SHA256_result[205]) );
  DFFHQX4 B_reg_14_ ( .D(n4684), .CK(clk), .Q(SHA256_result[206]) );
  DFFHQX4 B_reg_15_ ( .D(n4683), .CK(clk), .Q(SHA256_result[207]) );
  DFFHQX4 C_reg_0_ ( .D(n4666), .CK(clk), .Q(SHA256_result[160]) );
  DFFHQX4 C_reg_1_ ( .D(n4665), .CK(clk), .Q(SHA256_result[161]) );
  DFFHQX4 C_reg_2_ ( .D(n4664), .CK(clk), .Q(SHA256_result[162]) );
  DFFHQX4 C_reg_3_ ( .D(n4663), .CK(clk), .Q(SHA256_result[163]) );
  DFFHQX4 C_reg_4_ ( .D(n4662), .CK(clk), .Q(SHA256_result[164]) );
  DFFHQX4 C_reg_5_ ( .D(n4661), .CK(clk), .Q(SHA256_result[165]) );
  DFFHQX4 C_reg_6_ ( .D(n4660), .CK(clk), .Q(SHA256_result[166]) );
  DFFHQX4 C_reg_7_ ( .D(n4659), .CK(clk), .Q(SHA256_result[167]) );
  DFFHQX4 C_reg_8_ ( .D(n4658), .CK(clk), .Q(SHA256_result[168]) );
  DFFHQX4 C_reg_9_ ( .D(n4657), .CK(clk), .Q(SHA256_result[169]) );
  DFFHQX4 C_reg_12_ ( .D(n4654), .CK(clk), .Q(SHA256_result[172]) );
  DFFHQX4 C_reg_13_ ( .D(n4653), .CK(clk), .Q(SHA256_result[173]) );
  DFFHQX4 C_reg_14_ ( .D(n4652), .CK(clk), .Q(SHA256_result[174]) );
  DFFHQX4 C_reg_15_ ( .D(n4651), .CK(clk), .Q(SHA256_result[175]) );
  DFFHQX4 E_reg_0_ ( .D(n4570), .CK(clk), .Q(SHA256_result[96]) );
  DFFHQX4 E_reg_2_ ( .D(n4568), .CK(clk), .Q(SHA256_result[98]) );
  DFFHQX4 E_reg_4_ ( .D(n4566), .CK(clk), .Q(SHA256_result[100]) );
  DFFHQX4 E_reg_8_ ( .D(n4562), .CK(clk), .Q(SHA256_result[104]) );
  DFFHQX4 E_reg_9_ ( .D(n4561), .CK(clk), .Q(SHA256_result[105]) );
  DFFHQX4 E_reg_12_ ( .D(n4558), .CK(clk), .Q(SHA256_result[108]) );
  DFFHQX4 E_reg_13_ ( .D(n4557), .CK(clk), .Q(SHA256_result[109]) );
  DFFHQX4 E_reg_15_ ( .D(n4555), .CK(clk), .Q(SHA256_result[111]) );
  DFFHQX4 E_reg_16_ ( .D(n4554), .CK(clk), .Q(SHA256_result[112]) );
  DFFHQX4 E_reg_20_ ( .D(n4550), .CK(clk), .Q(SHA256_result[116]) );
  DFFHQX4 E_reg_21_ ( .D(n4549), .CK(clk), .Q(SHA256_result[117]) );
  DFFHQX4 E_reg_22_ ( .D(n4548), .CK(clk), .Q(SHA256_result[118]) );
  DFFHQX4 F_reg_1_ ( .D(n4442), .CK(clk), .Q(SHA256_result[65]) );
  DFFHQX4 F_reg_3_ ( .D(n4440), .CK(clk), .Q(SHA256_result[67]) );
  DFFHQX4 F_reg_4_ ( .D(n4439), .CK(clk), .Q(SHA256_result[68]) );
  DFFHQX4 F_reg_8_ ( .D(n4435), .CK(clk), .Q(SHA256_result[72]) );
  DFFHQX4 F_reg_9_ ( .D(n4434), .CK(clk), .Q(SHA256_result[73]) );
  DFFHQX4 F_reg_10_ ( .D(n4433), .CK(clk), .Q(SHA256_result[74]) );
  DFFHQX4 F_reg_11_ ( .D(n4432), .CK(clk), .Q(SHA256_result[75]) );
  DFFHQX4 F_reg_12_ ( .D(n4431), .CK(clk), .Q(SHA256_result[76]) );
  DFFHQX4 F_reg_13_ ( .D(n4430), .CK(clk), .Q(SHA256_result[77]) );
  DFFHQX4 F_reg_14_ ( .D(n4429), .CK(clk), .Q(SHA256_result[78]) );
  DFFHQX4 F_reg_15_ ( .D(n4428), .CK(clk), .Q(SHA256_result[79]) );
  DFFHQX4 G_reg_3_ ( .D(n4408), .CK(clk), .Q(SHA256_result[35]) );
  DFFHQX4 G_reg_6_ ( .D(n4405), .CK(clk), .Q(SHA256_result[38]) );
  DFFHQX4 G_reg_8_ ( .D(n4403), .CK(clk), .Q(SHA256_result[40]) );
  DFFHQX4 G_reg_11_ ( .D(n4400), .CK(clk), .Q(SHA256_result[43]) );
  DFFHQX4 G_reg_12_ ( .D(n4399), .CK(clk), .Q(SHA256_result[44]) );
  DFFHQX4 G_reg_13_ ( .D(n4398), .CK(clk), .Q(SHA256_result[45]) );
  DFFHQX4 G_reg_14_ ( .D(n4397), .CK(clk), .Q(SHA256_result[46]) );
  DFFHQX4 G_reg_15_ ( .D(n4396), .CK(clk), .Q(SHA256_result[47]) );
  AND2X2 U1409 ( .A(n3879), .B(n78), .Y(n3691) );
  AND2X2 U1410 ( .A(n3881), .B(n78), .Y(n3690) );
  AND2X2 U1412 ( .A(n3882), .B(n78), .Y(n3693) );
  AND2X2 U1413 ( .A(n3883), .B(n78), .Y(n3692) );
  AND2X2 U1415 ( .A(n3879), .B(n80), .Y(n3695) );
  AND2X2 U1416 ( .A(n3881), .B(n80), .Y(n3694) );
  AND2X2 U1418 ( .A(n3882), .B(n80), .Y(n3697) );
  AND2X2 U1419 ( .A(n3883), .B(n80), .Y(n3696) );
  AND2X2 U1422 ( .A(n3879), .B(n79), .Y(n3703) );
  AND2X2 U1423 ( .A(n3881), .B(n79), .Y(n3702) );
  AND2X2 U1425 ( .A(n3882), .B(n79), .Y(n3705) );
  AND2X2 U1426 ( .A(n3883), .B(n79), .Y(n3704) );
  AND2X2 U1428 ( .A(n3879), .B(n77), .Y(n3707) );
  AND2X2 U1429 ( .A(n3891), .B(n3892), .Y(n3879) );
  AND2X2 U1430 ( .A(n3881), .B(n77), .Y(n3706) );
  AND2X2 U1431 ( .A(n3891), .B(n3893), .Y(n3881) );
  AND2X2 U1433 ( .A(n3882), .B(n77), .Y(n3709) );
  AND2X2 U1434 ( .A(n3894), .B(n3892), .Y(n3882) );
  AND2X2 U1435 ( .A(n3883), .B(n77), .Y(n3708) );
  AND2X2 U1436 ( .A(n3894), .B(n3893), .Y(n3883) );
  AND2X2 U1439 ( .A(n78), .B(n3899), .Y(n3715) );
  AND2X2 U1440 ( .A(n78), .B(n3900), .Y(n3714) );
  AND2X2 U1442 ( .A(n78), .B(n3901), .Y(n3717) );
  AND2X2 U1443 ( .A(n78), .B(n3902), .Y(n3716) );
  AND2X2 U1445 ( .A(n80), .B(n3899), .Y(n3719) );
  AND2X2 U1446 ( .A(n80), .B(n3900), .Y(n3718) );
  AND2X2 U1448 ( .A(n80), .B(n3901), .Y(n3721) );
  AND2X2 U1449 ( .A(n80), .B(n3902), .Y(n3720) );
  AND2X2 U1452 ( .A(n3899), .B(n79), .Y(n3726) );
  AND2X2 U1453 ( .A(n79), .B(n3900), .Y(n3679) );
  AND2X2 U1455 ( .A(n3901), .B(n79), .Y(n3728) );
  AND2X2 U1456 ( .A(n3902), .B(n79), .Y(n3727) );
  AND2X2 U1458 ( .A(n77), .B(n3899), .Y(n3730) );
  AND2X2 U1459 ( .A(n3892), .B(n3907), .Y(n3899) );
  AND2X2 U1460 ( .A(n77), .B(n3900), .Y(n3729) );
  AND2X2 U1461 ( .A(n3893), .B(n3907), .Y(n3900) );
  AND2X2 U1463 ( .A(n77), .B(n3901), .Y(n3732) );
  AND2X2 U1464 ( .A(n3908), .B(n3892), .Y(n3901) );
  AND2X2 U1465 ( .A(read_counter[0]), .B(n1431), .Y(n3892) );
  AND2X2 U1466 ( .A(n77), .B(n3902), .Y(n3731) );
  AND2X2 U1467 ( .A(n3908), .B(n3893), .Y(n3902) );
  AND2X2 U1472 ( .A(n3917), .B(n78), .Y(n3742) );
  AND2X2 U1473 ( .A(n3918), .B(n78), .Y(n3741) );
  AND2X2 U1475 ( .A(n3919), .B(n78), .Y(n3744) );
  AND2X2 U1476 ( .A(n3920), .B(n78), .Y(n3743) );
  AND2X2 U1478 ( .A(n3917), .B(n80), .Y(n3746) );
  AND2X2 U1479 ( .A(n3918), .B(n80), .Y(n3745) );
  AND2X2 U1481 ( .A(n3919), .B(n80), .Y(n3748) );
  AND2X2 U1482 ( .A(n3920), .B(n80), .Y(n3747) );
  AND2X2 U1485 ( .A(n3917), .B(n79), .Y(n3754) );
  AND2X2 U1486 ( .A(n3918), .B(n79), .Y(n3753) );
  AND2X2 U1488 ( .A(n3919), .B(n79), .Y(n3756) );
  AND2X2 U1489 ( .A(n3920), .B(n79), .Y(n3755) );
  AND2X2 U1491 ( .A(n3917), .B(n77), .Y(n3758) );
  AND2X2 U1492 ( .A(n3925), .B(n3891), .Y(n3917) );
  AND2X2 U1493 ( .A(n3918), .B(n77), .Y(n3757) );
  AND2X2 U1494 ( .A(n3926), .B(n3891), .Y(n3918) );
  AND2X2 U1495 ( .A(read_counter[4]), .B(n1429), .Y(n3891) );
  AND2X2 U1497 ( .A(n3919), .B(n77), .Y(n3760) );
  AND2X2 U1498 ( .A(n3925), .B(n3894), .Y(n3919) );
  AND2X2 U1499 ( .A(n3920), .B(n77), .Y(n3759) );
  AND2X2 U1500 ( .A(n3926), .B(n3894), .Y(n3920) );
  AND2X2 U1501 ( .A(read_counter[4]), .B(read_counter[1]), .Y(n3894) );
  AND2X2 U1504 ( .A(n3931), .B(n78), .Y(n3766) );
  AND2X2 U1505 ( .A(n3932), .B(n78), .Y(n3765) );
  AND2X2 U1507 ( .A(n3933), .B(n78), .Y(n3768) );
  AND2X2 U1508 ( .A(n3934), .B(n78), .Y(n3767) );
  AND2X2 U1511 ( .A(n3931), .B(n80), .Y(n3770) );
  AND2X2 U1512 ( .A(n3932), .B(n80), .Y(n3769) );
  AND2X2 U1514 ( .A(n3933), .B(n80), .Y(n3772) );
  AND2X2 U1515 ( .A(n3934), .B(n80), .Y(n3771) );
  AND2X2 U1519 ( .A(n3931), .B(n79), .Y(n3778) );
  AND2X2 U1520 ( .A(n3932), .B(n79), .Y(n3777) );
  AND2X2 U1522 ( .A(n3933), .B(n79), .Y(n3780) );
  AND2X2 U1523 ( .A(n3934), .B(n79), .Y(n3779) );
  AND2X2 U1526 ( .A(n3931), .B(n77), .Y(n3782) );
  AND2X2 U1527 ( .A(n3925), .B(n3907), .Y(n3931) );
  AND2X2 U1528 ( .A(n3932), .B(n77), .Y(n3781) );
  AND2X2 U1529 ( .A(n3926), .B(n3907), .Y(n3932) );
  AND2X2 U1532 ( .A(n3933), .B(n77), .Y(n3784) );
  AND2X2 U1533 ( .A(n3925), .B(n3908), .Y(n3933) );
  AND2X2 U1534 ( .A(read_counter[0]), .B(read_counter[5]), .Y(n3925) );
  AND2X2 U1535 ( .A(n3934), .B(n77), .Y(n3783) );
  AND2X2 U1537 ( .A(n3926), .B(n3908), .Y(n3934) );
  CLKINVX4 U2229 ( .A(reset), .Y(n3114) );
  hash_core_DW01_inc_0 add_132 ( .A({round[6], n434, n318, n319, n431, n320, 
        n423}), .SUM({N158, N157, N156, N155, N154, N153, N152}) );
  hash_core_DW01_add_16 add_406 ( .A(next_A), .B(H0), .SUM({N1096, N1095, 
        N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, 
        N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, 
        N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065})
         );
  hash_core_DW01_add_24 add_0_root_add_0_root_add_126 ( .A(f3_A_32), .B({
        T2_32_31_, T2_32_30_, T2_32_29_, T2_32_28_, T2_32_27_, T2_32_26_, 
        T2_32_25_, T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_, T2_32_20_, 
        T2_32_19_, T2_32_18_, T2_32_17_, T2_32_16_, T2_32_15_, T2_32_14_, 
        T2_32_13_, T2_32_12_, T2_32_11_, T2_32_10_, T2_32_9_, T2_32_8_, 
        T2_32_7_, T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_, T2_32_2_, T2_32_1_, 
        T2_32_0_}), .SUM(next_A) );
  hash_core_DW01_add_26 add_125 ( .A(mux1), .B({T1_32[31:22], n17, T1_32[20:0]}), .SUM(next_E) );
  hash_core_DW01_add_29 add_378 ( .A({SHA256_result[63:57], n119, 
        SHA256_result[55:43], n159, n165, n184, n134, n143, n174, n140, n208, 
        n234, n164, n232}), .B(H7), .SUM({N872, N871, N870, N869, N868, N867, 
        N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, 
        N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, 
        N842, N841}) );
  hash_core_DW01_add_28 add_405 ( .A({n293, n294, n295, n296, n297, n298, n299, 
        n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, 
        SHA256_result[237:236], n15, n311, n312, n18, n219, n313, n314, 
        SHA256_result[228], n222, n315, n316, n317}), .B(H1), .SUM({N1064, 
        N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, 
        N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, 
        N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, 
        N1033}) );
  hash_core_DW01_add_33 add_380 ( .A({n106, n115, n110, n94, n123, n118, n244, 
        n103, n90, SHA256_result[118:116], n111, n291, SHA256_result[113:112], 
        n280, n203, n171, n146, n139, n127, n281, n210, n154, n136, n150, 
        SHA256_result[100], n283, n282, n158, n285}), .B(H5), .SUM({N936, N935, 
        N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, 
        N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, 
        N910, N909, N908, N907, N906, N905}) );
  hash_core_DW01_add_32 add_403 ( .A({SHA256_result[191:186], n86, 
        SHA256_result[184:179], n32, SHA256_result[177:160]}), .B(H3), .SUM({
        N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, 
        N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, 
        N977, N976, N975, N974, N973, N972, N971, N970, N969}) );
  hash_core_DW01_add_31 add_404 ( .A({SHA256_result[223:196], n100, 
        SHA256_result[194:193], n96}), .B(H2), .SUM({N1032, N1031, N1030, 
        N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, 
        N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, 
        N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001}) );
  hash_core_DW01_add_34 add_379 ( .A({SHA256_result[95:89], n31, 
        SHA256_result[87:75], n81, n11, n85, n167, n84, n130, 
        SHA256_result[68], n207, n213, n181, n239}), .B(H6), .SUM({N904, N903, 
        N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, 
        N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, 
        N878, N877, N876, N875, N874, N873}) );
  hash_core_DW01_add_27 add_0_root_add_0_root_add_118_2 ( .A(mux2), .B({N118, 
        N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, 
        N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, 
        N92, N91, N90, N89, N88, N87}), .SUM(M_w) );
  hash_core_DW01_add_35 add_1_root_add_0_root_add_118_2 ( .A(Kt), .B(Wt), 
        .SUM({N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, 
        N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, 
        N95, N94, N93, N92, N91, N90, N89, N88, N87}) );
  hash_core_DW01_add_38 add_0_root_add_0_root_add_121_2 ( .A(f4_E_32), .B({
        N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, 
        N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, 
        N126, N125, N124, N123, N122, N121, N120, N119}), .SUM(T1_32) );
  hash_core_DW01_add_40 add_1_root_add_0_root_add_126 ( .A(L), .B(f2_ABC_32), 
        .SUM({T2_32_31_, T2_32_30_, T2_32_29_, T2_32_28_, T2_32_27_, T2_32_26_, 
        T2_32_25_, T2_32_24_, T2_32_23_, T2_32_22_, T2_32_21_, T2_32_20_, 
        T2_32_19_, T2_32_18_, T2_32_17_, T2_32_16_, T2_32_15_, T2_32_14_, 
        T2_32_13_, T2_32_12_, T2_32_11_, T2_32_10_, T2_32_9_, T2_32_8_, 
        T2_32_7_, T2_32_6_, T2_32_5_, T2_32_4_, T2_32_3_, T2_32_2_, T2_32_1_, 
        T2_32_0_}) );
  hash_core_DW01_add_43 add_1_root_add_0_root_add_121_2 ( .A(M), .B({
        f1_EFG_32[31:1], n284}), .SUM({N150, N149, N148, N147, N146, N145, 
        N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, 
        N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, 
        N120, N119}) );
  hash_core_DW01_add_49 add_381 ( .A({next_E[31:27], n209, next_E[25:11], n186, 
        next_E[9:0]}), .B(H4), .SUM({N968, N967, N966, N965, N964, N963, N962, 
        N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, 
        N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, 
        N937}) );
  DFFHQX1 Kt_reg_31_ ( .D(N3164), .CK(clk), .Q(Kt[31]) );
  DFFHQX1 Kt_reg_30_ ( .D(N3163), .CK(clk), .Q(Kt[30]) );
  DFFTRX1 L_reg_31_ ( .D(T1_32[31]), .RN(n402), .CK(clk), .Q(L[31]) );
  DFFHQX1 Kt_reg_29_ ( .D(N3162), .CK(clk), .Q(Kt[29]) );
  DFFHQX1 read_counter_reg_5_ ( .D(N3584), .CK(clk), .Q(read_counter[5]) );
  DFFHQX1 read_counter_reg_1_ ( .D(N3580), .CK(clk), .Q(read_counter[1]) );
  DFFHQX1 read_counter_reg_2_ ( .D(N3581), .CK(clk), .Q(read_counter[2]) );
  DFFHQX1 read_counter_reg_3_ ( .D(N3582), .CK(clk), .Q(read_counter[3]) );
  DFFHQX1 read_counter_reg_4_ ( .D(N3583), .CK(clk), .Q(read_counter[4]) );
  DFFHQX1 read_counter_reg_0_ ( .D(N3579), .CK(clk), .Q(read_counter[0]) );
  DFFTRX1 L_reg_30_ ( .D(T1_32[30]), .RN(n402), .CK(clk), .Q(L[30]) );
  DFFTRX1 L_reg_29_ ( .D(T1_32[29]), .RN(n402), .CK(clk), .Q(L[29]) );
  DFFTRX1 L_reg_28_ ( .D(T1_32[28]), .RN(n402), .CK(clk), .Q(L[28]) );
  DFFHQX1 Kt_reg_27_ ( .D(N3160), .CK(clk), .Q(Kt[27]) );
  DFFHQX1 Kt_reg_26_ ( .D(N3159), .CK(clk), .Q(Kt[26]) );
  DFFHQX1 Kt_reg_24_ ( .D(N3157), .CK(clk), .Q(Kt[24]) );
  DFFHQX1 H0_reg_3_ ( .D(n4730), .CK(clk), .Q(H0[3]) );
  DFFTRX1 L_reg_26_ ( .D(T1_32[26]), .RN(n403), .CK(clk), .Q(L[26]) );
  DFFTRX1 L_reg_24_ ( .D(T1_32[24]), .RN(n403), .CK(clk), .Q(L[24]) );
  DFFHQX1 Kt_reg_23_ ( .D(N3156), .CK(clk), .Q(Kt[23]) );
  DFFHQX1 Kt_reg_22_ ( .D(N3155), .CK(clk), .Q(Kt[22]) );
  DFFHQX1 Kt_reg_21_ ( .D(N3154), .CK(clk), .Q(Kt[21]) );
  DFFHQX1 Kt_reg_20_ ( .D(N3153), .CK(clk), .Q(Kt[20]) );
  DFFHQX1 Kt_reg_19_ ( .D(N3152), .CK(clk), .Q(Kt[19]) );
  DFFHQX1 Kt_reg_18_ ( .D(N3151), .CK(clk), .Q(Kt[18]) );
  DFFHQX1 Kt_reg_17_ ( .D(N3150), .CK(clk), .Q(Kt[17]) );
  DFFHQX1 Kt_reg_16_ ( .D(N3149), .CK(clk), .Q(Kt[16]) );
  DFFTRX2 round_reg_3_ ( .D(N155), .RN(n4250), .CK(clk), .Q(round[3]), .QN(
        n2938) );
  DFFTRX2 round_reg_4_ ( .D(N156), .RN(n4250), .CK(clk), .Q(round[4]), .QN(
        n2925) );
  DFFHQXL A_reg_26_ ( .D(n4738), .CK(clk), .Q(SHA256_result[250]) );
  DFFHQXL A_reg_29_ ( .D(n4735), .CK(clk), .Q(SHA256_result[253]) );
  DFFHQXL A_reg_30_ ( .D(n4734), .CK(clk), .Q(SHA256_result[254]) );
  DFFHQXL A_reg_31_ ( .D(n4733), .CK(clk), .Q(SHA256_result[255]) );
  DFFHQX1 Kt_reg_15_ ( .D(N3148), .CK(clk), .Q(Kt[15]) );
  DFFHQX1 Kt_reg_14_ ( .D(N3147), .CK(clk), .Q(Kt[14]) );
  DFFHQX1 Kt_reg_13_ ( .D(N3146), .CK(clk), .Q(Kt[13]) );
  DFFHQX1 Kt_reg_12_ ( .D(N3145), .CK(clk), .Q(Kt[12]) );
  DFFHQX1 Kt_reg_11_ ( .D(N3144), .CK(clk), .Q(Kt[11]) );
  DFFHQX1 Kt_reg_10_ ( .D(N3143), .CK(clk), .Q(Kt[10]) );
  DFFHQX1 Kt_reg_9_ ( .D(N3142), .CK(clk), .Q(Kt[9]) );
  DFFHQX1 Kt_reg_8_ ( .D(N3141), .CK(clk), .Q(Kt[8]) );
  DFFHQX1 Kt_reg_4_ ( .D(N3137), .CK(clk), .Q(Kt[4]) );
  DFFHQX1 A_reg_18_ ( .D(n4746), .CK(clk), .Q(SHA256_result[242]) );
  DFFHQXL A_reg_19_ ( .D(n4745), .CK(clk), .Q(SHA256_result[243]) );
  DFFHQX1 A_reg_21_ ( .D(n4743), .CK(clk), .Q(SHA256_result[245]) );
  DFFHQXL A_reg_22_ ( .D(n4742), .CK(clk), .Q(SHA256_result[246]) );
  DFFHQXL A_reg_23_ ( .D(n4741), .CK(clk), .Q(SHA256_result[247]) );
  DFFHQXL A_reg_24_ ( .D(n4740), .CK(clk), .Q(SHA256_result[248]) );
  DFFHQXL A_reg_25_ ( .D(n4739), .CK(clk), .Q(SHA256_result[249]) );
  DFFHQXL A_reg_27_ ( .D(n4737), .CK(clk), .Q(SHA256_result[251]) );
  DFFHQXL A_reg_28_ ( .D(n4736), .CK(clk), .Q(SHA256_result[252]) );
  DFFHQXL E_reg_18_ ( .D(n4552), .CK(clk), .Q(SHA256_result[114]) );
  DFFTRX1 M_reg_21_ ( .D(M_w[21]), .RN(n401), .CK(clk), .Q(M[21]) );
  DFFTRX1 M_reg_20_ ( .D(M_w[20]), .RN(n401), .CK(clk), .Q(M[20]) );
  DFFTRX1 L_reg_18_ ( .D(n169), .RN(n403), .CK(clk), .Q(L[18]) );
  DFFTRX1 L_reg_15_ ( .D(T1_32[15]), .RN(n404), .CK(clk), .Q(L[15]) );
  DFFTRX1 M_reg_17_ ( .D(M_w[17]), .RN(n404), .CK(clk), .Q(M[17]) );
  DFFTRX1 L_reg_7_ ( .D(T1_32[7]), .RN(n404), .CK(clk), .Q(L[7]) );
  DFFHQX1 Kt_reg_7_ ( .D(N3140), .CK(clk), .Q(Kt[7]) );
  DFFHQX1 Kt_reg_6_ ( .D(N3139), .CK(clk), .Q(Kt[6]) );
  DFFHQX1 Kt_reg_5_ ( .D(N3138), .CK(clk), .Q(Kt[5]) );
  DFFHQX1 Kt_reg_3_ ( .D(N3136), .CK(clk), .Q(Kt[3]) );
  DFFHQX1 Kt_reg_2_ ( .D(N3135), .CK(clk), .Q(Kt[2]) );
  DFFHQX1 Kt_reg_0_ ( .D(N3133), .CK(clk), .Q(Kt[0]) );
  DFFTRX1 L_reg_6_ ( .D(T1_32[6]), .RN(n404), .CK(clk), .Q(L[6]) );
  DFFTRX1 output_valid_reg ( .D(output_enable), .RN(n3114), .CK(clk), .Q(
        output_valid) );
  DFFHQX1 digest_reg_3_ ( .D(N3578), .CK(clk), .Q(digest[3]) );
  DFFHQX1 digest_reg_2_ ( .D(N3577), .CK(clk), .Q(digest[2]) );
  DFFHQX1 digest_reg_1_ ( .D(N3576), .CK(clk), .Q(digest[1]) );
  DFFHQX1 digest_reg_0_ ( .D(N3575), .CK(clk), .Q(digest[0]) );
  DFFHQXL D_reg_11_ ( .D(n4623), .CK(clk), .Q(SHA256_result[139]) );
  DFFHQXL D_reg_2_ ( .D(n4632), .CK(clk), .Q(SHA256_result[130]) );
  DFFHQXL F_reg_24_ ( .D(n4419), .CK(clk), .Q(SHA256_result[88]) );
  DFFHQXL A_reg_20_ ( .D(n4744), .CK(clk), .Q(SHA256_result[244]) );
  DFFHQXL D_reg_0_ ( .D(n4634), .CK(clk), .Q(SHA256_result[128]) );
  DFFHQX4 mux_control_reg_0_ ( .D(n4700), .CK(clk), .Q(mux_control_0_) );
  DFFTRX1 round_reg_6_ ( .D(N158), .RN(n4250), .CK(clk), .Q(round[6]), .QN(
        n2878) );
  DFFHQX1 A_reg_16_ ( .D(n4748), .CK(clk), .Q(SHA256_result[240]) );
  DFFHQXL H2_reg_31_ ( .D(n4475), .CK(clk), .Q(H2[31]) );
  DFFHQXL H6_reg_31_ ( .D(n4348), .CK(clk), .Q(H6[31]) );
  DFFHQXL H4_reg_31_ ( .D(n4507), .CK(clk), .Q(H4[31]) );
  DFFHQXL H0_reg_31_ ( .D(n4702), .CK(clk), .Q(H0[31]) );
  DFFHQXL H5_reg_31_ ( .D(n4316), .CK(clk), .Q(H5[31]) );
  DFFHQXL H3_reg_31_ ( .D(n4571), .CK(clk), .Q(H3[31]) );
  DFFHQXL H7_reg_31_ ( .D(n4252), .CK(clk), .Q(H7[31]) );
  DFFHQXL H1_reg_31_ ( .D(n4444), .CK(clk), .Q(H1[31]) );
  DFFHQXL H1_reg_30_ ( .D(n4445), .CK(clk), .Q(H1[30]) );
  DFFHQXL H5_reg_30_ ( .D(n4317), .CK(clk), .Q(H5[30]) );
  DFFHQXL H5_reg_29_ ( .D(n4318), .CK(clk), .Q(H5[29]) );
  DFFHQXL H2_reg_30_ ( .D(n4476), .CK(clk), .Q(H2[30]) );
  DFFHQXL H6_reg_29_ ( .D(n4350), .CK(clk), .Q(H6[29]) );
  DFFHQXL H6_reg_30_ ( .D(n4349), .CK(clk), .Q(H6[30]) );
  DFFHQXL H3_reg_30_ ( .D(n4572), .CK(clk), .Q(H3[30]) );
  DFFHQXL H2_reg_29_ ( .D(n4477), .CK(clk), .Q(H2[29]) );
  DFFHQXL H3_reg_29_ ( .D(n4573), .CK(clk), .Q(H3[29]) );
  DFFHQXL H7_reg_30_ ( .D(n4253), .CK(clk), .Q(H7[30]) );
  DFFHQXL H0_reg_28_ ( .D(n4705), .CK(clk), .Q(H0[28]) );
  DFFHQXL H4_reg_29_ ( .D(n4509), .CK(clk), .Q(H4[29]) );
  DFFHQXL H_reg_29_ ( .D(n4285), .CK(clk), .Q(SHA256_result[29]) );
  DFFHQXL H_reg_31_ ( .D(n4283), .CK(clk), .Q(SHA256_result[31]) );
  DFFHQXL H_reg_28_ ( .D(n4286), .CK(clk), .Q(SHA256_result[28]) );
  DFFHQXL H_reg_30_ ( .D(n4284), .CK(clk), .Q(SHA256_result[30]) );
  DFFHQXL H4_reg_30_ ( .D(n4508), .CK(clk), .Q(H4[30]) );
  DFFHQXL H0_reg_29_ ( .D(n4704), .CK(clk), .Q(H0[29]) );
  DFFHQXL H4_reg_28_ ( .D(n4510), .CK(clk), .Q(H4[28]) );
  DFFHQXL H0_reg_30_ ( .D(n4703), .CK(clk), .Q(H0[30]) );
  DFFHQXL Kt_reg_28_ ( .D(N3161), .CK(clk), .Q(Kt[28]) );
  DFFHQXL H7_reg_29_ ( .D(n4254), .CK(clk), .Q(H7[29]) );
  DFFHQXL H3_reg_28_ ( .D(n4574), .CK(clk), .Q(H3[28]) );
  DFFHQXL H1_reg_28_ ( .D(n4447), .CK(clk), .Q(H1[28]) );
  DFFHQXL H1_reg_29_ ( .D(n4446), .CK(clk), .Q(H1[29]) );
  DFFHQXL H5_reg_28_ ( .D(n4319), .CK(clk), .Q(H5[28]) );
  DFFHQXL H6_reg_28_ ( .D(n4351), .CK(clk), .Q(H6[28]) );
  DFFHQXL H7_reg_28_ ( .D(n4255), .CK(clk), .Q(H7[28]) );
  DFFHQXL H0_reg_27_ ( .D(n4706), .CK(clk), .Q(H0[27]) );
  DFFHQXL H0_reg_21_ ( .D(n4712), .CK(clk), .Q(H0[21]) );
  DFFHQXL H2_reg_28_ ( .D(n4478), .CK(clk), .Q(H2[28]) );
  DFFHQXL H0_reg_23_ ( .D(n4710), .CK(clk), .Q(H0[23]) );
  DFFHQXL H4_reg_15_ ( .D(n4523), .CK(clk), .Q(H4[15]) );
  DFFHQXL H4_reg_14_ ( .D(n4524), .CK(clk), .Q(H4[14]) );
  DFFHQXL H4_reg_24_ ( .D(n4514), .CK(clk), .Q(H4[24]) );
  DFFHQXL H_reg_24_ ( .D(n4290), .CK(clk), .Q(SHA256_result[24]) );
  DFFHQXL H_reg_27_ ( .D(n4287), .CK(clk), .Q(SHA256_result[27]) );
  DFFHQXL H0_reg_22_ ( .D(n4711), .CK(clk), .Q(H0[22]) );
  DFFHQXL H4_reg_8_ ( .D(n4530), .CK(clk), .Q(H4[8]) );
  DFFHQXL H4_reg_23_ ( .D(n4515), .CK(clk), .Q(H4[23]) );
  DFFHQXL D_reg_30_ ( .D(n4604), .CK(clk), .Q(SHA256_result[158]) );
  DFFHQXL D_reg_31_ ( .D(n4603), .CK(clk), .Q(SHA256_result[159]) );
  DFFHQXL H4_reg_22_ ( .D(n4516), .CK(clk), .Q(H4[22]) );
  DFFHQXL H4_reg_27_ ( .D(n4511), .CK(clk), .Q(H4[27]) );
  DFFHQXL H0_reg_20_ ( .D(n4713), .CK(clk), .Q(H0[20]) );
  DFFHQXL H0_reg_24_ ( .D(n4709), .CK(clk), .Q(H0[24]) );
  DFFHQXL H4_reg_21_ ( .D(n4517), .CK(clk), .Q(H4[21]) );
  DFFHQXL H4_reg_13_ ( .D(n4525), .CK(clk), .Q(H4[13]) );
  DFFHQXL H4_reg_19_ ( .D(n4519), .CK(clk), .Q(H4[19]) );
  DFFHQXL H4_reg_16_ ( .D(n4522), .CK(clk), .Q(H4[16]) );
  DFFHQXL H0_reg_26_ ( .D(n4707), .CK(clk), .Q(H0[26]) );
  DFFHQXL H0_reg_25_ ( .D(n4708), .CK(clk), .Q(H0[25]) );
  DFFHQXL H4_reg_20_ ( .D(n4518), .CK(clk), .Q(H4[20]) );
  DFFHQXL H4_reg_26_ ( .D(n4512), .CK(clk), .Q(H4[26]) );
  DFFHQXL H4_reg_25_ ( .D(n4513), .CK(clk), .Q(H4[25]) );
  DFFHQXL H2_reg_24_ ( .D(n4482), .CK(clk), .Q(H2[24]) );
  DFFHQXL H5_reg_26_ ( .D(n4321), .CK(clk), .Q(H5[26]) );
  DFFHQXL H3_reg_27_ ( .D(n4575), .CK(clk), .Q(H3[27]) );
  DFFHQXL H2_reg_26_ ( .D(n4480), .CK(clk), .Q(H2[26]) );
  DFFHQXL H6_reg_26_ ( .D(n4353), .CK(clk), .Q(H6[26]) );
  DFFHQXL H1_reg_24_ ( .D(n4451), .CK(clk), .Q(H1[24]) );
  DFFHQXL H3_reg_24_ ( .D(n4578), .CK(clk), .Q(H3[24]) );
  DFFHQXL H3_reg_26_ ( .D(n4576), .CK(clk), .Q(H3[26]) );
  DFFHQXL H5_reg_24_ ( .D(n4323), .CK(clk), .Q(H5[24]) );
  DFFHQXL H5_reg_25_ ( .D(n4322), .CK(clk), .Q(H5[25]) );
  DFFHQXL H6_reg_24_ ( .D(n4355), .CK(clk), .Q(H6[24]) );
  DFFHQXL H1_reg_27_ ( .D(n4448), .CK(clk), .Q(H1[27]) );
  DFFHQXL H2_reg_27_ ( .D(n4479), .CK(clk), .Q(H2[27]) );
  DFFHQXL H5_reg_27_ ( .D(n4320), .CK(clk), .Q(H5[27]) );
  DFFHQXL H6_reg_27_ ( .D(n4352), .CK(clk), .Q(H6[27]) );
  DFFHQXL H7_reg_27_ ( .D(n4256), .CK(clk), .Q(H7[27]) );
  DFFHQXL H4_reg_3_ ( .D(n4535), .CK(clk), .Q(H4[3]) );
  DFFHQXL H0_reg_17_ ( .D(n4716), .CK(clk), .Q(H0[17]) );
  DFFHQXL H0_reg_18_ ( .D(n4715), .CK(clk), .Q(H0[18]) );
  DFFHQXL H_reg_20_ ( .D(n4294), .CK(clk), .Q(SHA256_result[20]) );
  DFFHQXL H0_reg_15_ ( .D(n4718), .CK(clk), .Q(H0[15]) );
  DFFHQXL H0_reg_19_ ( .D(n4714), .CK(clk), .Q(H0[19]) );
  DFFHQXL H4_reg_9_ ( .D(n4529), .CK(clk), .Q(H4[9]) );
  DFFHQXL H_reg_26_ ( .D(n4288), .CK(clk), .Q(SHA256_result[26]) );
  DFFHQXL H_reg_21_ ( .D(n4293), .CK(clk), .Q(SHA256_result[21]) );
  DFFHQXL H_reg_22_ ( .D(n4292), .CK(clk), .Q(SHA256_result[22]) );
  DFFHQXL H_reg_23_ ( .D(n4291), .CK(clk), .Q(SHA256_result[23]) );
  DFFHQXL H_reg_25_ ( .D(n4289), .CK(clk), .Q(SHA256_result[25]) );
  DFFHQXL H4_reg_10_ ( .D(n4528), .CK(clk), .Q(H4[10]) );
  DFFHQXL H0_reg_14_ ( .D(n4719), .CK(clk), .Q(H0[14]) );
  DFFHQXL H4_reg_2_ ( .D(n4536), .CK(clk), .Q(H4[2]) );
  DFFHQXL H4_reg_0_ ( .D(n4538), .CK(clk), .Q(H4[0]) );
  DFFHQXL D_reg_28_ ( .D(n4606), .CK(clk), .Q(SHA256_result[156]) );
  DFFHQXL D_reg_27_ ( .D(n4607), .CK(clk), .Q(SHA256_result[155]) );
  DFFHQXL D_reg_29_ ( .D(n4605), .CK(clk), .Q(SHA256_result[157]) );
  DFFHQXL D_reg_26_ ( .D(n4608), .CK(clk), .Q(SHA256_result[154]) );
  DFFHQXL H0_reg_11_ ( .D(n4722), .CK(clk), .Q(H0[11]) );
  DFFHQXL H0_reg_9_ ( .D(n4724), .CK(clk), .Q(H0[9]) );
  DFFHQXL H0_reg_10_ ( .D(n4723), .CK(clk), .Q(H0[10]) );
  DFFHQXL H4_reg_17_ ( .D(n4521), .CK(clk), .Q(H4[17]) );
  DFFHQXL H4_reg_4_ ( .D(n4534), .CK(clk), .Q(H4[4]) );
  DFFHQXL H0_reg_12_ ( .D(n4721), .CK(clk), .Q(H0[12]) );
  DFFHQXL H0_reg_8_ ( .D(n4725), .CK(clk), .Q(H0[8]) );
  DFFHQXL H4_reg_7_ ( .D(n4531), .CK(clk), .Q(H4[7]) );
  DFFHQXL H4_reg_5_ ( .D(n4533), .CK(clk), .Q(H4[5]) );
  DFFHQXL H4_reg_6_ ( .D(n4532), .CK(clk), .Q(H4[6]) );
  DFFHQXL H0_reg_16_ ( .D(n4717), .CK(clk), .Q(H0[16]) );
  DFFHQXL H0_reg_13_ ( .D(n4720), .CK(clk), .Q(H0[13]) );
  DFFHQXL F_reg_31_ ( .D(n4412), .CK(clk), .Q(SHA256_result[95]) );
  DFFHQXL H4_reg_12_ ( .D(n4526), .CK(clk), .Q(H4[12]) );
  DFFHQXL H4_reg_18_ ( .D(n4520), .CK(clk), .Q(H4[18]) );
  DFFHQXL H4_reg_11_ ( .D(n4527), .CK(clk), .Q(H4[11]) );
  DFFHQXL C_reg_31_ ( .D(n4635), .CK(clk), .Q(SHA256_result[191]) );
  DFFHQXL G_reg_31_ ( .D(n4380), .CK(clk), .Q(SHA256_result[63]) );
  DFFHQXL B_reg_31_ ( .D(n4667), .CK(clk), .Q(SHA256_result[223]) );
  DFFHQXL Kt_reg_25_ ( .D(N3158), .CK(clk), .Q(Kt[25]) );
  DFFHQXL H1_reg_20_ ( .D(n4455), .CK(clk), .Q(H1[20]) );
  DFFHQXL H1_reg_26_ ( .D(n4449), .CK(clk), .Q(H1[26]) );
  DFFHQXL H2_reg_20_ ( .D(n4486), .CK(clk), .Q(H2[20]) );
  DFFHQXL H2_reg_25_ ( .D(n4481), .CK(clk), .Q(H2[25]) );
  DFFHQXL H5_reg_20_ ( .D(n4327), .CK(clk), .Q(H5[20]) );
  DFFHQXL H5_reg_21_ ( .D(n4326), .CK(clk), .Q(H5[21]) );
  DFFHQXL H5_reg_22_ ( .D(n4325), .CK(clk), .Q(H5[22]) );
  DFFHQXL H6_reg_20_ ( .D(n4359), .CK(clk), .Q(H6[20]) );
  DFFHQXL H6_reg_21_ ( .D(n4358), .CK(clk), .Q(H6[21]) );
  DFFHQXL H6_reg_22_ ( .D(n4357), .CK(clk), .Q(H6[22]) );
  DFFHQXL H7_reg_26_ ( .D(n4257), .CK(clk), .Q(H7[26]) );
  DFFHQXL H3_reg_20_ ( .D(n4582), .CK(clk), .Q(H3[20]) );
  DFFHQXL H3_reg_21_ ( .D(n4581), .CK(clk), .Q(H3[21]) );
  DFFHQXL H3_reg_25_ ( .D(n4577), .CK(clk), .Q(H3[25]) );
  DFFHQXL H1_reg_19_ ( .D(n4456), .CK(clk), .Q(H1[19]) );
  DFFHQXL H1_reg_23_ ( .D(n4452), .CK(clk), .Q(H1[23]) );
  DFFHQXL H2_reg_23_ ( .D(n4483), .CK(clk), .Q(H2[23]) );
  DFFHQXL H5_reg_19_ ( .D(n4328), .CK(clk), .Q(H5[19]) );
  DFFHQXL H6_reg_19_ ( .D(n4360), .CK(clk), .Q(H6[19]) );
  DFFHQXL H5_reg_23_ ( .D(n4324), .CK(clk), .Q(H5[23]) );
  DFFHQXL H3_reg_23_ ( .D(n4579), .CK(clk), .Q(H3[23]) );
  DFFHQXL H1_reg_22_ ( .D(n4453), .CK(clk), .Q(H1[22]) );
  DFFHQXL H2_reg_21_ ( .D(n4485), .CK(clk), .Q(H2[21]) );
  DFFHQXL H2_reg_22_ ( .D(n4484), .CK(clk), .Q(H2[22]) );
  DFFHQXL H1_reg_25_ ( .D(n4450), .CK(clk), .Q(H1[25]) );
  DFFHQXL H3_reg_22_ ( .D(n4580), .CK(clk), .Q(H3[22]) );
  DFFHQXL H6_reg_25_ ( .D(n4354), .CK(clk), .Q(H6[25]) );
  DFFHQXL H7_reg_24_ ( .D(n4259), .CK(clk), .Q(H7[24]) );
  DFFHQXL H7_reg_25_ ( .D(n4258), .CK(clk), .Q(H7[25]) );
  DFFHQXL H2_reg_19_ ( .D(n4487), .CK(clk), .Q(H2[19]) );
  DFFHQXL H3_reg_19_ ( .D(n4583), .CK(clk), .Q(H3[19]) );
  DFFHQXL H6_reg_23_ ( .D(n4356), .CK(clk), .Q(H6[23]) );
  DFFHQXL H7_reg_23_ ( .D(n4260), .CK(clk), .Q(H7[23]) );
  DFFHQXL H4_reg_1_ ( .D(n4537), .CK(clk), .Q(H4[1]) );
  DFFHQXL H0_reg_6_ ( .D(n4727), .CK(clk), .Q(H0[6]) );
  DFFHQXL H_reg_15_ ( .D(n4299), .CK(clk), .Q(SHA256_result[15]) );
  DFFHQXL H_reg_14_ ( .D(n4300), .CK(clk), .Q(SHA256_result[14]) );
  DFFHQXL H_reg_12_ ( .D(n4302), .CK(clk), .Q(SHA256_result[12]) );
  DFFHQXL H_reg_13_ ( .D(n4301), .CK(clk), .Q(SHA256_result[13]) );
  DFFHQXL H_reg_16_ ( .D(n4298), .CK(clk), .Q(SHA256_result[16]) );
  DFFHQXL H_reg_17_ ( .D(n4297), .CK(clk), .Q(SHA256_result[17]) );
  DFFHQXL H_reg_18_ ( .D(n4296), .CK(clk), .Q(SHA256_result[18]) );
  DFFHQXL H_reg_19_ ( .D(n4295), .CK(clk), .Q(SHA256_result[19]) );
  DFFHQXL D_reg_20_ ( .D(n4614), .CK(clk), .Q(SHA256_result[148]) );
  DFFHQXL D_reg_21_ ( .D(n4613), .CK(clk), .Q(SHA256_result[149]) );
  DFFHQXL D_reg_23_ ( .D(n4611), .CK(clk), .Q(SHA256_result[151]) );
  DFFHQXL D_reg_25_ ( .D(n4609), .CK(clk), .Q(SHA256_result[153]) );
  DFFHQXL D_reg_22_ ( .D(n4612), .CK(clk), .Q(SHA256_result[150]) );
  DFFHQXL D_reg_24_ ( .D(n4610), .CK(clk), .Q(SHA256_result[152]) );
  DFFHQXL H0_reg_7_ ( .D(n4726), .CK(clk), .Q(H0[7]) );
  DFFHQXL H0_reg_4_ ( .D(n4729), .CK(clk), .Q(H0[4]) );
  DFFHQXL H0_reg_5_ ( .D(n4728), .CK(clk), .Q(H0[5]) );
  DFFHQXL F_reg_30_ ( .D(n4413), .CK(clk), .Q(SHA256_result[94]) );
  DFFHQXL B_reg_30_ ( .D(n4668), .CK(clk), .Q(SHA256_result[222]) );
  DFFHQXL C_reg_30_ ( .D(n4636), .CK(clk), .Q(SHA256_result[190]) );
  DFFHQXL G_reg_30_ ( .D(n4381), .CK(clk), .Q(SHA256_result[62]) );
  DFFHQXL D_reg_9_ ( .D(n4625), .CK(clk), .Q(SHA256_result[137]) );
  DFFHQXL H_reg_2_ ( .D(n4312), .CK(clk), .Q(SHA256_result[2]) );
  DFFHQXL H_reg_3_ ( .D(n4311), .CK(clk), .Q(SHA256_result[3]) );
  DFFHQXL H2_reg_16_ ( .D(n4490), .CK(clk), .Q(H2[16]) );
  DFFHQXL H6_reg_18_ ( .D(n4361), .CK(clk), .Q(H6[18]) );
  DFFHQXL H5_reg_17_ ( .D(n4330), .CK(clk), .Q(H5[17]) );
  DFFHQXL H7_reg_20_ ( .D(n4263), .CK(clk), .Q(H7[20]) );
  DFFHQXL H7_reg_16_ ( .D(n4267), .CK(clk), .Q(H7[16]) );
  DFFHQXL H7_reg_18_ ( .D(n4265), .CK(clk), .Q(H7[18]) );
  DFFHQXL H7_reg_17_ ( .D(n4266), .CK(clk), .Q(H7[17]) );
  DFFHQXL H7_reg_19_ ( .D(n4264), .CK(clk), .Q(H7[19]) );
  DFFHQXL H5_reg_0_ ( .D(n4347), .CK(clk), .Q(H5[0]) );
  DFFHQXL H1_reg_17_ ( .D(n4458), .CK(clk), .Q(H1[17]) );
  DFFHQXL H1_reg_18_ ( .D(n4457), .CK(clk), .Q(H1[18]) );
  DFFHQXL H1_reg_21_ ( .D(n4454), .CK(clk), .Q(H1[21]) );
  DFFHQXL H2_reg_17_ ( .D(n4489), .CK(clk), .Q(H2[17]) );
  DFFHQXL H2_reg_18_ ( .D(n4488), .CK(clk), .Q(H2[18]) );
  DFFHQXL H5_reg_18_ ( .D(n4329), .CK(clk), .Q(H5[18]) );
  DFFHQXL H6_reg_16_ ( .D(n4363), .CK(clk), .Q(H6[16]) );
  DFFHQXL H6_reg_17_ ( .D(n4362), .CK(clk), .Q(H6[17]) );
  DFFHQXL H1_reg_16_ ( .D(n4459), .CK(clk), .Q(H1[16]) );
  DFFHQXL H3_reg_16_ ( .D(n4586), .CK(clk), .Q(H3[16]) );
  DFFHQXL H3_reg_17_ ( .D(n4585), .CK(clk), .Q(H3[17]) );
  DFFHQXL H3_reg_18_ ( .D(n4584), .CK(clk), .Q(H3[18]) );
  DFFHQXL H5_reg_16_ ( .D(n4331), .CK(clk), .Q(H5[16]) );
  DFFHQXL H7_reg_21_ ( .D(n4262), .CK(clk), .Q(H7[21]) );
  DFFHQXL H7_reg_22_ ( .D(n4261), .CK(clk), .Q(H7[22]) );
  DFFHQXL H0_reg_0_ ( .D(n4765), .CK(clk), .Q(H0[0]) );
  DFFHQXL H0_reg_1_ ( .D(n4732), .CK(clk), .Q(H0[1]) );
  DFFHQXL H_reg_7_ ( .D(n4307), .CK(clk), .Q(SHA256_result[7]) );
  DFFHQXL H_reg_9_ ( .D(n4305), .CK(clk), .Q(SHA256_result[9]) );
  DFFHQXL D_reg_13_ ( .D(n4621), .CK(clk), .Q(SHA256_result[141]) );
  DFFHQXL H_reg_11_ ( .D(n4303), .CK(clk), .Q(SHA256_result[11]) );
  DFFHQXL H_reg_10_ ( .D(n4304), .CK(clk), .Q(SHA256_result[10]) );
  DFFHQXL H_reg_8_ ( .D(n4306), .CK(clk), .Q(SHA256_result[8]) );
  DFFHQXL D_reg_14_ ( .D(n4620), .CK(clk), .Q(SHA256_result[142]) );
  DFFHQXL D_reg_15_ ( .D(n4619), .CK(clk), .Q(SHA256_result[143]) );
  DFFHQXL D_reg_12_ ( .D(n4622), .CK(clk), .Q(SHA256_result[140]) );
  DFFHQXL H0_reg_2_ ( .D(n4731), .CK(clk), .Q(H0[2]) );
  DFFHQXL D_reg_16_ ( .D(n4618), .CK(clk), .Q(SHA256_result[144]) );
  DFFHQXL D_reg_17_ ( .D(n4617), .CK(clk), .Q(SHA256_result[145]) );
  DFFHQXL D_reg_19_ ( .D(n4615), .CK(clk), .Q(SHA256_result[147]) );
  DFFHQXL D_reg_18_ ( .D(n4616), .CK(clk), .Q(SHA256_result[146]) );
  DFFHQXL F_reg_29_ ( .D(n4414), .CK(clk), .Q(SHA256_result[93]) );
  DFFHQXL B_reg_28_ ( .D(n4670), .CK(clk), .Q(SHA256_result[220]) );
  DFFHQXL B_reg_29_ ( .D(n4669), .CK(clk), .Q(SHA256_result[221]) );
  DFFHQXL C_reg_29_ ( .D(n4637), .CK(clk), .Q(SHA256_result[189]) );
  DFFHQXL C_reg_28_ ( .D(n4638), .CK(clk), .Q(SHA256_result[188]) );
  DFFHQX1 H_reg_6_ ( .D(n4308), .CK(clk), .Q(SHA256_result[6]) );
  DFFHQX1 H7_reg_6_ ( .D(n4277), .CK(clk), .Q(H7[6]) );
  DFFHQX1 H7_reg_2_ ( .D(n4281), .CK(clk), .Q(H7[2]) );
  DFFHQX1 H7_reg_5_ ( .D(n4278), .CK(clk), .Q(H7[5]) );
  DFFHQX1 C_reg_24_ ( .D(n4642), .CK(clk), .Q(SHA256_result[184]) );
  DFFHQX1 B_reg_24_ ( .D(n4674), .CK(clk), .Q(SHA256_result[216]) );
  DFFHQX1 G_reg_27_ ( .D(n4384), .CK(clk), .Q(SHA256_result[59]) );
  DFFHQX1 F_reg_25_ ( .D(n4418), .CK(clk), .Q(SHA256_result[89]) );
  DFFTRXL M_reg_29_ ( .D(M_w[29]), .RN(n401), .CK(clk), .Q(M[29]) );
  DFFTRXL M_reg_28_ ( .D(M_w[28]), .RN(n401), .CK(clk), .Q(M[28]) );
  DFFTRXL M_reg_30_ ( .D(M_w[30]), .RN(n401), .CK(clk), .Q(M[30]) );
  DFFTRXL M_reg_24_ ( .D(M_w[24]), .RN(n401), .CK(clk), .Q(M[24]) );
  DFFTRXL M_reg_27_ ( .D(M_w[27]), .RN(n401), .CK(clk), .Q(M[27]) );
  DFFHQXL H5_reg_15_ ( .D(n4332), .CK(clk), .Q(H5[15]) );
  DFFHQXL H3_reg_0_ ( .D(n4602), .CK(clk), .Q(H3[0]) );
  DFFHQXL H5_reg_3_ ( .D(n4344), .CK(clk), .Q(H5[3]) );
  DFFHQXL H5_reg_2_ ( .D(n4345), .CK(clk), .Q(H5[2]) );
  DFFHQXL H2_reg_0_ ( .D(n4506), .CK(clk), .Q(H2[0]) );
  DFFHQXL H3_reg_3_ ( .D(n4599), .CK(clk), .Q(H3[3]) );
  DFFHQXL H2_reg_3_ ( .D(n4503), .CK(clk), .Q(H2[3]) );
  DFFHQXL H3_reg_2_ ( .D(n4600), .CK(clk), .Q(H3[2]) );
  DFFHQXL H6_reg_0_ ( .D(n4379), .CK(clk), .Q(H6[0]) );
  DFFHQXL H2_reg_2_ ( .D(n4504), .CK(clk), .Q(H2[2]) );
  DFFHQXL H5_reg_11_ ( .D(n4336), .CK(clk), .Q(H5[11]) );
  DFFHQXL G_reg_29_ ( .D(n4382), .CK(clk), .Q(SHA256_result[61]) );
  DFFHQX1 H7_reg_14_ ( .D(n4269), .CK(clk), .Q(H7[14]) );
  DFFHQX1 H7_reg_8_ ( .D(n4275), .CK(clk), .Q(H7[8]) );
  DFFHQX1 H7_reg_10_ ( .D(n4273), .CK(clk), .Q(H7[10]) );
  DFFHQX1 H7_reg_11_ ( .D(n4272), .CK(clk), .Q(H7[11]) );
  DFFHQX1 H7_reg_15_ ( .D(n4268), .CK(clk), .Q(H7[15]) );
  DFFHQX1 D_reg_1_ ( .D(n4633), .CK(clk), .Q(SHA256_result[129]) );
  DFFX4 F_reg_0_ ( .D(n4443), .CK(clk), .Q(n238), .QN(n237) );
  DFFTRXL M_reg_31_ ( .D(M_w[31]), .RN(n401), .CK(clk), .Q(M[31]) );
  DFFHQXL D_reg_7_ ( .D(n4627), .CK(clk), .Q(SHA256_result[135]) );
  DFFHQXL D_reg_6_ ( .D(n4628), .CK(clk), .Q(SHA256_result[134]) );
  DFFHQXL H_reg_5_ ( .D(n4309), .CK(clk), .Q(SHA256_result[5]) );
  DFFHQXL H_reg_4_ ( .D(n4310), .CK(clk), .Q(SHA256_result[4]) );
  DFFHQXL D_reg_10_ ( .D(n4624), .CK(clk), .Q(SHA256_result[138]) );
  DFFHQXL D_reg_8_ ( .D(n4626), .CK(clk), .Q(SHA256_result[136]) );
  DFFHQX1 F_reg_26_ ( .D(n4417), .CK(clk), .Q(SHA256_result[90]) );
  DFFX4 G_reg_0_ ( .D(n4411), .CK(clk), .Q(n231), .QN(n230) );
  DFFHQX1 G_reg_26_ ( .D(n4385), .CK(clk), .Q(SHA256_result[58]) );
  DFFTRXL M_reg_26_ ( .D(M_w[26]), .RN(n401), .CK(clk), .Q(M[26]) );
  DFFTRXL M_reg_25_ ( .D(M_w[25]), .RN(n401), .CK(clk), .Q(M[25]) );
  DFFHQXL F_reg_28_ ( .D(n4415), .CK(clk), .Q(SHA256_result[92]) );
  DFFHQXL G_reg_28_ ( .D(n4383), .CK(clk), .Q(SHA256_result[60]) );
  DFFHQX1 D_reg_4_ ( .D(n4630), .CK(clk), .Q(SHA256_result[132]) );
  DFFHQX1 D_reg_5_ ( .D(n4629), .CK(clk), .Q(SHA256_result[133]) );
  DFFHQX1 D_reg_3_ ( .D(n4631), .CK(clk), .Q(SHA256_result[131]) );
  DFFHQX1 H_reg_1_ ( .D(n4313), .CK(clk), .Q(SHA256_result[1]) );
  DFFHQX1 H_reg_0_ ( .D(n4314), .CK(clk), .Q(SHA256_result[0]) );
  DFFHQX1 H1_reg_8_ ( .D(n4467), .CK(clk), .Q(H1[8]) );
  DFFHQX1 H1_reg_12_ ( .D(n4463), .CK(clk), .Q(H1[12]) );
  DFFHQX1 H7_reg_7_ ( .D(n4276), .CK(clk), .Q(H7[7]) );
  DFFHQX1 H7_reg_9_ ( .D(n4274), .CK(clk), .Q(H7[9]) );
  DFFHQX1 H7_reg_12_ ( .D(n4271), .CK(clk), .Q(H7[12]) );
  DFFHQX1 H7_reg_13_ ( .D(n4270), .CK(clk), .Q(H7[13]) );
  DFFHQX1 H2_reg_1_ ( .D(n4505), .CK(clk), .Q(H2[1]) );
  DFFHQX1 H2_reg_4_ ( .D(n4502), .CK(clk), .Q(H2[4]) );
  DFFHQX1 H2_reg_6_ ( .D(n4500), .CK(clk), .Q(H2[6]) );
  DFFHQX1 H2_reg_14_ ( .D(n4492), .CK(clk), .Q(H2[14]) );
  DFFHQX1 H3_reg_1_ ( .D(n4601), .CK(clk), .Q(H3[1]) );
  DFFHQX1 H3_reg_4_ ( .D(n4598), .CK(clk), .Q(H3[4]) );
  DFFHQX1 H3_reg_6_ ( .D(n4596), .CK(clk), .Q(H3[6]) );
  DFFHQX1 H3_reg_14_ ( .D(n4588), .CK(clk), .Q(H3[14]) );
  DFFHQX1 H5_reg_4_ ( .D(n4343), .CK(clk), .Q(H5[4]) );
  DFFHQX1 H5_reg_6_ ( .D(n4341), .CK(clk), .Q(H5[6]) );
  DFFHQX1 H5_reg_14_ ( .D(n4333), .CK(clk), .Q(H5[14]) );
  DFFHQX1 H6_reg_4_ ( .D(n4375), .CK(clk), .Q(H6[4]) );
  DFFHQX1 H6_reg_6_ ( .D(n4373), .CK(clk), .Q(H6[6]) );
  DFFHQX1 H6_reg_14_ ( .D(n4365), .CK(clk), .Q(H6[14]) );
  DFFHQX1 H7_reg_1_ ( .D(n4282), .CK(clk), .Q(H7[1]) );
  DFFHQX1 H7_reg_4_ ( .D(n4279), .CK(clk), .Q(H7[4]) );
  DFFHQX1 H1_reg_0_ ( .D(n4699), .CK(clk), .Q(H1[0]) );
  DFFHQX1 H1_reg_2_ ( .D(n4473), .CK(clk), .Q(H1[2]) );
  DFFHQX1 H1_reg_7_ ( .D(n4468), .CK(clk), .Q(H1[7]) );
  DFFHQX1 H1_reg_9_ ( .D(n4466), .CK(clk), .Q(H1[9]) );
  DFFHQX1 H1_reg_10_ ( .D(n4465), .CK(clk), .Q(H1[10]) );
  DFFHQX1 H1_reg_11_ ( .D(n4464), .CK(clk), .Q(H1[11]) );
  DFFHQX1 H1_reg_13_ ( .D(n4462), .CK(clk), .Q(H1[13]) );
  DFFHQX1 H1_reg_15_ ( .D(n4460), .CK(clk), .Q(H1[15]) );
  DFFHQX1 H2_reg_5_ ( .D(n4501), .CK(clk), .Q(H2[5]) );
  DFFHQX1 H2_reg_7_ ( .D(n4499), .CK(clk), .Q(H2[7]) );
  DFFHQX1 H2_reg_8_ ( .D(n4498), .CK(clk), .Q(H2[8]) );
  DFFHQX1 H2_reg_9_ ( .D(n4497), .CK(clk), .Q(H2[9]) );
  DFFHQX1 H2_reg_10_ ( .D(n4496), .CK(clk), .Q(H2[10]) );
  DFFHQX1 H2_reg_11_ ( .D(n4495), .CK(clk), .Q(H2[11]) );
  DFFHQX1 H2_reg_12_ ( .D(n4494), .CK(clk), .Q(H2[12]) );
  DFFHQX1 H2_reg_13_ ( .D(n4493), .CK(clk), .Q(H2[13]) );
  DFFHQX1 H2_reg_15_ ( .D(n4491), .CK(clk), .Q(H2[15]) );
  DFFHQX1 H3_reg_5_ ( .D(n4597), .CK(clk), .Q(H3[5]) );
  DFFHQX1 H3_reg_7_ ( .D(n4595), .CK(clk), .Q(H3[7]) );
  DFFHQX1 H3_reg_8_ ( .D(n4594), .CK(clk), .Q(H3[8]) );
  DFFHQX1 H3_reg_9_ ( .D(n4593), .CK(clk), .Q(H3[9]) );
  DFFHQX1 H3_reg_10_ ( .D(n4592), .CK(clk), .Q(H3[10]) );
  DFFHQX1 H3_reg_12_ ( .D(n4590), .CK(clk), .Q(H3[12]) );
  DFFHQX1 H3_reg_13_ ( .D(n4589), .CK(clk), .Q(H3[13]) );
  DFFHQX1 H3_reg_15_ ( .D(n4587), .CK(clk), .Q(H3[15]) );
  DFFHQX1 H5_reg_5_ ( .D(n4342), .CK(clk), .Q(H5[5]) );
  DFFHQX1 H5_reg_8_ ( .D(n4339), .CK(clk), .Q(H5[8]) );
  DFFHQX1 H5_reg_9_ ( .D(n4338), .CK(clk), .Q(H5[9]) );
  DFFHQX1 H5_reg_10_ ( .D(n4337), .CK(clk), .Q(H5[10]) );
  DFFHQX1 H5_reg_12_ ( .D(n4335), .CK(clk), .Q(H5[12]) );
  DFFHQX1 H5_reg_13_ ( .D(n4334), .CK(clk), .Q(H5[13]) );
  DFFHQX1 H6_reg_2_ ( .D(n4377), .CK(clk), .Q(H6[2]) );
  DFFHQX1 H6_reg_3_ ( .D(n4376), .CK(clk), .Q(H6[3]) );
  DFFHQX1 H6_reg_5_ ( .D(n4374), .CK(clk), .Q(H6[5]) );
  DFFHQX1 H6_reg_7_ ( .D(n4372), .CK(clk), .Q(H6[7]) );
  DFFHQX1 H6_reg_8_ ( .D(n4371), .CK(clk), .Q(H6[8]) );
  DFFHQX1 H6_reg_9_ ( .D(n4370), .CK(clk), .Q(H6[9]) );
  DFFHQX1 H6_reg_10_ ( .D(n4369), .CK(clk), .Q(H6[10]) );
  DFFHQX1 H6_reg_11_ ( .D(n4368), .CK(clk), .Q(H6[11]) );
  DFFHQX1 H6_reg_12_ ( .D(n4367), .CK(clk), .Q(H6[12]) );
  DFFHQX1 H6_reg_13_ ( .D(n4366), .CK(clk), .Q(H6[13]) );
  DFFHQX1 H6_reg_15_ ( .D(n4364), .CK(clk), .Q(H6[15]) );
  DFFHQX1 H7_reg_0_ ( .D(n4315), .CK(clk), .Q(H7[0]) );
  DFFHQX1 H7_reg_3_ ( .D(n4280), .CK(clk), .Q(H7[3]) );
  DFFHQX1 B_reg_26_ ( .D(n4672), .CK(clk), .Q(SHA256_result[218]) );
  DFFHQX1 B_reg_27_ ( .D(n4671), .CK(clk), .Q(SHA256_result[219]) );
  DFFHQX1 C_reg_26_ ( .D(n4640), .CK(clk), .Q(SHA256_result[186]) );
  DFFHQX1 F_reg_27_ ( .D(n4416), .CK(clk), .Q(SHA256_result[91]) );
  DFFHQX1 C_reg_27_ ( .D(n4639), .CK(clk), .Q(SHA256_result[187]) );
  DFFTRX1 round_reg_1_ ( .D(N153), .RN(n4250), .CK(clk), .Q(round[1]), .QN(
        n2946) );
  DFFTRX1 round_reg_2_ ( .D(N154), .RN(n4250), .CK(clk), .Q(round[2]), .QN(
        n2943) );
  DFFTRX1 round_reg_0_ ( .D(N152), .RN(n4250), .CK(clk), .Q(round[0]), .QN(
        n2947) );
  DFFTRX1 M_reg_23_ ( .D(M_w[23]), .RN(n401), .CK(clk), .Q(M[23]) );
  DFFTRX1 M_reg_22_ ( .D(M_w[22]), .RN(n401), .CK(clk), .Q(M[22]) );
  DFFTRX1 M_reg_16_ ( .D(M_w[16]), .RN(n403), .CK(clk), .Q(M[16]) );
  DFFX4 A_reg_3_ ( .D(n4761), .CK(clk), .Q(n221), .QN(n220) );
  DFFTRX2 L_reg_5_ ( .D(T1_32[5]), .RN(n404), .CK(clk), .Q(L[5]) );
  DFFTRX2 L_reg_1_ ( .D(T1_32[1]), .RN(n403), .CK(clk), .Q(L[1]) );
  DFFX4 F_reg_2_ ( .D(n4441), .CK(clk), .Q(n212), .QN(n211) );
  DFFHQXL H1_reg_1_ ( .D(n4474), .CK(clk), .Q(H1[1]) );
  DFFHQXL H1_reg_4_ ( .D(n4471), .CK(clk), .Q(H1[4]) );
  DFFHQXL H1_reg_6_ ( .D(n4469), .CK(clk), .Q(H1[6]) );
  DFFHQXL H1_reg_3_ ( .D(n4472), .CK(clk), .Q(H1[3]) );
  DFFHQXL H1_reg_5_ ( .D(n4470), .CK(clk), .Q(H1[5]) );
  DFFHQXL H3_reg_11_ ( .D(n4591), .CK(clk), .Q(H3[11]) );
  DFFX4 G_reg_5_ ( .D(n4406), .CK(clk), .Q(n173), .QN(n172) );
  DFFX4 F_reg_7_ ( .D(n4436), .CK(clk), .Q(n167), .QN(n168) );
  DFFX4 G_reg_9_ ( .D(n4402), .CK(clk), .Q(n165), .QN(n166) );
  DFFX4 G_reg_1_ ( .D(n4410), .CK(clk), .Q(n163), .QN(n162) );
  DFFX4 G_reg_10_ ( .D(n4401), .CK(clk), .Q(n159), .QN(n160) );
  DFFX4 E_reg_1_ ( .D(n4569), .CK(clk), .Q(n157), .QN(n156) );
  DFFX4 E_reg_7_ ( .D(n4563), .CK(clk), .Q(n153), .QN(n152) );
  DFFHQX4 G_reg_2_ ( .D(n4409), .CK(clk), .Q(n151) );
  DFFX4 E_reg_5_ ( .D(n4565), .CK(clk), .Q(n149), .QN(n148) );
  DFFX4 G_reg_7_ ( .D(n4404), .CK(clk), .Q(n133), .QN(n132) );
  DFFX4 F_reg_5_ ( .D(n4438), .CK(clk), .Q(n129), .QN(n128) );
  DFFX4 E_reg_10_ ( .D(n4560), .CK(clk), .Q(n126), .QN(n125) );
  DFFXL E_reg_27_ ( .D(n4543), .CK(clk), .Q(n122), .QN(n121) );
  DFFX1 G_reg_24_ ( .D(n4387), .CK(clk), .Q(n119), .QN(n120) );
  DFFXL E_reg_26_ ( .D(n4544), .CK(clk), .Q(n117), .QN(n116) );
  DFFXL E_reg_30_ ( .D(n4540), .CK(clk), .Q(n114), .QN(n113) );
  DFFX4 E_reg_19_ ( .D(n4551), .CK(clk), .Q(n111), .QN(n112) );
  DFFXL E_reg_29_ ( .D(n4541), .CK(clk), .Q(n109), .QN(n108) );
  DFFXL E_reg_31_ ( .D(n4539), .CK(clk), .Q(n105), .QN(n104) );
  DFFXL E_reg_24_ ( .D(n4546), .CK(clk), .Q(n102), .QN(n101) );
  DFFX4 B_reg_3_ ( .D(n4695), .CK(clk), .Q(n99), .QN(n98) );
  DFFX4 B_reg_0_ ( .D(n4698), .CK(clk), .Q(n96), .QN(n97) );
  DFFXL E_reg_28_ ( .D(n4542), .CK(clk), .Q(n93), .QN(n92) );
  DFFX4 E_reg_23_ ( .D(n4547), .CK(clk), .Q(n90), .QN(n91) );
  DFFX4 E_reg_6_ ( .D(n4564), .CK(clk), .Q(SHA256_result[102]), .QN(n135) );
  DFFX4 F_reg_6_ ( .D(n4437), .CK(clk), .Q(n83), .QN(n82) );
  DFFX4 B_reg_2_ ( .D(n4696), .CK(clk), .Q(SHA256_result[194]), .QN(n1308) );
  DFFHQXL H5_reg_7_ ( .D(n4340), .CK(clk), .Q(H5[7]) );
  DFFHQXL H6_reg_1_ ( .D(n4378), .CK(clk), .Q(H6[1]) );
  DFFX4 E_reg_17_ ( .D(n4553), .CK(clk), .Q(SHA256_result[113]), .QN(n1367) );
  DFFHQX1 B_reg_25_ ( .D(n4673), .CK(clk), .Q(SHA256_result[217]) );
  DFFHQX2 B_reg_16_ ( .D(n4682), .CK(clk), .Q(SHA256_result[208]) );
  DFFHQX2 B_reg_20_ ( .D(n4678), .CK(clk), .Q(SHA256_result[212]) );
  DFFHQX2 B_reg_23_ ( .D(n4675), .CK(clk), .Q(SHA256_result[215]) );
  DFFHQX2 B_reg_19_ ( .D(n4679), .CK(clk), .Q(SHA256_result[211]) );
  DFFX2 A_reg_7_ ( .D(n4757), .CK(clk), .Q(n218), .QN(n217) );
  DFFX2 E_reg_11_ ( .D(n4559), .CK(clk), .Q(n138), .QN(n137) );
  DFFX1 mux_control_reg_1_ ( .D(n4701), .CK(clk), .QN(n439) );
  DFFX4 G_reg_4_ ( .D(n4407), .CK(clk), .Q(n73), .QN(n72) );
  DFFX4 E_reg_3_ ( .D(n4567), .CK(clk), .Q(n68), .QN(n67) );
  DFFTRX1 M_reg_19_ ( .D(M_w[19]), .RN(n404), .CK(clk), .Q(M[19]) );
  DFFTRX1 M_reg_18_ ( .D(M_w[18]), .RN(n256), .CK(clk), .Q(M[18]) );
  DFFTRX1 M_reg_15_ ( .D(M_w[15]), .RN(n256), .CK(clk), .Q(M[15]) );
  DFFTRX1 M_reg_14_ ( .D(M_w[14]), .RN(n256), .CK(clk), .Q(M[14]) );
  DFFTRX1 M_reg_13_ ( .D(M_w[13]), .RN(n256), .CK(clk), .Q(M[13]) );
  DFFTRX1 M_reg_12_ ( .D(M_w[12]), .RN(n403), .CK(clk), .Q(M[12]) );
  DFFTRX1 M_reg_11_ ( .D(M_w[11]), .RN(n256), .CK(clk), .Q(M[11]) );
  DFFTRX2 M_reg_9_ ( .D(M_w[9]), .RN(n401), .CK(clk), .Q(M[9]) );
  DFFTRX2 M_reg_6_ ( .D(M_w[6]), .RN(n402), .CK(clk), .Q(M[6]) );
  DFFTRX2 M_reg_5_ ( .D(M_w[5]), .RN(n402), .CK(clk), .Q(M[5]) );
  DFFTRX2 M_reg_4_ ( .D(M_w[4]), .RN(n402), .CK(clk), .Q(M[4]) );
  DFFTRX2 M_reg_2_ ( .D(M_w[2]), .RN(n402), .CK(clk), .Q(M[2]) );
  DFFTRX2 M_reg_1_ ( .D(M_w[1]), .RN(n402), .CK(clk), .Q(M[1]) );
  DFFTRX2 M_reg_0_ ( .D(M_w[0]), .RN(n402), .CK(clk), .Q(M[0]) );
  DFFHQX2 A_reg_10_ ( .D(n4754), .CK(clk), .Q(SHA256_result[234]) );
  DFFHQX2 A_reg_14_ ( .D(n4750), .CK(clk), .Q(SHA256_result[238]) );
  DFFHQX1 A_reg_17_ ( .D(n4747), .CK(clk), .Q(SHA256_result[241]) );
  DFFHQX2 B_reg_17_ ( .D(n4681), .CK(clk), .Q(SHA256_result[209]) );
  DFFHQX2 C_reg_17_ ( .D(n4649), .CK(clk), .Q(SHA256_result[177]) );
  DFFHQX2 E_reg_14_ ( .D(n4556), .CK(clk), .Q(SHA256_result[110]) );
  DFFHQX2 F_reg_16_ ( .D(n4427), .CK(clk), .Q(SHA256_result[80]) );
  DFFHQX2 F_reg_17_ ( .D(n4426), .CK(clk), .Q(SHA256_result[81]) );
  DFFHQX2 F_reg_21_ ( .D(n4422), .CK(clk), .Q(SHA256_result[85]) );
  DFFHQX2 F_reg_22_ ( .D(n4421), .CK(clk), .Q(SHA256_result[86]) );
  DFFHQX1 F_reg_23_ ( .D(n4420), .CK(clk), .Q(SHA256_result[87]) );
  DFFHQX2 G_reg_16_ ( .D(n4395), .CK(clk), .Q(SHA256_result[48]) );
  DFFHQX2 G_reg_17_ ( .D(n4394), .CK(clk), .Q(SHA256_result[49]) );
  DFFHQX2 G_reg_18_ ( .D(n4393), .CK(clk), .Q(SHA256_result[50]) );
  DFFHQX2 G_reg_20_ ( .D(n4391), .CK(clk), .Q(SHA256_result[52]) );
  DFFHQX2 G_reg_21_ ( .D(n4390), .CK(clk), .Q(SHA256_result[53]) );
  DFFHQX2 G_reg_22_ ( .D(n4389), .CK(clk), .Q(SHA256_result[54]) );
  DFFTRX2 L_reg_3_ ( .D(T1_32[3]), .RN(n401), .CK(clk), .Q(L[3]) );
  DFFTRX2 L_reg_4_ ( .D(T1_32[4]), .RN(n404), .CK(clk), .Q(L[4]) );
  DFFHQX2 C_reg_23_ ( .D(n4643), .CK(clk), .Q(SHA256_result[183]) );
  DFFHQX2 C_reg_22_ ( .D(n4644), .CK(clk), .Q(SHA256_result[182]) );
  DFFHQX2 C_reg_20_ ( .D(n4646), .CK(clk), .Q(SHA256_result[180]) );
  DFFHQX2 C_reg_21_ ( .D(n4645), .CK(clk), .Q(SHA256_result[181]) );
  DFFHQX2 C_reg_16_ ( .D(n4650), .CK(clk), .Q(SHA256_result[176]) );
  DFFTRX1 L_reg_0_ ( .D(T1_32[0]), .RN(n404), .CK(clk), .Q(L[0]) );
  DFFHQX2 B_reg_22_ ( .D(n4676), .CK(clk), .Q(SHA256_result[214]) );
  DFFHQX2 B_reg_21_ ( .D(n4677), .CK(clk), .Q(SHA256_result[213]) );
  DFFTRX2 M_reg_3_ ( .D(M_w[3]), .RN(n402), .CK(clk), .Q(M[3]) );
  DFFHQX1 H5_reg_1_ ( .D(n4346), .CK(clk), .Q(H5[1]) );
  DFFTRX1 L_reg_14_ ( .D(T1_32[14]), .RN(n404), .CK(clk), .Q(L[14]) );
  DFFTRX1 L_reg_13_ ( .D(n194), .RN(n404), .CK(clk), .Q(L[13]) );
  DFFTRX1 L_reg_11_ ( .D(T1_32[11]), .RN(n404), .CK(clk), .Q(L[11]) );
  DFFTRX1 L_reg_10_ ( .D(n175), .RN(n404), .CK(clk), .Q(L[10]) );
  DFFTRX1 L_reg_23_ ( .D(n12), .RN(n403), .CK(clk), .Q(L[23]) );
  DFFTRX1 L_reg_17_ ( .D(n71), .RN(n403), .CK(clk), .Q(L[17]) );
  DFFTRX1 L_reg_25_ ( .D(n155), .RN(n403), .CK(clk), .Q(L[25]) );
  DFFTRX1 L_reg_9_ ( .D(T1_32[9]), .RN(n404), .CK(clk), .Q(L[9]) );
  DFFHQX1 H1_reg_14_ ( .D(n4461), .CK(clk), .Q(H1[14]) );
  DFFTRX1 L_reg_8_ ( .D(n161), .RN(n404), .CK(clk), .Q(L[8]) );
  DFFTRX1 L_reg_19_ ( .D(T1_32[19]), .RN(n403), .CK(clk), .Q(L[19]) );
  DFFTRX1 L_reg_16_ ( .D(T1_32[16]), .RN(n403), .CK(clk), .Q(L[16]) );
  DFFTRX1 L_reg_12_ ( .D(T1_32[12]), .RN(n404), .CK(clk), .Q(L[12]) );
  DFFHQX1 C_reg_18_ ( .D(n4648), .CK(clk), .Q(SHA256_result[178]) );
  DFFTRX1 L_reg_2_ ( .D(T1_32[2]), .RN(n402), .CK(clk), .Q(L[2]) );
  DFFTRX1 L_reg_20_ ( .D(T1_32[20]), .RN(n403), .CK(clk), .Q(L[20]) );
  DFFTRX1 L_reg_22_ ( .D(T1_32[22]), .RN(n403), .CK(clk), .Q(L[22]) );
  DFFX1 C_reg_25_ ( .D(n4641), .CK(clk), .Q(n86), .QN(n87) );
  DFFTRX1 round_reg_5_ ( .D(N157), .RN(n4250), .CK(clk), .Q(round[5]), .QN(
        n2906) );
  DFFTRX1 L_reg_21_ ( .D(n17), .RN(n403), .CK(clk), .Q(L[21]) );
  DFFHQX4 F_reg_20_ ( .D(n4423), .CK(clk), .Q(SHA256_result[84]) );
  DFFHQX4 G_reg_19_ ( .D(n4392), .CK(clk), .Q(SHA256_result[51]) );
  DFFHQX4 B_reg_18_ ( .D(n4680), .CK(clk), .Q(SHA256_result[210]) );
  DFFHQX4 G_reg_25_ ( .D(n4386), .CK(clk), .Q(SHA256_result[57]) );
  DFFHQX4 G_reg_23_ ( .D(n4388), .CK(clk), .Q(SHA256_result[55]) );
  DFFHQX4 C_reg_11_ ( .D(n4655), .CK(clk), .Q(SHA256_result[171]) );
  DFFX4 E_reg_25_ ( .D(n4545), .CK(clk), .Q(n244), .QN(n243) );
  DFFHQX2 C_reg_19_ ( .D(n4647), .CK(clk), .Q(SHA256_result[179]) );
  DFFTRX2 M_reg_8_ ( .D(M_w[8]), .RN(n402), .CK(clk), .Q(M[8]) );
  DFFHQX4 C_reg_10_ ( .D(n4656), .CK(clk), .Q(SHA256_result[170]) );
  DFFHQX2 Kt_reg_1_ ( .D(N3134), .CK(clk), .Q(Kt[1]) );
  DFFHQX2 F_reg_19_ ( .D(n4424), .CK(clk), .Q(SHA256_result[83]) );
  DFFTRX2 M_reg_10_ ( .D(M_w[10]), .RN(n256), .CK(clk), .Q(M[10]) );
  DFFHQX2 F_reg_18_ ( .D(n4425), .CK(clk), .Q(SHA256_result[82]) );
  DFFTRX2 L_reg_27_ ( .D(T1_32[27]), .RN(n403), .CK(clk), .Q(L[27]) );
  OAI2BB1X4 U3 ( .A0N(n807), .A1N(N967), .B0(n701), .Y(n4540) );
  INVX1 U4 ( .A(n690), .Y(n11) );
  INVX4 U5 ( .A(SHA256_result[73]), .Y(n690) );
  NAND3BX1 U15 ( .AN(n447), .B(n1221), .C(n423), .Y(n798) );
  DLY1X1 U16 ( .A(next_E[22]), .Y(n198) );
  OAI211X1 U17 ( .A0(n334), .A1(n121), .B0(n615), .C0(n614), .Y(n4416) );
  AOI21XL U18 ( .A0(n343), .A1(SHA256_result[30]), .B0(n328), .Y(n451) );
  AOI21XL U19 ( .A0(n343), .A1(n111), .B0(n328), .Y(n730) );
  AOI21XL U20 ( .A0(SHA256_result[75]), .A1(n342), .B0(n328), .Y(n648) );
  AOI21XL U21 ( .A0(SHA256_result[77]), .A1(n342), .B0(n328), .Y(n643) );
  AOI21XL U22 ( .A0(SHA256_result[78]), .A1(n342), .B0(n328), .Y(n641) );
  NOR3X1 U23 ( .A(n444), .B(n1246), .C(n811), .Y(n445) );
  NAND4X4 U24 ( .A(n717), .B(n718), .C(n802), .D(n716), .Y(n4546) );
  NAND4X2 U25 ( .A(n1128), .B(n1127), .C(n384), .D(n1126), .Y(n4745) );
  DLY1X1 U26 ( .A(T1_32[23]), .Y(n12) );
  NAND2X2 U27 ( .A(n229), .B(n177), .Y(n4545) );
  AOI2BB1X2 U28 ( .A0N(n2878), .A1N(n3580), .B0(n3577), .Y(n3579) );
  INVX16 U29 ( .A(n3517), .Y(n1244) );
  INVX20 U30 ( .A(n75), .Y(n419) );
  NAND2X4 U31 ( .A(N961), .B(n807), .Y(n717) );
  OAI2BB1X4 U32 ( .A0N(SHA256_result[199]), .A1N(n218), .B0(n1076), .Y(
        f2_ABC_32[7]) );
  OAI21X4 U33 ( .A0(n317), .A1(n96), .B0(SHA256_result[160]), .Y(n1083) );
  BUFX16 U34 ( .A(SHA256_result[224]), .Y(n317) );
  NAND2X4 U35 ( .A(n1085), .B(n1084), .Y(n4733) );
  CLKBUFX3 U36 ( .A(next_E[25]), .Y(n188) );
  INVX8 U37 ( .A(SHA256_result[45]), .Y(n684) );
  INVX8 U38 ( .A(n145), .Y(n146) );
  OAI21X1 U39 ( .A0(n300), .A1(SHA256_result[216]), .B0(SHA256_result[184]), 
        .Y(n1059) );
  BUFX4 U40 ( .A(SHA256_result[235]), .Y(n14) );
  BUFX1 U41 ( .A(SHA256_result[235]), .Y(n15) );
  BUFX4 U42 ( .A(SHA256_result[235]), .Y(n16) );
  MX2X1 U43 ( .A(SHA256_result[51]), .B(SHA256_result[83]), .S0(n111), .Y(
        f1_EFG_32[19]) );
  DLY1X1 U44 ( .A(T1_32[13]), .Y(n194) );
  INVX8 U45 ( .A(n1243), .Y(n1221) );
  CLKINVX3 U46 ( .A(n3115), .Y(n421) );
  DLY1X1 U47 ( .A(T1_32[17]), .Y(n71) );
  BUFX16 U48 ( .A(T1_32[21]), .Y(n17) );
  AOI22X2 U49 ( .A0(N1087), .A1(n353), .B0(n302), .B1(n247), .Y(n1121) );
  CLKINVX8 U50 ( .A(SHA256_result[43]), .Y(n688) );
  XOR3X2 U51 ( .A(SHA256_result[102]), .B(n139), .C(n244), .Y(f4_E_32[0]) );
  INVX1 U52 ( .A(round[0]), .Y(n430) );
  INVX8 U53 ( .A(SHA256_result[65]), .Y(n698) );
  NAND2X4 U54 ( .A(n1117), .B(n1116), .Y(n4741) );
  AOI22X4 U55 ( .A0(N1088), .A1(n353), .B0(n301), .B1(n247), .Y(n1117) );
  INVX4 U56 ( .A(SHA256_result[75]), .Y(n687) );
  DLY1X1 U57 ( .A(T1_32[10]), .Y(n175) );
  INVX8 U58 ( .A(SHA256_result[74]), .Y(n689) );
  INVX2 U59 ( .A(n802), .Y(n328) );
  INVX1 U60 ( .A(n802), .Y(n329) );
  INVX8 U61 ( .A(n73), .Y(n1210) );
  OAI21X2 U62 ( .A0(n299), .A1(SHA256_result[217]), .B0(n86), .Y(n1058) );
  BUFX16 U63 ( .A(SHA256_result[232]), .Y(n18) );
  MX2X2 U64 ( .A(SHA256_result[57]), .B(SHA256_result[89]), .S0(n244), .Y(
        f1_EFG_32[25]) );
  NAND2X2 U65 ( .A(n3377), .B(n811), .Y(n816) );
  NAND2X2 U66 ( .A(n1221), .B(round[6]), .Y(n811) );
  NOR2X2 U67 ( .A(n3503), .B(n3574), .Y(n3377) );
  OAI21X2 U68 ( .A0(n14), .A1(SHA256_result[203]), .B0(SHA256_result[171]), 
        .Y(n1072) );
  BUFX12 U69 ( .A(SHA256_result[242]), .Y(n306) );
  AOI221XL U70 ( .A0(n318), .A1(n1224), .B0(n258), .B1(n320), .C0(n4096), .Y(
        n4156) );
  CLKBUFX8 U71 ( .A(round[4]), .Y(n318) );
  INVX12 U72 ( .A(n359), .Y(n354) );
  INVX3 U73 ( .A(n373), .Y(n359) );
  INVX1 U74 ( .A(n396), .Y(n20) );
  INVX8 U75 ( .A(n398), .Y(n21) );
  INVX12 U76 ( .A(n394), .Y(n22) );
  INVX12 U77 ( .A(n392), .Y(n23) );
  INVX4 U78 ( .A(n393), .Y(n24) );
  INVX4 U79 ( .A(n391), .Y(n25) );
  INVX4 U80 ( .A(n397), .Y(n26) );
  INVX20 U81 ( .A(n396), .Y(n27) );
  INVX8 U82 ( .A(n395), .Y(n28) );
  INVXL U83 ( .A(n1200), .Y(n29) );
  INVX1 U84 ( .A(n20), .Y(n30) );
  INVX1 U85 ( .A(n288), .Y(n396) );
  INVX16 U86 ( .A(n380), .Y(n390) );
  INVXL U87 ( .A(n386), .Y(n380) );
  NAND2X2 U88 ( .A(N962), .B(n807), .Y(n229) );
  OAI21X4 U89 ( .A0(SHA256_result[200]), .A1(n18), .B0(SHA256_result[168]), 
        .Y(n1075) );
  OAI2BB1X4 U90 ( .A0N(SHA256_result[200]), .A1N(n18), .B0(n1075), .Y(
        f2_ABC_32[8]) );
  MX2X4 U91 ( .A(SHA256_result[55]), .B(SHA256_result[87]), .S0(n90), .Y(
        f1_EFG_32[23]) );
  AOI21X1 U92 ( .A0(n344), .A1(SHA256_result[55]), .B0(n326), .Y(n547) );
  BUFX3 U93 ( .A(SHA256_result[88]), .Y(n31) );
  AOI21X1 U94 ( .A0(n344), .A1(SHA256_result[57]), .B0(n326), .Y(n541) );
  XOR3X4 U95 ( .A(n154), .B(n147), .C(n117), .Y(f4_E_32[1]) );
  INVX4 U96 ( .A(n145), .Y(n147) );
  OAI21X4 U97 ( .A0(SHA256_result[210]), .A1(n306), .B0(n32), .Y(n1065) );
  BUFX8 U98 ( .A(SHA256_result[178]), .Y(n32) );
  MX2X4 U99 ( .A(SHA256_result[52]), .B(SHA256_result[84]), .S0(
        SHA256_result[116]), .Y(f1_EFG_32[20]) );
  OAI21X4 U100 ( .A0(SHA256_result[209]), .A1(n307), .B0(SHA256_result[177]), 
        .Y(n1066) );
  OAI2BB1X4 U101 ( .A0N(SHA256_result[209]), .A1N(n307), .B0(n1066), .Y(
        f2_ABC_32[17]) );
  BUFX12 U102 ( .A(SHA256_result[241]), .Y(n307) );
  MX2X2 U103 ( .A(SHA256_result[54]), .B(SHA256_result[86]), .S0(
        SHA256_result[118]), .Y(f1_EFG_32[22]) );
  BUFX3 U104 ( .A(SHA256_result[252]), .Y(n296) );
  AND2X2 U105 ( .A(first_block_core), .B(n815), .Y(n261) );
  INVX1 U106 ( .A(n230), .Y(n232) );
  CLKINVX3 U107 ( .A(n795), .Y(n336) );
  BUFX3 U108 ( .A(SHA256_result[251]), .Y(n297) );
  CLKBUFX8 U109 ( .A(SHA256_result[249]), .Y(n299) );
  BUFX3 U110 ( .A(SHA256_result[248]), .Y(n300) );
  CLKINVX3 U111 ( .A(n423), .Y(n422) );
  NOR2BX1 U112 ( .AN(n4070), .B(n434), .Y(n3955) );
  CLKINVX3 U113 ( .A(n802), .Y(n326) );
  CLKINVX3 U114 ( .A(n346), .Y(n344) );
  CLKINVX3 U115 ( .A(n802), .Y(n327) );
  CLKINVX3 U116 ( .A(n346), .Y(n343) );
  INVX4 U117 ( .A(SHA256_result[110]), .Y(n746) );
  CLKINVX3 U118 ( .A(n346), .Y(n342) );
  INVX4 U119 ( .A(n338), .Y(n332) );
  INVX1 U120 ( .A(n322), .Y(n176) );
  CLKINVX3 U121 ( .A(n346), .Y(n345) );
  INVX2 U122 ( .A(n360), .Y(n353) );
  OAI21X2 U123 ( .A0(SHA256_result[212]), .A1(n304), .B0(SHA256_result[180]), 
        .Y(n1063) );
  OAI2BB1X2 U124 ( .A0N(SHA256_result[206]), .A1N(n310), .B0(n1069), .Y(
        f2_ABC_32[14]) );
  OAI21X2 U125 ( .A0(SHA256_result[206]), .A1(n310), .B0(SHA256_result[174]), 
        .Y(n1069) );
  OAI21X2 U126 ( .A0(SHA256_result[204]), .A1(SHA256_result[236]), .B0(
        SHA256_result[172]), .Y(n1071) );
  OAI2BB1X2 U127 ( .A0N(SHA256_result[201]), .A1N(n312), .B0(n1074), .Y(
        f2_ABC_32[9]) );
  MX2X2 U128 ( .A(SHA256_result[53]), .B(SHA256_result[85]), .S0(
        SHA256_result[117]), .Y(f1_EFG_32[21]) );
  CLKBUFX8 U129 ( .A(f1_EFG_32[0]), .Y(n284) );
  NAND3X2 U130 ( .A(n3578), .B(n3564), .C(n3579), .Y(n3503) );
  CLKINVX3 U131 ( .A(n152), .Y(n154) );
  CLKINVX3 U132 ( .A(n2943), .Y(n428) );
  INVX4 U133 ( .A(SHA256_result[35]), .Y(n1212) );
  BUFX1 U134 ( .A(SHA256_result[98]), .Y(n282) );
  NAND2X1 U135 ( .A(round[6]), .B(n1219), .Y(n447) );
  NAND2X1 U136 ( .A(n261), .B(n816), .Y(n1198) );
  INVX1 U137 ( .A(n1186), .Y(n373) );
  INVX1 U138 ( .A(n443), .Y(n812) );
  NAND2X1 U139 ( .A(n4057), .B(n4249), .Y(n3378) );
  INVX4 U140 ( .A(n173), .Y(n1208) );
  INVX4 U141 ( .A(n133), .Y(n692) );
  INVX4 U142 ( .A(SHA256_result[44]), .Y(n686) );
  INVX4 U143 ( .A(SHA256_result[46]), .Y(n682) );
  CLKINVX3 U144 ( .A(n95), .Y(n1246) );
  CLKBUFX8 U145 ( .A(SHA256_result[244]), .Y(n304) );
  BUFX4 U146 ( .A(SHA256_result[245]), .Y(n303) );
  NAND2X2 U147 ( .A(n249), .B(n2938), .Y(n1300) );
  BUFX3 U148 ( .A(SHA256_result[254]), .Y(n294) );
  BUFX3 U149 ( .A(SHA256_result[253]), .Y(n295) );
  BUFX3 U150 ( .A(SHA256_result[250]), .Y(n298) );
  AOI222XL U151 ( .A0(n258), .A1(n4000), .B0(n4055), .B1(n4056), .C0(n319), 
        .C1(n4015), .Y(n4048) );
  INVX16 U152 ( .A(n421), .Y(n420) );
  NOR2X2 U153 ( .A(round[0]), .B(n319), .Y(n4042) );
  INVX2 U154 ( .A(SHA256_result[78]), .Y(n681) );
  INVX1 U155 ( .A(n183), .Y(n184) );
  BUFX3 U156 ( .A(SHA256_result[38]), .Y(n143) );
  CLKBUFX8 U157 ( .A(SHA256_result[114]), .Y(n291) );
  INVX4 U158 ( .A(SHA256_result[108]), .Y(n145) );
  BUFX3 U159 ( .A(n282), .Y(n185) );
  INVX12 U160 ( .A(n798), .Y(n807) );
  INVX1 U161 ( .A(N937), .Y(n797) );
  CLKINVX3 U162 ( .A(n381), .Y(n389) );
  BUFX8 U163 ( .A(SHA256_result[238]), .Y(n310) );
  INVX8 U164 ( .A(n400), .Y(n399) );
  INVX1 U165 ( .A(n1201), .Y(n400) );
  NAND2X1 U166 ( .A(n1223), .B(n433), .Y(n809) );
  INVX1 U167 ( .A(n178), .Y(n177) );
  NAND2BX1 U168 ( .AN(n179), .B(n714), .Y(n178) );
  OAI21XL U169 ( .A0(n28), .A1(n1106), .B0(n990), .Y(n992) );
  NAND2X2 U170 ( .A(N954), .B(n807), .Y(n735) );
  OAI211X1 U171 ( .A0(n411), .A1(n162), .B0(n3203), .C0(n419), .Y(n4378) );
  OAI211X1 U172 ( .A0(n412), .A1(n131), .B0(n3184), .C0(n419), .Y(n4340) );
  NAND2X2 U173 ( .A(n190), .B(n76), .Y(n4547) );
  NAND2X2 U174 ( .A(N960), .B(n807), .Y(n190) );
  INVX1 U175 ( .A(n196), .Y(n195) );
  INVX1 U176 ( .A(n192), .Y(n191) );
  INVX1 U177 ( .A(n200), .Y(n199) );
  OAI211X1 U178 ( .A0(n335), .A1(n131), .B0(n587), .C0(n586), .Y(n4404) );
  OAI211X1 U179 ( .A0(n335), .A1(n211), .B0(n600), .C0(n599), .Y(n4409) );
  NAND3X1 U180 ( .A(n248), .B(n773), .C(n772), .Y(n4563) );
  BUFX3 U181 ( .A(T1_32[8]), .Y(n161) );
  BUFX3 U182 ( .A(T1_32[25]), .Y(n155) );
  OAI21XL U183 ( .A0(n23), .A1(n1119), .B0(n998), .Y(n1000) );
  OAI21XL U184 ( .A0(n420), .A1(n860), .B0(n859), .Y(n4593) );
  OAI21XL U185 ( .A0(n420), .A1(n867), .B0(n866), .Y(n4595) );
  OAI21XL U186 ( .A0(n420), .A1(n937), .B0(n936), .Y(n4495) );
  OAI21XL U187 ( .A0(n420), .A1(n941), .B0(n940), .Y(n4496) );
  OAI21XL U188 ( .A0(n420), .A1(n951), .B0(n950), .Y(n4499) );
  OAI21XL U189 ( .A0(n420), .A1(n82), .B0(n661), .Y(n4341) );
  OAI21XL U190 ( .A0(n420), .A1(n668), .B0(n667), .Y(n4343) );
  OAI21XL U191 ( .A0(n420), .A1(n870), .B0(n869), .Y(n4596) );
  AOI21X1 U192 ( .A0(SHA256_result[0]), .A1(n342), .B0(n326), .Y(n524) );
  OAI21XL U193 ( .A0(n27), .A1(n964), .B0(n881), .Y(n883) );
  OAI21XL U194 ( .A0(n21), .A1(n957), .B0(n873), .Y(n875) );
  OAI21XL U195 ( .A0(n27), .A1(n960), .B0(n877), .Y(n879) );
  OAI21XL U196 ( .A0(n25), .A1(n947), .B0(n863), .Y(n865) );
  OAI21XL U197 ( .A0(n22), .A1(n969), .B0(n888), .Y(n890) );
  OAI21XL U198 ( .A0(n420), .A1(n885), .B0(n884), .Y(n4600) );
  OAI21XL U199 ( .A0(n420), .A1(n964), .B0(n963), .Y(n4503) );
  OAI211X1 U200 ( .A0(n407), .A1(n211), .B0(n3186), .C0(n419), .Y(n4345) );
  OAI21XL U201 ( .A0(n420), .A1(n892), .B0(n891), .Y(n4602) );
  AOI21X1 U202 ( .A0(n344), .A1(SHA256_result[59]), .B0(n326), .Y(n535) );
  OAI21XL U203 ( .A0(n23), .A1(n1111), .B0(n993), .Y(n995) );
  OAI211X1 U204 ( .A0(n333), .A1(n141), .B0(n520), .C0(n519), .Y(n4312) );
  OAI21XL U205 ( .A0(n24), .A1(n1051), .B0(n977), .Y(n979) );
  OAI21XL U206 ( .A0(n420), .A1(n125), .B0(n760), .Y(n4528) );
  OAI211X1 U207 ( .A0(n406), .A1(n763), .B0(n3314), .C0(n419), .Y(n4529) );
  OAI221XL U208 ( .A0(n287), .A1(n480), .B0(n1393), .B1(n795), .C0(n479), .Y(
        n4294) );
  OAI21XL U209 ( .A0(n420), .A1(n768), .B0(n767), .Y(n4530) );
  AOI21X1 U210 ( .A0(n343), .A1(SHA256_result[28]), .B0(n329), .Y(n456) );
  OAI21XL U211 ( .A0(n420), .A1(n104), .B0(n804), .Y(n4507) );
  AOI222XL U212 ( .A0(n3954), .A1(n253), .B0(n4225), .B1(n432), .C0(n4239), 
        .C1(n425), .Y(n4235) );
  AOI222XL U213 ( .A0(n4149), .A1(n425), .B0(n253), .B1(n257), .C0(n1289), 
        .C1(n422), .Y(n4195) );
  BUFX3 U214 ( .A(T1_32[18]), .Y(n169) );
  NAND2X1 U215 ( .A(n1097), .B(n1096), .Y(n4736) );
  AOI2BB2X1 U216 ( .B0(N1093), .B1(n353), .A0N(n1095), .A1N(n204), .Y(n1097)
         );
  NAND4X2 U217 ( .A(n1100), .B(n1101), .C(n381), .D(n1099), .Y(n4737) );
  AOI221X1 U218 ( .A0(n3954), .A1(n422), .B0(n3960), .B1(n258), .C0(n4170), 
        .Y(n4169) );
  OAI21XL U219 ( .A0(n420), .A1(n220), .B0(n1184), .Y(n4730) );
  OAI221XL U220 ( .A0(n287), .A1(n551), .B0(n1378), .B1(n330), .C0(n550), .Y(
        n4389) );
  OAI211X1 U221 ( .A0(n330), .A1(n683), .B0(n573), .C0(n572), .Y(n4398) );
  AOI21X1 U222 ( .A0(SHA256_result[44]), .A1(n342), .B0(n327), .Y(n574) );
  AOI21X1 U223 ( .A0(n208), .A1(n342), .B0(n327), .Y(n596) );
  OAI221XL U224 ( .A0(n287), .A1(n627), .B0(n1370), .B1(n795), .C0(n626), .Y(
        n4422) );
  NAND2X1 U225 ( .A(n728), .B(n727), .Y(n4550) );
  AOI2BB2X2 U226 ( .B0(N957), .B1(n807), .A0N(n180), .A1N(n1369), .Y(n728) );
  NAND2X1 U227 ( .A(n741), .B(n740), .Y(n4554) );
  AOI22X2 U228 ( .A0(N953), .A1(n807), .B0(SHA256_result[112]), .B1(n323), .Y(
        n741) );
  INVX1 U229 ( .A(n322), .Y(n187) );
  NAND4X1 U230 ( .A(n749), .B(n748), .C(n802), .D(n747), .Y(n4556) );
  NAND2X1 U231 ( .A(N951), .B(n807), .Y(n748) );
  NAND3X1 U232 ( .A(n252), .B(n753), .C(n752), .Y(n4557) );
  OAI222XL U233 ( .A0(n28), .A1(n939), .B0(n367), .B1(n938), .C0(n351), .C1(
        n937), .Y(n4655) );
  OAI21XL U234 ( .A0(n21), .A1(n1151), .B0(n1021), .Y(n1023) );
  OAI21XL U235 ( .A0(n22), .A1(n1154), .B0(n1024), .Y(n1026) );
  OAI21XL U236 ( .A0(n22), .A1(n1158), .B0(n1027), .Y(n1029) );
  OAI21XL U237 ( .A0(n23), .A1(n217), .B0(n1032), .Y(n1034) );
  NAND4X1 U238 ( .A(n1138), .B(n1137), .C(n383), .D(n1136), .Y(n4749) );
  NAND2X1 U239 ( .A(N1080), .B(n357), .Y(n1137) );
  OAI21XL U240 ( .A0(n24), .A1(n1160), .B0(n1159), .Y(n1162) );
  OAI21XL U241 ( .A0(n24), .A1(n1172), .B0(n1171), .Y(n1174) );
  OAI21XL U242 ( .A0(n26), .A1(n1177), .B0(n1176), .Y(n1179) );
  OAI21XL U243 ( .A0(n21), .A1(n1190), .B0(n1189), .Y(n1192) );
  OAI21XL U244 ( .A0(n23), .A1(n1195), .B0(n1194), .Y(n1197) );
  OAI21XL U245 ( .A0(n24), .A1(n1199), .B0(n380), .Y(n1204) );
  AOI21X1 U246 ( .A0(n323), .A1(SHA256_result[31]), .B0(n445), .Y(n446) );
  INVX1 U247 ( .A(n67), .Y(n69) );
  CLKBUFX2 U248 ( .A(n69), .Y(n283) );
  DLY1X1 U249 ( .A(next_E[27]), .Y(n70) );
  INVX1 U250 ( .A(n72), .Y(n74) );
  NOR2X1 U251 ( .A(n809), .B(n253), .Y(n3580) );
  NOR2X2 U252 ( .A(n2946), .B(n430), .Y(n253) );
  CLKINVX3 U253 ( .A(n435), .Y(n434) );
  INVX2 U254 ( .A(n413), .Y(n412) );
  CLKINVX3 U255 ( .A(n416), .Y(n407) );
  INVX2 U256 ( .A(n415), .Y(n408) );
  INVX1 U257 ( .A(n323), .Y(n180) );
  CLKINVX3 U258 ( .A(n107), .Y(n406) );
  CLKINVX3 U259 ( .A(n338), .Y(n331) );
  CLKINVX3 U260 ( .A(n339), .Y(n330) );
  NAND2X2 U261 ( .A(n261), .B(n450), .Y(n802) );
  INVX1 U262 ( .A(n415), .Y(n409) );
  CLKINVX3 U263 ( .A(n336), .Y(n335) );
  CLKINVX3 U264 ( .A(n135), .Y(n136) );
  INVX1 U265 ( .A(mux_control_0_), .Y(n436) );
  CLKINVX3 U266 ( .A(n247), .Y(n204) );
  INVX1 U267 ( .A(n125), .Y(n127) );
  INVX4 U268 ( .A(n325), .Y(n323) );
  CLKINVX3 U269 ( .A(n325), .Y(n322) );
  INVX1 U270 ( .A(n414), .Y(n410) );
  INVX1 U271 ( .A(n1244), .Y(n414) );
  CLKINVX3 U272 ( .A(n337), .Y(n333) );
  AND2X2 U273 ( .A(first_block_core), .B(n414), .Y(n75) );
  BUFX3 U274 ( .A(round[3]), .Y(n319) );
  CLKINVX3 U275 ( .A(n336), .Y(n334) );
  INVX1 U276 ( .A(n334), .Y(n340) );
  INVX1 U277 ( .A(n262), .Y(n3116) );
  NOR2X1 U278 ( .A(n226), .B(n189), .Y(n76) );
  INVX1 U279 ( .A(n374), .Y(n358) );
  NOR2X2 U280 ( .A(n1430), .B(read_counter[3]), .Y(n77) );
  AND2X2 U281 ( .A(read_counter[3]), .B(n1430), .Y(n78) );
  NOR2X2 U282 ( .A(read_counter[3]), .B(read_counter[2]), .Y(n79) );
  AND2X2 U283 ( .A(read_counter[3]), .B(read_counter[2]), .Y(n80) );
  INVX1 U284 ( .A(round[5]), .Y(n435) );
  INVX1 U285 ( .A(n125), .Y(n202) );
  CLKINVX3 U286 ( .A(n220), .Y(n222) );
  CLKINVX3 U287 ( .A(n170), .Y(n171) );
  CLKINVX3 U288 ( .A(n217), .Y(n219) );
  INVX1 U289 ( .A(n128), .Y(n130) );
  BUFX3 U290 ( .A(SHA256_result[255]), .Y(n293) );
  BUFX16 U291 ( .A(SHA256_result[111]), .Y(n280) );
  BUFX16 U292 ( .A(n3116), .Y(n205) );
  INVXL U293 ( .A(n689), .Y(n81) );
  BUFX3 U294 ( .A(SHA256_result[104]), .Y(n210) );
  INVX1 U295 ( .A(n82), .Y(n84) );
  BUFX3 U296 ( .A(SHA256_result[105]), .Y(n281) );
  BUFX3 U297 ( .A(SHA256_result[72]), .Y(n85) );
  INVX4 U298 ( .A(SHA256_result[72]), .Y(n691) );
  INVX1 U299 ( .A(n1181), .Y(n88) );
  INVX4 U300 ( .A(SHA256_result[67]), .Y(n696) );
  INVX1 U301 ( .A(n208), .Y(n89) );
  BUFX3 U302 ( .A(n144), .Y(n208) );
  NAND2X2 U303 ( .A(n724), .B(n723), .Y(n4548) );
  INVX1 U304 ( .A(n92), .Y(n94) );
  BUFX8 U305 ( .A(n1200), .Y(n288) );
  AOI22X4 U306 ( .A0(N1091), .A1(n353), .B0(n298), .B1(n247), .Y(n1105) );
  NAND2X4 U307 ( .A(N1092), .B(n357), .Y(n1100) );
  NOR2BX2 U308 ( .AN(n1223), .B(n2947), .Y(n95) );
  CLKINVX2 U309 ( .A(n1300), .Y(n1223) );
  AOI2BB2X4 U310 ( .B0(N958), .B1(n807), .A0N(n324), .A1N(n1370), .Y(n726) );
  INVX1 U311 ( .A(n98), .Y(n100) );
  INVX1 U312 ( .A(n101), .Y(n103) );
  INVX1 U313 ( .A(n104), .Y(n106) );
  INVXL U314 ( .A(n1244), .Y(n107) );
  INVXL U315 ( .A(n414), .Y(n411) );
  NOR3XL U316 ( .A(n3116), .B(n3577), .C(n3578), .Y(n3517) );
  INVXL U317 ( .A(n1244), .Y(n415) );
  INVXL U318 ( .A(n1244), .Y(n413) );
  INVXL U319 ( .A(n1244), .Y(n416) );
  INVX1 U320 ( .A(n108), .Y(n110) );
  NAND2X2 U321 ( .A(n3378), .B(n3377), .Y(n450) );
  INVX1 U322 ( .A(n113), .Y(n115) );
  INVX1 U323 ( .A(SHA256_result[112]), .Y(n739) );
  INVX1 U324 ( .A(n116), .Y(n118) );
  CLKINVX3 U325 ( .A(n121), .Y(n123) );
  INVXL U326 ( .A(n1186), .Y(n124) );
  OR3X2 U327 ( .A(n809), .B(n808), .C(n811), .Y(n1186) );
  MXI2X4 U328 ( .A(n683), .B(n684), .S0(n170), .Y(f1_EFG_32[13]) );
  INVX4 U329 ( .A(SHA256_result[76]), .Y(n685) );
  INVX1 U330 ( .A(n167), .Y(n131) );
  DLY1X1 U331 ( .A(SHA256_result[100]), .Y(n292) );
  INVX1 U332 ( .A(n132), .Y(n134) );
  CLKINVX8 U333 ( .A(n137), .Y(n139) );
  INVXL U334 ( .A(n1210), .Y(n140) );
  INVX1 U335 ( .A(n234), .Y(n141) );
  INVXL U336 ( .A(n1214), .Y(n234) );
  INVX4 U337 ( .A(n151), .Y(n1214) );
  INVX4 U338 ( .A(SHA256_result[77]), .Y(n683) );
  NAND2BX4 U339 ( .AN(n3577), .B(output_enable), .Y(n3564) );
  INVXL U340 ( .A(n696), .Y(n142) );
  INVXL U341 ( .A(n1212), .Y(n144) );
  CLKINVX2 U342 ( .A(n358), .Y(n357) );
  NAND2XL U343 ( .A(N985), .B(n354), .Y(n844) );
  NAND2XL U344 ( .A(N981), .B(n354), .Y(n852) );
  NAND2XL U345 ( .A(N983), .B(n354), .Y(n848) );
  NAND2XL U346 ( .A(N984), .B(n354), .Y(n846) );
  NAND2XL U347 ( .A(N991), .B(n354), .Y(n832) );
  NAND2XL U348 ( .A(N986), .B(n354), .Y(n842) );
  NAND2XL U349 ( .A(N987), .B(n354), .Y(n840) );
  NAND2XL U350 ( .A(N988), .B(n354), .Y(n838) );
  NAND2XL U351 ( .A(N993), .B(n354), .Y(n828) );
  NAND2XL U352 ( .A(N1015), .B(n354), .Y(n930) );
  INVX1 U353 ( .A(n211), .Y(n213) );
  INVX4 U354 ( .A(n212), .Y(n697) );
  AOI21X1 U355 ( .A0(SHA256_result[46]), .A1(n342), .B0(n327), .Y(n569) );
  CLKBUFX2 U356 ( .A(SHA256_result[96]), .Y(n285) );
  CLKINVX3 U357 ( .A(n148), .Y(n150) );
  AOI21XL U358 ( .A0(n343), .A1(SHA256_result[113]), .B0(n329), .Y(n736) );
  CLKINVX3 U359 ( .A(n156), .Y(n158) );
  NAND2X2 U360 ( .A(n745), .B(n744), .Y(n4555) );
  INVX1 U361 ( .A(n162), .Y(n164) );
  OAI21XL U362 ( .A0(n420), .A1(n152), .B0(n771), .Y(n4531) );
  INVX4 U363 ( .A(SHA256_result[109]), .Y(n170) );
  INVX1 U364 ( .A(n172), .Y(n174) );
  OAI211X1 U365 ( .A0(n333), .A1(n698), .B0(n602), .C0(n601), .Y(n4410) );
  OR2X4 U366 ( .A(n3577), .B(output_enable), .Y(n1243) );
  AND2X2 U367 ( .A(n3503), .B(n3564), .Y(n262) );
  AOI2BB2X4 U368 ( .B0(N959), .B1(n807), .A0N(n722), .A1N(n176), .Y(n724) );
  AND2X1 U369 ( .A(n244), .B(n323), .Y(n179) );
  AOI22X2 U370 ( .A0(N1076), .A1(n353), .B0(n16), .B1(n247), .Y(n1153) );
  NAND4X4 U371 ( .A(n1088), .B(n1089), .C(n384), .D(n1087), .Y(n4734) );
  INVXL U372 ( .A(n698), .Y(n181) );
  OAI21XL U373 ( .A0(n420), .A1(n698), .B0(n675), .Y(n4346) );
  INVX4 U374 ( .A(n163), .Y(n182) );
  INVX4 U375 ( .A(SHA256_result[40]), .Y(n183) );
  AOI21XL U376 ( .A0(next_E[30]), .A1(n336), .B0(n700), .Y(n701) );
  OAI211X1 U377 ( .A0(n333), .A1(n128), .B0(n592), .C0(n591), .Y(n4406) );
  NAND2X2 U378 ( .A(n1153), .B(n1152), .Y(n4753) );
  NAND2X1 U379 ( .A(N972), .B(n371), .Y(n881) );
  NAND2X2 U380 ( .A(N1094), .B(n357), .Y(n1092) );
  NAND2X4 U381 ( .A(N1095), .B(n357), .Y(n1088) );
  NAND2X1 U382 ( .A(n94), .B(n345), .Y(n706) );
  BUFX8 U383 ( .A(next_E[10]), .Y(n186) );
  AOI2BB2X4 U384 ( .B0(N952), .B1(n807), .A0N(n743), .A1N(n187), .Y(n745) );
  INVX8 U385 ( .A(n324), .Y(n321) );
  NAND2X2 U386 ( .A(n1105), .B(n1104), .Y(n4738) );
  INVX1 U387 ( .A(n720), .Y(n189) );
  BUFX16 U388 ( .A(next_E[26]), .Y(n209) );
  NAND2X4 U389 ( .A(N955), .B(n807), .Y(n732) );
  OAI2BB1X4 U390 ( .A0N(n807), .A1N(N968), .B0(n806), .Y(n4539) );
  NAND2X4 U391 ( .A(n233), .B(n191), .Y(n4544) );
  NAND2BX1 U392 ( .AN(n193), .B(n712), .Y(n192) );
  AND2X1 U393 ( .A(n118), .B(n323), .Y(n193) );
  NAND2X4 U394 ( .A(n214), .B(n195), .Y(n4541) );
  NAND2BX1 U395 ( .AN(n197), .B(n704), .Y(n196) );
  AND2X1 U396 ( .A(n110), .B(n323), .Y(n197) );
  OAI211X2 U397 ( .A0(n332), .A1(n734), .B0(n733), .C0(n732), .Y(n4552) );
  NAND4X2 U398 ( .A(n1093), .B(n1092), .C(n383), .D(n1091), .Y(n4735) );
  INVX3 U399 ( .A(n1198), .Y(n386) );
  NAND2X4 U400 ( .A(n235), .B(n199), .Y(n4543) );
  NAND2BX1 U401 ( .AN(n201), .B(n710), .Y(n200) );
  AND2X1 U402 ( .A(n123), .B(n323), .Y(n201) );
  NAND2X4 U403 ( .A(N963), .B(n807), .Y(n233) );
  NAND3X2 U404 ( .A(n251), .B(n762), .C(n761), .Y(n4560) );
  CLKINVX8 U405 ( .A(n746), .Y(n203) );
  AOI2BB2X4 U406 ( .B0(N1096), .B1(n353), .A0N(n1051), .A1N(n204), .Y(n1085)
         );
  CLKINVX3 U407 ( .A(n439), .Y(n437) );
  OAI211X2 U408 ( .A0(n331), .A1(n737), .B0(n735), .C0(n736), .Y(n4553) );
  OAI211X1 U409 ( .A0(n1311), .A1(n24), .B0(n956), .C0(n955), .Y(n4660) );
  OAI211X1 U410 ( .A0(n1310), .A1(n27), .B0(n959), .C0(n958), .Y(n4661) );
  OAI211X1 U411 ( .A0(n1317), .A1(n28), .B0(n928), .C0(n927), .Y(n4651) );
  OAI211X1 U412 ( .A0(n1315), .A1(n24), .B0(n932), .C0(n931), .Y(n4653) );
  OAI211X1 U413 ( .A0(n1307), .A1(n23), .B0(n971), .C0(n970), .Y(n4665) );
  OAI211X1 U414 ( .A0(n1322), .A1(n28), .B0(n915), .C0(n914), .Y(n4645) );
  OAI211X1 U415 ( .A0(n1320), .A1(n23), .B0(n919), .C0(n918), .Y(n4647) );
  OAI211X1 U416 ( .A0(n411), .A1(n1205), .B0(n3576), .C0(n419), .Y(n4765) );
  OAI211X1 U417 ( .A0(n407), .A1(n969), .B0(n3305), .C0(n419), .Y(n4505) );
  OAI211X1 U418 ( .A0(n406), .A1(n1317), .B0(n419), .C0(n3280), .Y(n4460) );
  OAI211X1 U419 ( .A0(n412), .A1(n1315), .B0(n419), .C0(n3281), .Y(n4462) );
  OAI211X1 U420 ( .A0(n406), .A1(n939), .B0(n419), .C0(n3282), .Y(n4464) );
  OAI211X1 U421 ( .A0(n406), .A1(n943), .B0(n419), .C0(n3283), .Y(n4465) );
  OAI211X1 U422 ( .A0(n1244), .A1(n1313), .B0(n419), .C0(n3284), .Y(n4466) );
  OAI211X1 U423 ( .A0(n408), .A1(n953), .B0(n419), .C0(n3285), .Y(n4468) );
  OAI211X1 U424 ( .A0(n409), .A1(n1308), .B0(n419), .C0(n3286), .Y(n4473) );
  OAI211X1 U425 ( .A0(n412), .A1(n1331), .B0(n419), .C0(n3296), .Y(n4491) );
  OAI211X1 U426 ( .A0(n406), .A1(n1330), .B0(n419), .C0(n3297), .Y(n4492) );
  OAI211X1 U427 ( .A0(n1244), .A1(n1329), .B0(n419), .C0(n3298), .Y(n4493) );
  OAI211X1 U428 ( .A0(n408), .A1(n1388), .B0(n419), .C0(n3195), .Y(n4364) );
  NAND2X4 U429 ( .A(N956), .B(n807), .Y(n729) );
  INVXL U430 ( .A(n142), .Y(n206) );
  CLKINVX3 U431 ( .A(n206), .Y(n207) );
  OAI2BB1X4 U432 ( .A0N(SHA256_result[211]), .A1N(n305), .B0(n1064), .Y(
        f2_ABC_32[19]) );
  OAI21X4 U433 ( .A0(SHA256_result[211]), .A1(n305), .B0(SHA256_result[179]), 
        .Y(n1064) );
  OAI211X2 U434 ( .A0(n330), .A1(n731), .B0(n729), .C0(n730), .Y(n4551) );
  OAI211X1 U435 ( .A0(n1227), .A1(n26), .B0(n1014), .C0(n1013), .Y(n4683) );
  OAI211X1 U436 ( .A0(n1318), .A1(n22), .B0(n923), .C0(n922), .Y(n4649) );
  OAI211X1 U437 ( .A0(n1309), .A1(n22), .B0(n962), .C0(n961), .Y(n4662) );
  OAI211X1 U438 ( .A0(n1229), .A1(n25), .B0(n1010), .C0(n1009), .Y(n4681) );
  OAI211X1 U439 ( .A0(n1323), .A1(n24), .B0(n913), .C0(n912), .Y(n4644) );
  OAI211X1 U440 ( .A0(n1233), .A1(n21), .B0(n1002), .C0(n1001), .Y(n4677) );
  OAI211X1 U441 ( .A0(n1230), .A1(n28), .B0(n1008), .C0(n1007), .Y(n4680) );
  OAI211X1 U442 ( .A0(n1228), .A1(n24), .B0(n1012), .C0(n1011), .Y(n4682) );
  OAI211X1 U443 ( .A0(n1235), .A1(n26), .B0(n903), .C0(n902), .Y(n4639) );
  OAI211X1 U444 ( .A0(n1234), .A1(n25), .B0(n905), .C0(n904), .Y(n4640) );
  NAND2X4 U445 ( .A(n726), .B(n725), .Y(n4549) );
  NAND2X4 U446 ( .A(n812), .B(n816), .Y(n247) );
  NAND2X4 U447 ( .A(N964), .B(n807), .Y(n235) );
  OAI21X4 U448 ( .A0(SHA256_result[213]), .A1(n303), .B0(SHA256_result[181]), 
        .Y(n1062) );
  OAI2BB1X4 U449 ( .A0N(SHA256_result[213]), .A1N(n303), .B0(n1062), .Y(
        f2_ABC_32[21]) );
  NAND4X4 U450 ( .A(n707), .B(n708), .C(n802), .D(n706), .Y(n4542) );
  NAND2X4 U451 ( .A(N965), .B(n807), .Y(n707) );
  OAI2BB1X4 U452 ( .A0N(SHA256_result[214]), .A1N(n302), .B0(n1061), .Y(
        f2_ABC_32[22]) );
  OAI21X4 U453 ( .A0(n302), .A1(SHA256_result[214]), .B0(SHA256_result[182]), 
        .Y(n1061) );
  OAI2BB1X4 U454 ( .A0N(SHA256_result[215]), .A1N(n301), .B0(n1060), .Y(
        f2_ABC_32[23]) );
  OAI21X4 U455 ( .A0(n301), .A1(SHA256_result[215]), .B0(SHA256_result[183]), 
        .Y(n1060) );
  OAI2BB1X4 U456 ( .A0N(SHA256_result[210]), .A1N(n306), .B0(n1065), .Y(
        f2_ABC_32[18]) );
  NAND2X1 U457 ( .A(n247), .B(SHA256_result[176]), .Y(n924) );
  OAI2BB1X4 U458 ( .A0N(SHA256_result[212]), .A1N(n304), .B0(n1063), .Y(
        f2_ABC_32[20]) );
  NAND3BX4 U459 ( .AN(n810), .B(n450), .C(n441), .Y(n795) );
  INVX2 U460 ( .A(n795), .Y(n339) );
  INVX2 U461 ( .A(n795), .Y(n338) );
  INVX2 U462 ( .A(n795), .Y(n337) );
  NOR2X2 U463 ( .A(n435), .B(n318), .Y(n259) );
  NOR2X1 U464 ( .A(n2906), .B(n426), .Y(n258) );
  OAI21X4 U465 ( .A0(SHA256_result[208]), .A1(n308), .B0(SHA256_result[176]), 
        .Y(n1067) );
  OAI2BB1X4 U466 ( .A0N(SHA256_result[208]), .A1N(n308), .B0(n1067), .Y(
        f2_ABC_32[16]) );
  NAND2X4 U467 ( .A(N966), .B(n807), .Y(n214) );
  AND2X2 U468 ( .A(n90), .B(n323), .Y(n226) );
  NOR2X2 U469 ( .A(n1302), .B(n434), .Y(n4012) );
  INVX1 U470 ( .A(n4227), .Y(n1296) );
  BUFX12 U471 ( .A(SHA256_result[225]), .Y(n316) );
  AOI21XL U472 ( .A0(next_E[31]), .A1(n338), .B0(n805), .Y(n806) );
  OAI2BB1X4 U473 ( .A0N(SHA256_result[193]), .A1N(n316), .B0(n1082), .Y(
        f2_ABC_32[1]) );
  NAND2X1 U474 ( .A(n322), .B(SHA256_result[29]), .Y(n454) );
  NAND2X2 U475 ( .A(N872), .B(n286), .Y(n444) );
  OAI21X1 U476 ( .A0(n1403), .A1(n335), .B0(n446), .Y(n4283) );
  BUFX8 U477 ( .A(SHA256_result[243]), .Y(n305) );
  OAI211X1 U478 ( .A0(n331), .A1(n152), .B0(n660), .C0(n659), .Y(n4436) );
  OAI211X1 U479 ( .A0(n335), .A1(n784), .B0(n672), .C0(n671), .Y(n4440) );
  OAI211X1 U480 ( .A0(n335), .A1(n788), .B0(n674), .C0(n673), .Y(n4441) );
  OAI211X1 U481 ( .A0(n330), .A1(n148), .B0(n666), .C0(n665), .Y(n4438) );
  OAI211X1 U482 ( .A0(n332), .A1(n156), .B0(n677), .C0(n676), .Y(n4442) );
  OAI211X1 U483 ( .A0(n330), .A1(n768), .B0(n658), .C0(n657), .Y(n4435) );
  OAI211X1 U484 ( .A0(n333), .A1(n135), .B0(n663), .C0(n662), .Y(n4437) );
  OAI211X1 U485 ( .A0(n334), .A1(n780), .B0(n670), .C0(n669), .Y(n4439) );
  OAI2BB1X4 U486 ( .A0N(n99), .A1N(n221), .B0(n1080), .Y(f2_ABC_32[3]) );
  OAI21X4 U487 ( .A0(n221), .A1(n99), .B0(SHA256_result[163]), .Y(n1080) );
  INVX1 U488 ( .A(n237), .Y(n239) );
  INVXL U489 ( .A(n288), .Y(n397) );
  INVX1 U490 ( .A(n3954), .Y(n1298) );
  INVX1 U491 ( .A(n4088), .Y(n1257) );
  MXI2XL U492 ( .A(n885), .B(n967), .S0(n437), .Y(mux1[2]) );
  AOI21XL U493 ( .A0(n292), .A1(n341), .B0(n329), .Y(n781) );
  NAND2X1 U494 ( .A(N941), .B(n807), .Y(n782) );
  AOI21XL U495 ( .A0(n150), .A1(n341), .B0(n329), .Y(n777) );
  INVX1 U496 ( .A(n428), .Y(n426) );
  AOI21XL U497 ( .A0(n257), .A1(n286), .B0(n3950), .Y(n4179) );
  MX2X1 U498 ( .A(SHA256_result[139]), .B(SHA256_result[171]), .S0(n437), .Y(
        mux1[11]) );
  OAI211XL U499 ( .A0(n333), .A1(n796), .B0(n680), .C0(n679), .Y(n4443) );
  INVX1 U500 ( .A(SHA256_result[128]), .Y(n892) );
  MX2X1 U501 ( .A(SHA256_result[140]), .B(SHA256_result[172]), .S0(n437), .Y(
        mux1[12]) );
  AOI21XL U502 ( .A0(n344), .A1(SHA256_result[8]), .B0(n326), .Y(n504) );
  NAND2XL U503 ( .A(n1291), .B(n1276), .Y(n4113) );
  NAND2XL U504 ( .A(n1223), .B(n286), .Y(n442) );
  NOR2BX1 U505 ( .AN(n3564), .B(n815), .Y(n449) );
  INVX1 U506 ( .A(n405), .Y(n402) );
  INVX1 U507 ( .A(n405), .Y(n404) );
  NAND4XL U508 ( .A(n3999), .B(n4104), .C(n1291), .D(n3971), .Y(n4100) );
  NAND4XL U509 ( .A(n4184), .B(n4093), .C(n1291), .D(n1295), .Y(n4212) );
  NAND3XL U510 ( .A(n4151), .B(n4093), .C(n3958), .Y(n4237) );
  NAND2X1 U511 ( .A(N1081), .B(n357), .Y(n1134) );
  NAND4X1 U512 ( .A(n1135), .B(n1134), .C(n382), .D(n1133), .Y(n4748) );
  NAND3BX1 U513 ( .AN(n1179), .B(n382), .C(n1178), .Y(n4759) );
  OR2X2 U514 ( .A(n324), .B(n137), .Y(n250) );
  NAND2X1 U515 ( .A(next_A[13]), .B(n30), .Y(n1144) );
  MXI2X1 U516 ( .A(n887), .B(n969), .S0(n437), .Y(mux1[1]) );
  MXI2X1 U517 ( .A(n892), .B(n973), .S0(n437), .Y(mux1[0]) );
  OR2X2 U518 ( .A(n324), .B(n768), .Y(n254) );
  INVX4 U519 ( .A(n4159), .Y(n1295) );
  NOR3XL U520 ( .A(n4158), .B(n4137), .C(n4159), .Y(n4153) );
  AOI211XL U521 ( .A0(n3990), .A1(n425), .B0(n4136), .C0(n4120), .Y(n4135) );
  AOI211XL U522 ( .A0(n4024), .A1(n429), .B0(n4163), .C0(n1250), .Y(n4162) );
  NOR4XL U523 ( .A(n4066), .B(n3990), .C(n4244), .D(n4245), .Y(n4243) );
  NAND3BXL U524 ( .AN(n4074), .B(n1278), .C(n4094), .Y(n4144) );
  AOI2BB1XL U525 ( .A0N(n3989), .A1N(n3990), .B0(n426), .Y(n3987) );
  CLKINVX8 U526 ( .A(n4107), .Y(n1262) );
  OAI21XL U527 ( .A0(first_block_core), .A1(n448), .B0(n3564), .Y(n443) );
  OAI2BB1XL U528 ( .A0N(n447), .A1N(n440), .B0(n1221), .Y(n810) );
  NAND2XL U529 ( .A(n3964), .B(n258), .Y(n4019) );
  NOR2XL U530 ( .A(n259), .B(n260), .Y(n3948) );
  AOI22XL U531 ( .A0(n3745), .A1(n307), .B0(n3746), .B1(n303), .Y(n3854) );
  AOI22XL U532 ( .A0(n3745), .A1(n306), .B0(n3746), .B1(n302), .Y(n3812) );
  AOI22XL U533 ( .A0(n3745), .A1(n305), .B0(n3746), .B1(n301), .Y(n3738) );
  AND3X1 U534 ( .A(n259), .B(n4026), .C(n4016), .Y(n4028) );
  OAI211X1 U535 ( .A0(n1205), .A1(n21), .B0(n1049), .C0(n1048), .Y(n4698) );
  AOI21XL U536 ( .A0(n399), .A1(SHA256_result[157]), .B0(n387), .Y(n817) );
  NAND2XL U537 ( .A(n247), .B(SHA256_result[180]), .Y(n916) );
  OAI211X1 U538 ( .A0(n331), .A1(n739), .B0(n638), .C0(n637), .Y(n4427) );
  OAI211X1 U539 ( .A0(n332), .A1(n170), .B0(n644), .C0(n643), .Y(n4430) );
  OAI211X1 U540 ( .A0(n333), .A1(n91), .B0(n623), .C0(n622), .Y(n4420) );
  OAI211X1 U541 ( .A0(n335), .A1(n722), .B0(n625), .C0(n624), .Y(n4421) );
  NAND2X1 U542 ( .A(SHA256_result[6]), .B(n322), .Y(n510) );
  OAI2BB2X1 U543 ( .B0(n420), .B1(n1371), .A0N(H5[15]), .A1N(n205), .Y(n4332)
         );
  OAI2BB2X1 U544 ( .B0(n420), .B1(n1316), .A0N(H1[14]), .A1N(n205), .Y(n4461)
         );
  OAI2BB2X1 U545 ( .B0(n420), .B1(n1314), .A0N(H1[12]), .A1N(n205), .Y(n4463)
         );
  OAI2BB2X1 U546 ( .B0(n420), .B1(n1312), .A0N(H1[8]), .A1N(n205), .Y(n4467)
         );
  OAI2BB2X1 U547 ( .B0(n420), .B1(n1311), .A0N(H1[6]), .A1N(n205), .Y(n4469)
         );
  OAI2BB2X1 U548 ( .B0(n420), .B1(n1310), .A0N(H1[5]), .A1N(n205), .Y(n4470)
         );
  OAI2BB2X1 U549 ( .B0(n420), .B1(n1309), .A0N(H1[4]), .A1N(n205), .Y(n4471)
         );
  OAI2BB2X1 U550 ( .B0(n420), .B1(n98), .A0N(H1[3]), .A1N(n205), .Y(n4472) );
  OAI2BB2X1 U551 ( .B0(n420), .B1(n1307), .A0N(H1[1]), .A1N(n205), .Y(n4474)
         );
  OAI2BB2X1 U552 ( .B0(n420), .B1(n1415), .A0N(H7[18]), .A1N(n205), .Y(n4265)
         );
  OAI2BB2X1 U553 ( .B0(n420), .B1(n1414), .A0N(H7[17]), .A1N(n205), .Y(n4266)
         );
  OAI2BB2X1 U554 ( .B0(n420), .B1(n1413), .A0N(H7[16]), .A1N(n205), .Y(n4267)
         );
  OAI2BB2X1 U555 ( .B0(n420), .B1(n1410), .A0N(H7[13]), .A1N(n205), .Y(n4270)
         );
  OAI2BB2X1 U556 ( .B0(n420), .B1(n1409), .A0N(H7[12]), .A1N(n205), .Y(n4271)
         );
  OAI2BB2X1 U557 ( .B0(n420), .B1(n1406), .A0N(H7[9]), .A1N(n205), .Y(n4274)
         );
  OAI2BB2X1 U558 ( .B0(n420), .B1(n1404), .A0N(H7[7]), .A1N(n205), .Y(n4276)
         );
  OAI2BB2X1 U559 ( .B0(n420), .B1(n1366), .A0N(H3[30]), .A1N(n205), .Y(n4572)
         );
  OAI2BB2X1 U560 ( .B0(n420), .B1(n1364), .A0N(H3[28]), .A1N(n205), .Y(n4574)
         );
  OAI2BB2X1 U561 ( .B0(n420), .B1(n1363), .A0N(H3[27]), .A1N(n205), .Y(n4575)
         );
  OAI2BB2X1 U562 ( .B0(n420), .B1(n1361), .A0N(H3[25]), .A1N(n205), .Y(n4577)
         );
  OAI2BB2X1 U563 ( .B0(n420), .B1(n1359), .A0N(H3[23]), .A1N(n205), .Y(n4579)
         );
  OAI2BB2X1 U564 ( .B0(n420), .B1(n1357), .A0N(H3[21]), .A1N(n205), .Y(n4581)
         );
  OAI2BB2X1 U565 ( .B0(n420), .B1(n1356), .A0N(H3[20]), .A1N(n205), .Y(n4582)
         );
  OAI2BB2X1 U566 ( .B0(n420), .B1(n1347), .A0N(H3[11]), .A1N(n205), .Y(n4591)
         );
  OAI2BB2X1 U567 ( .B0(n420), .B1(n1233), .A0N(H0[21]), .A1N(n205), .Y(n4712)
         );
  OAI2BB2X1 U568 ( .B0(n420), .B1(n1232), .A0N(H0[20]), .A1N(n205), .Y(n4713)
         );
  OAI2BB2X1 U569 ( .B0(n420), .B1(n1230), .A0N(H0[18]), .A1N(n205), .Y(n4715)
         );
  OAI2BB2X1 U570 ( .B0(n420), .B1(n1229), .A0N(H0[17]), .A1N(n205), .Y(n4716)
         );
  AOI21XL U571 ( .A0(n399), .A1(SHA256_result[174]), .B0(n385), .Y(n929) );
  NAND2XL U572 ( .A(H6[28]), .B(n205), .Y(n3187) );
  NAND2XL U573 ( .A(H6[27]), .B(n205), .Y(n3188) );
  NAND2XL U574 ( .A(H6[25]), .B(n205), .Y(n3190) );
  NAND2XL U575 ( .A(H5[25]), .B(n205), .Y(n3177) );
  NAND2XL U576 ( .A(H1[25]), .B(n205), .Y(n3273) );
  NAND2XL U577 ( .A(H1[24]), .B(n205), .Y(n3274) );
  NAND2XL U578 ( .A(H4[18]), .B(n205), .Y(n3310) );
  OAI211X1 U579 ( .A0(n335), .A1(n125), .B0(n652), .C0(n651), .Y(n4433) );
  NAND2X1 U580 ( .A(n336), .B(SHA256_result[92]), .Y(n534) );
  CLKBUFX8 U581 ( .A(SHA256_result[240]), .Y(n308) );
  NAND2XL U582 ( .A(H5[27]), .B(n205), .Y(n3176) );
  NAND2XL U583 ( .A(H5[28]), .B(n205), .Y(n3175) );
  NOR2X1 U584 ( .A(n2925), .B(n434), .Y(n260) );
  NOR2XL U585 ( .A(n2938), .B(n426), .Y(n4014) );
  AOI211XL U586 ( .A0(n249), .A1(n286), .B0(n4032), .C0(n1222), .Y(n4157) );
  AND4X1 U587 ( .A(n3943), .B(n1260), .C(n1281), .D(n1295), .Y(n3941) );
  MX2XL U588 ( .A(SHA256_result[13]), .B(SHA256_result[45]), .S0(
        mux_control_0_), .Y(mux2[13]) );
  MX2XL U589 ( .A(SHA256_result[12]), .B(SHA256_result[44]), .S0(
        mux_control_0_), .Y(mux2[12]) );
  INVX1 U590 ( .A(SHA256_result[130]), .Y(n885) );
  NOR2X4 U591 ( .A(n1246), .B(n431), .Y(n3963) );
  INVXL U592 ( .A(n249), .Y(n1305) );
  NAND2XL U593 ( .A(n249), .B(n423), .Y(n3992) );
  NOR2X4 U594 ( .A(n318), .B(round[5]), .Y(n249) );
  INVXL U595 ( .A(n386), .Y(n382) );
  INVXL U596 ( .A(n385), .Y(n379) );
  INVXL U597 ( .A(n385), .Y(n378) );
  INVXL U598 ( .A(n288), .Y(n395) );
  INVXL U599 ( .A(n751), .Y(n324) );
  INVXL U600 ( .A(n288), .Y(n394) );
  INVXL U601 ( .A(n288), .Y(n391) );
  INVXL U602 ( .A(n288), .Y(n392) );
  INVXL U603 ( .A(n288), .Y(n393) );
  INVXL U604 ( .A(n288), .Y(n398) );
  NAND2BXL U605 ( .AN(n4075), .B(n1296), .Y(n4073) );
  NAND2XL U606 ( .A(n247), .B(SHA256_result[215]), .Y(n996) );
  NAND2XL U607 ( .A(n247), .B(SHA256_result[212]), .Y(n1003) );
  NAND2BXL U608 ( .AN(n810), .B(n816), .Y(n1200) );
  NAND3BXL U609 ( .AN(n815), .B(n816), .C(n3564), .Y(n1201) );
  NAND2XL U610 ( .A(n449), .B(n450), .Y(n800) );
  OR2XL U611 ( .A(n180), .B(n152), .Y(n248) );
  NOR2XL U612 ( .A(n1296), .B(n425), .Y(n3988) );
  AOI211XL U613 ( .A0(n427), .A1(n3955), .B0(n4043), .C0(n4072), .Y(n4240) );
  NAND2XL U614 ( .A(n1296), .B(n1259), .Y(n4226) );
  NOR2XL U615 ( .A(n1251), .B(n1303), .Y(n4009) );
  NOR2XL U616 ( .A(n426), .B(n1279), .Y(n4025) );
  NAND2XL U617 ( .A(n4012), .B(n4103), .Y(n4104) );
  NOR2XL U618 ( .A(n1302), .B(n431), .Y(n4030) );
  OAI211XL U619 ( .A0(n425), .A1(n1302), .B0(n1257), .C0(n1276), .Y(n4231) );
  AOI21XL U620 ( .A0(n1301), .A1(n3958), .B0(n808), .Y(n4001) );
  AOI22XL U621 ( .A0(n430), .A1(n286), .B0(n431), .B1(n3960), .Y(n4082) );
  NOR2XL U622 ( .A(n1302), .B(n1282), .Y(n3961) );
  NOR2XL U623 ( .A(n4026), .B(n1302), .Y(n3998) );
  AOI21XL U624 ( .A0(n1305), .A1(n3958), .B0(n1251), .Y(n4145) );
  AOI21XL U625 ( .A0(n4082), .A1(n1251), .B0(n1306), .Y(n4080) );
  OAI2BB1XL U626 ( .A0N(n3944), .A1N(n4083), .B0(n1279), .Y(n3949) );
  NAND2XL U627 ( .A(n294), .B(n399), .Y(n1087) );
  NAND2XL U628 ( .A(next_A[30]), .B(n30), .Y(n1089) );
  NAND2XL U629 ( .A(next_A[27]), .B(n30), .Y(n1101) );
  NAND2XL U630 ( .A(n297), .B(n399), .Y(n1099) );
  MXI2XL U631 ( .A(n876), .B(n960), .S0(n437), .Y(mux1[4]) );
  MXI2XL U632 ( .A(n880), .B(n964), .S0(n437), .Y(mux1[3]) );
  INVXL U633 ( .A(next_A[3]), .Y(n1187) );
  INVXL U634 ( .A(n247), .Y(n352) );
  AOI21XL U635 ( .A0(n343), .A1(n291), .B0(n329), .Y(n733) );
  INVXL U636 ( .A(next_E[3]), .Y(n787) );
  NAND2XL U637 ( .A(N939), .B(n807), .Y(n790) );
  INVXL U638 ( .A(next_E[1]), .Y(n794) );
  NAND3X4 U639 ( .A(n250), .B(n759), .C(n758), .Y(n4559) );
  NAND2XL U640 ( .A(n399), .B(n305), .Y(n1126) );
  NAND2XL U641 ( .A(N1084), .B(n357), .Y(n1127) );
  NAND2XL U642 ( .A(n399), .B(n309), .Y(n1136) );
  NAND2XL U643 ( .A(n399), .B(n310), .Y(n1139) );
  NAND2XL U644 ( .A(n295), .B(n399), .Y(n1091) );
  NAND2XL U645 ( .A(next_A[29]), .B(n30), .Y(n1093) );
  NAND2XL U646 ( .A(n299), .B(n399), .Y(n1107) );
  OR2X2 U647 ( .A(n324), .B(n125), .Y(n251) );
  OR2X2 U648 ( .A(n324), .B(n170), .Y(n252) );
  NAND2XL U649 ( .A(n29), .B(next_A[17]), .Y(n1131) );
  NAND2BXL U650 ( .AN(n23), .B(next_A[28]), .Y(n1096) );
  NAND2BXL U651 ( .AN(n21), .B(next_A[24]), .Y(n1112) );
  AOI22XL U652 ( .A0(N1089), .A1(n353), .B0(n300), .B1(n247), .Y(n1113) );
  NAND2BXL U653 ( .AN(n24), .B(next_A[20]), .Y(n1124) );
  AOI22XL U654 ( .A0(N1085), .A1(n353), .B0(n247), .B1(n304), .Y(n1125) );
  MXI2XL U655 ( .A(n870), .B(n954), .S0(n437), .Y(mux1[6]) );
  MXI2XL U656 ( .A(n867), .B(n951), .S0(n437), .Y(mux1[7]) );
  MXI2XL U657 ( .A(n872), .B(n957), .S0(n437), .Y(mux1[5]) );
  NOR2XL U658 ( .A(n1300), .B(n2946), .Y(n4004) );
  NOR2XL U659 ( .A(n798), .B(n797), .Y(n799) );
  NAND3XL U660 ( .A(n803), .B(n802), .C(n801), .Y(n4570) );
  NAND2XL U661 ( .A(next_E[0]), .B(n337), .Y(n803) );
  NAND2XL U662 ( .A(n312), .B(n399), .Y(n1161) );
  NAND2XL U663 ( .A(n313), .B(n399), .Y(n1173) );
  INVXL U664 ( .A(next_A[6]), .Y(n1172) );
  NAND2XL U665 ( .A(n315), .B(n399), .Y(n1191) );
  NAND2XL U666 ( .A(n314), .B(n399), .Y(n1178) );
  NAND2XL U667 ( .A(n316), .B(n399), .Y(n1196) );
  INVXL U668 ( .A(next_A[1]), .Y(n1195) );
  NAND2XL U669 ( .A(n317), .B(n399), .Y(n1203) );
  NAND2XL U670 ( .A(N1065), .B(n355), .Y(n1202) );
  NAND4XL U671 ( .A(n766), .B(n765), .C(n802), .D(n764), .Y(n4561) );
  NAND2XL U672 ( .A(n399), .B(SHA256_result[237]), .Y(n1142) );
  NAND2XL U673 ( .A(n399), .B(n308), .Y(n1133) );
  NAND3X1 U674 ( .A(n254), .B(n770), .C(n769), .Y(n4562) );
  AOI21XL U675 ( .A0(n136), .A1(n341), .B0(n329), .Y(n774) );
  MXI2XL U676 ( .A(n862), .B(n947), .S0(n437), .Y(mux1[8]) );
  MXI2XL U677 ( .A(n860), .B(n944), .S0(n437), .Y(mux1[9]) );
  MXI2XL U678 ( .A(n855), .B(n941), .S0(n437), .Y(mux1[10]) );
  OR2X4 U679 ( .A(n320), .B(n432), .Y(n255) );
  NOR2XL U680 ( .A(n426), .B(n320), .Y(n4055) );
  AOI31XL U681 ( .A0(n3502), .A1(n3578), .A2(n1245), .B0(n1243), .Y(n4250) );
  CLKINVX2 U682 ( .A(n433), .Y(n431) );
  NOR2XL U683 ( .A(round[0]), .B(n320), .Y(n4103) );
  NAND2XL U684 ( .A(n318), .B(n258), .Y(n3958) );
  AOI22XL U685 ( .A0(n1265), .A1(n286), .B0(n3960), .B1(n259), .Y(n4020) );
  NOR2XL U686 ( .A(n809), .B(n320), .Y(n4248) );
  OAI22XL U687 ( .A0(n3502), .A1(n1243), .B0(n3501), .B1(n436), .Y(n4700) );
  OAI22XL U688 ( .A0(n3378), .A1(n1243), .B0(n3501), .B1(n439), .Y(n4701) );
  AOI221XL U689 ( .A0(n4041), .A1(n434), .B0(n253), .B1(n258), .C0(n4155), .Y(
        n4154) );
  NOR3XL U690 ( .A(n4164), .B(n4057), .C(n4074), .Y(n4161) );
  AOI22XL U691 ( .A0(n260), .A1(n4026), .B0(n253), .B1(n4014), .Y(n4202) );
  NOR3XL U692 ( .A(n3961), .B(n1262), .C(n4056), .Y(n4168) );
  AOI222XL U693 ( .A0(n253), .A1(n4140), .B0(n4059), .B1(n1223), .C0(n4132), 
        .C1(n422), .Y(n4133) );
  AOI211XL U694 ( .A0(n4059), .A1(n260), .B0(n4044), .C0(n1262), .Y(n4045) );
  NOR4BXL U695 ( .AN(n3971), .B(n4057), .C(n3988), .D(n4058), .Y(n4046) );
  AOI211XL U696 ( .A0(n3986), .A1(n422), .B0(n3987), .C0(n3988), .Y(n3980) );
  AOI31XL U697 ( .A0(n429), .A1(n427), .A2(n4011), .B0(n4123), .Y(n4115) );
  AOI211XL U698 ( .A0(n4118), .A1(n286), .B0(n4119), .C0(n4120), .Y(n4117) );
  AOI211XL U699 ( .A0(n4063), .A1(n320), .B0(n4064), .C0(n4065), .Y(n4062) );
  AOI21XL U700 ( .A0(n429), .A1(n4073), .B0(n4074), .Y(n4060) );
  AOI22XL U701 ( .A0(n3973), .A1(n259), .B0(n434), .B1(n4042), .Y(n4034) );
  AOI22XL U702 ( .A0(n4043), .A1(n318), .B0(n4044), .B1(n320), .Y(n4033) );
  AOI211XL U703 ( .A0(n4036), .A1(n286), .B0(n4037), .C0(n4038), .Y(n4035) );
  NOR2XL U704 ( .A(n1277), .B(n320), .Y(n4058) );
  NAND2XL U705 ( .A(n260), .B(n286), .Y(n4094) );
  AOI211XL U706 ( .A0(n260), .A1(n319), .B0(n259), .C0(n3960), .Y(n3957) );
  NOR2XL U707 ( .A(n2946), .B(n4107), .Y(n4072) );
  NOR2XL U708 ( .A(n1251), .B(n318), .Y(n4039) );
  NOR2XL U709 ( .A(n1275), .B(n320), .Y(n4150) );
  AOI222XL U710 ( .A0(n4055), .A1(n1223), .B0(n4132), .B1(n429), .C0(n260), 
        .C1(n4014), .Y(n4241) );
  AND4X1 U711 ( .A(n4183), .B(n1279), .C(n1273), .D(n4184), .Y(n4182) );
  AOI22XL U712 ( .A0(n4044), .A1(n422), .B0(n4159), .B1(n2946), .Y(n4174) );
  AOI222XL U713 ( .A0(n4012), .A1(n4055), .B0(n3973), .B1(n257), .C0(n1224), 
        .C1(n4140), .Y(n4175) );
  AOI222XL U714 ( .A0(n4012), .A1(n422), .B0(n4013), .B1(n434), .C0(n260), 
        .C1(n4014), .Y(n4006) );
  AOI211XL U715 ( .A0(n3973), .A1(n249), .B0(n3975), .C0(n3976), .Y(n3967) );
  AOI21XL U716 ( .A0(n1289), .A1(n429), .B0(n3978), .Y(n3966) );
  AOI31XL U717 ( .A0(n319), .A1(n286), .A2(n434), .B0(n1264), .Y(n3970) );
  NAND2BXL U718 ( .AN(n2946), .B(n2947), .Y(n808) );
  NAND4XL U719 ( .A(n4104), .B(n3985), .C(n1278), .D(n1246), .Y(n4244) );
  NOR2XL U720 ( .A(n2947), .B(n319), .Y(n3960) );
  INVX1 U721 ( .A(n266), .Y(n417) );
  NAND2XL U722 ( .A(n257), .B(n258), .Y(n3999) );
  INVX1 U723 ( .A(n266), .Y(n418) );
  NAND2XL U724 ( .A(n253), .B(n4016), .Y(n4010) );
  NOR3XL U725 ( .A(n2946), .B(n431), .C(n4086), .Y(n3969) );
  NOR2XL U726 ( .A(n4086), .B(n320), .Y(n3997) );
  AOI21XL U727 ( .A0(n3985), .A1(n4124), .B0(n427), .Y(n4123) );
  AOI2BB1XL U728 ( .A0N(n4011), .A1N(n3997), .B0(n429), .Y(n4218) );
  AOI21XL U729 ( .A0(n4124), .A1(n1283), .B0(n431), .Y(n4199) );
  AOI2BB1XL U730 ( .A0N(n257), .A1N(n3965), .B0(n1251), .Y(n3975) );
  AOI22XL U731 ( .A0(n3741), .A1(n316), .B0(n3742), .B1(n314), .Y(n3856) );
  AOI22XL U732 ( .A0(n3741), .A1(n315), .B0(n3742), .B1(n313), .Y(n3814) );
  AOI22XL U733 ( .A0(n3743), .A1(n15), .B0(n3744), .B1(n309), .Y(n3739) );
  AOI22XL U734 ( .A0(n3743), .A1(n311), .B0(n3744), .B1(n310), .Y(n3813) );
  AOI22XL U735 ( .A0(n3743), .A1(n312), .B0(n3744), .B1(SHA256_result[237]), 
        .Y(n3855) );
  INVX1 U736 ( .A(n320), .Y(n425) );
  NOR3XL U737 ( .A(n1280), .B(n434), .C(n432), .Y(n4138) );
  NAND2XL U738 ( .A(n3946), .B(n249), .Y(n4052) );
  INVXL U739 ( .A(n309), .Y(n1227) );
  INVXL U740 ( .A(SHA256_result[237]), .Y(n1225) );
  INVXL U741 ( .A(n317), .Y(n1205) );
  INVXL U742 ( .A(n292), .Y(n780) );
  INVXL U743 ( .A(n310), .Y(n1226) );
  INVXL U744 ( .A(n313), .Y(n1170) );
  INVXL U745 ( .A(n314), .Y(n1175) );
  INVXL U746 ( .A(n316), .Y(n1193) );
  INVXL U747 ( .A(n311), .Y(n1154) );
  INVXL U748 ( .A(n312), .Y(n1158) );
  INVXL U749 ( .A(n315), .Y(n1188) );
  INVXL U750 ( .A(SHA256_result[236]), .Y(n1146) );
  INVXL U751 ( .A(n15), .Y(n1151) );
  OAI211XL U752 ( .A0(n406), .A1(n1408), .B0(n419), .C0(n3128), .Y(n4272) );
  INVXL U753 ( .A(SHA256_result[11]), .Y(n1408) );
  NAND2XL U754 ( .A(H7[11]), .B(n205), .Y(n3128) );
  OAI211XL U755 ( .A0(n407), .A1(n1407), .B0(n419), .C0(n3129), .Y(n4273) );
  INVXL U756 ( .A(SHA256_result[10]), .Y(n1407) );
  NAND2XL U757 ( .A(H7[10]), .B(n205), .Y(n3129) );
  OAI211XL U758 ( .A0(n412), .A1(n1405), .B0(n419), .C0(n3130), .Y(n4275) );
  INVXL U759 ( .A(SHA256_result[8]), .Y(n1405) );
  NAND2XL U760 ( .A(H7[8]), .B(n205), .Y(n3130) );
  INVXL U761 ( .A(SHA256_result[60]), .Y(n1400) );
  INVXL U762 ( .A(SHA256_result[59]), .Y(n1399) );
  INVXL U763 ( .A(SHA256_result[57]), .Y(n1397) );
  NAND2XL U764 ( .A(H6[15]), .B(n205), .Y(n3195) );
  INVXL U765 ( .A(SHA256_result[92]), .Y(n1384) );
  INVXL U766 ( .A(SHA256_result[91]), .Y(n1383) );
  INVXL U767 ( .A(SHA256_result[89]), .Y(n1381) );
  INVXL U768 ( .A(n291), .Y(n1368) );
  OAI211XL U769 ( .A0(n407), .A1(n1351), .B0(n419), .C0(n3389), .Y(n4587) );
  NAND2XL U770 ( .A(H3[15]), .B(n205), .Y(n3389) );
  OAI211XL U771 ( .A0(n412), .A1(n1350), .B0(n419), .C0(n3390), .Y(n4588) );
  NAND2XL U772 ( .A(H3[14]), .B(n205), .Y(n3390) );
  OAI211XL U773 ( .A0(n407), .A1(n1349), .B0(n419), .C0(n3391), .Y(n4589) );
  INVXL U774 ( .A(SHA256_result[141]), .Y(n1349) );
  NAND2XL U775 ( .A(H3[13]), .B(n205), .Y(n3391) );
  OAI211XL U776 ( .A0(n410), .A1(n1348), .B0(n419), .C0(n3392), .Y(n4590) );
  NAND2XL U777 ( .A(H3[12]), .B(n205), .Y(n3392) );
  NAND2XL U778 ( .A(H2[15]), .B(n205), .Y(n3296) );
  NAND2XL U779 ( .A(H2[14]), .B(n205), .Y(n3297) );
  NAND2XL U780 ( .A(H2[13]), .B(n205), .Y(n3298) );
  INVXL U781 ( .A(SHA256_result[217]), .Y(n1326) );
  INVXL U782 ( .A(SHA256_result[216]), .Y(n1325) );
  NAND2XL U783 ( .A(H1[15]), .B(n205), .Y(n3280) );
  NAND2XL U784 ( .A(H1[13]), .B(n205), .Y(n3281) );
  NAND2XL U785 ( .A(H1[11]), .B(n205), .Y(n3282) );
  NAND2XL U786 ( .A(H1[10]), .B(n205), .Y(n3283) );
  NAND2XL U787 ( .A(H1[9]), .B(n205), .Y(n3284) );
  NAND2XL U788 ( .A(H1[7]), .B(n205), .Y(n3285) );
  NAND2XL U789 ( .A(H1[2]), .B(n205), .Y(n3286) );
  OAI211XL U790 ( .A0(n408), .A1(n97), .B0(n419), .C0(n3500), .Y(n4699) );
  NAND2XL U791 ( .A(H1[0]), .B(n205), .Y(n3500) );
  OAI21X4 U792 ( .A0(SHA256_result[193]), .A1(n316), .B0(SHA256_result[161]), 
        .Y(n1082) );
  NAND2XL U793 ( .A(H5[14]), .B(n205), .Y(n3181) );
  NAND2XL U794 ( .A(H5[13]), .B(n205), .Y(n3182) );
  NAND2XL U795 ( .A(H5[11]), .B(n205), .Y(n3183) );
  NAND2XL U796 ( .A(H5[7]), .B(n205), .Y(n3184) );
  NAND2XL U797 ( .A(H5[3]), .B(n205), .Y(n3185) );
  NAND2XL U798 ( .A(H5[2]), .B(n205), .Y(n3186) );
  NAND2XL U799 ( .A(H6[14]), .B(n205), .Y(n3196) );
  NAND2XL U800 ( .A(H6[12]), .B(n205), .Y(n3197) );
  NAND2XL U801 ( .A(H6[11]), .B(n205), .Y(n3198) );
  NAND2XL U802 ( .A(H6[8]), .B(n205), .Y(n3199) );
  NAND2XL U803 ( .A(H6[7]), .B(n205), .Y(n3200) );
  NAND2XL U804 ( .A(H6[5]), .B(n205), .Y(n3201) );
  NAND2XL U805 ( .A(H6[3]), .B(n205), .Y(n3202) );
  NAND2XL U806 ( .A(H6[1]), .B(n205), .Y(n3203) );
  NAND2XL U807 ( .A(H6[0]), .B(n205), .Y(n3204) );
  NAND2XL U808 ( .A(H7[1]), .B(n205), .Y(n521) );
  NAND2XL U809 ( .A(H6[13]), .B(n205), .Y(n571) );
  NAND2XL U810 ( .A(H6[10]), .B(n205), .Y(n578) );
  NAND2XL U811 ( .A(H6[9]), .B(n205), .Y(n581) );
  NAND2XL U812 ( .A(H6[6]), .B(n205), .Y(n588) );
  NAND2XL U813 ( .A(H6[4]), .B(n205), .Y(n593) );
  NAND2XL U814 ( .A(H6[2]), .B(n205), .Y(n598) );
  NAND2XL U815 ( .A(H5[12]), .B(n205), .Y(n645) );
  NAND2XL U816 ( .A(H5[10]), .B(n205), .Y(n650) );
  NAND2XL U817 ( .A(H5[9]), .B(n205), .Y(n653) );
  NAND2XL U818 ( .A(H5[8]), .B(n205), .Y(n656) );
  NAND2XL U819 ( .A(H5[6]), .B(n205), .Y(n661) );
  NAND2XL U820 ( .A(H5[5]), .B(n205), .Y(n664) );
  NAND2XL U821 ( .A(H5[4]), .B(n205), .Y(n667) );
  NAND2XL U822 ( .A(H5[1]), .B(n205), .Y(n675) );
  NAND2XL U823 ( .A(H5[0]), .B(n205), .Y(n678) );
  NAND2XL U824 ( .A(H3[9]), .B(n205), .Y(n859) );
  NAND2XL U825 ( .A(H3[7]), .B(n205), .Y(n866) );
  NAND2XL U826 ( .A(H3[6]), .B(n205), .Y(n869) );
  NAND2XL U827 ( .A(H3[2]), .B(n205), .Y(n884) );
  NAND2XL U828 ( .A(H3[0]), .B(n205), .Y(n891) );
  NAND2XL U829 ( .A(H2[11]), .B(n205), .Y(n936) );
  NAND2XL U830 ( .A(H2[10]), .B(n205), .Y(n940) );
  NAND2XL U831 ( .A(H2[7]), .B(n205), .Y(n950) );
  NAND2XL U832 ( .A(H2[3]), .B(n205), .Y(n963) );
  NAND2XL U833 ( .A(H2[2]), .B(n205), .Y(n966) );
  NAND2XL U834 ( .A(H2[0]), .B(n205), .Y(n972) );
  OAI211XL U835 ( .A0(n408), .A1(n1193), .B0(n3519), .C0(n419), .Y(n4732) );
  NAND2XL U836 ( .A(H0[1]), .B(n205), .Y(n3519) );
  NAND2XL U837 ( .A(H0[0]), .B(n205), .Y(n3576) );
  OAI211XL U838 ( .A0(n407), .A1(n855), .B0(n3393), .C0(n419), .Y(n4592) );
  NAND2XL U839 ( .A(H3[10]), .B(n205), .Y(n3393) );
  OAI211XL U840 ( .A0(n412), .A1(n862), .B0(n3394), .C0(n419), .Y(n4594) );
  NAND2XL U841 ( .A(H3[8]), .B(n205), .Y(n3394) );
  OAI211XL U842 ( .A0(n410), .A1(n872), .B0(n3395), .C0(n419), .Y(n4597) );
  NAND2XL U843 ( .A(H3[5]), .B(n205), .Y(n3395) );
  OAI211XL U844 ( .A0(n1244), .A1(n876), .B0(n3396), .C0(n419), .Y(n4598) );
  NAND2XL U845 ( .A(H3[4]), .B(n205), .Y(n3396) );
  OAI211XL U846 ( .A0(n406), .A1(n880), .B0(n3397), .C0(n419), .Y(n4599) );
  NAND2XL U847 ( .A(H3[3]), .B(n205), .Y(n3397) );
  OAI211XL U848 ( .A0(n407), .A1(n887), .B0(n3398), .C0(n419), .Y(n4601) );
  NAND2XL U849 ( .A(H3[1]), .B(n205), .Y(n3398) );
  OAI211XL U850 ( .A0(n410), .A1(n933), .B0(n3299), .C0(n419), .Y(n4494) );
  NAND2XL U851 ( .A(H2[12]), .B(n205), .Y(n3299) );
  OAI211XL U852 ( .A0(n408), .A1(n944), .B0(n3300), .C0(n419), .Y(n4497) );
  NAND2XL U853 ( .A(H2[9]), .B(n205), .Y(n3300) );
  OAI211XL U854 ( .A0(n410), .A1(n947), .B0(n3301), .C0(n419), .Y(n4498) );
  NAND2XL U855 ( .A(H2[8]), .B(n205), .Y(n3301) );
  OAI211XL U856 ( .A0(n412), .A1(n954), .B0(n3302), .C0(n419), .Y(n4500) );
  NAND2XL U857 ( .A(H2[6]), .B(n205), .Y(n3302) );
  OAI211XL U858 ( .A0(n410), .A1(n957), .B0(n3303), .C0(n419), .Y(n4501) );
  NAND2XL U859 ( .A(H2[5]), .B(n205), .Y(n3303) );
  OAI211XL U860 ( .A0(n407), .A1(n960), .B0(n3304), .C0(n419), .Y(n4502) );
  NAND2XL U861 ( .A(H2[4]), .B(n205), .Y(n3304) );
  NAND2XL U862 ( .A(H2[1]), .B(n205), .Y(n3305) );
  OAI211XL U863 ( .A0(n412), .A1(n1412), .B0(n419), .C0(n3126), .Y(n4268) );
  NAND2XL U864 ( .A(H7[15]), .B(n205), .Y(n3126) );
  OAI211XL U865 ( .A0(n411), .A1(n1411), .B0(n419), .C0(n3127), .Y(n4269) );
  NAND2XL U866 ( .A(H7[14]), .B(n205), .Y(n3127) );
  OAI211XL U867 ( .A0(n408), .A1(n113), .B0(n3306), .C0(n419), .Y(n4508) );
  OAI211XL U868 ( .A0(n1244), .A1(n705), .B0(n3307), .C0(n419), .Y(n4510) );
  OAI211XL U869 ( .A0(n409), .A1(n715), .B0(n3308), .C0(n419), .Y(n4514) );
  OAI211XL U870 ( .A0(n408), .A1(n746), .B0(n3312), .C0(n419), .Y(n4524) );
  OAI211XL U871 ( .A0(n409), .A1(n145), .B0(n3313), .C0(n419), .Y(n4526) );
  OAI211XL U872 ( .A0(n412), .A1(n1211), .B0(n3131), .C0(n419), .Y(n4279) );
  NAND2XL U873 ( .A(H7[4]), .B(n205), .Y(n3131) );
  OAI211XL U874 ( .A0(n407), .A1(n1213), .B0(n3132), .C0(n419), .Y(n4280) );
  NAND2XL U875 ( .A(H7[3]), .B(n205), .Y(n3132) );
  OAI211XL U876 ( .A0(n412), .A1(n1218), .B0(n3173), .C0(n419), .Y(n4315) );
  NAND2XL U877 ( .A(H7[0]), .B(n205), .Y(n3173) );
  INVXL U878 ( .A(SHA256_result[9]), .Y(n1406) );
  INVXL U879 ( .A(SHA256_result[7]), .Y(n1404) );
  INVXL U880 ( .A(SHA256_result[90]), .Y(n1382) );
  NAND2XL U881 ( .A(n247), .B(SHA256_result[139]), .Y(n853) );
  NAND2XL U882 ( .A(n247), .B(n86), .Y(n906) );
  NAND2XL U883 ( .A(n247), .B(SHA256_result[184]), .Y(n908) );
  NAND2XL U884 ( .A(n247), .B(SHA256_result[183]), .Y(n910) );
  INVXL U885 ( .A(SHA256_result[208]), .Y(n925) );
  NAND2XL U886 ( .A(n247), .B(SHA256_result[218]), .Y(n988) );
  NAND2XL U887 ( .A(n321), .B(SHA256_result[26]), .Y(n462) );
  NAND2XL U888 ( .A(n323), .B(SHA256_result[20]), .Y(n479) );
  NAND2XL U889 ( .A(n322), .B(SHA256_result[19]), .Y(n481) );
  NAND2XL U890 ( .A(n322), .B(SHA256_result[18]), .Y(n483) );
  NAND2XL U891 ( .A(n322), .B(SHA256_result[17]), .Y(n485) );
  NAND2XL U892 ( .A(n321), .B(SHA256_result[16]), .Y(n487) );
  NAND2XL U893 ( .A(n322), .B(SHA256_result[62]), .Y(n528) );
  NAND2XL U894 ( .A(n322), .B(SHA256_result[61]), .Y(n530) );
  OAI22XL U895 ( .A0(round[6]), .A1(n3580), .B0(n4251), .B1(n2878), .Y(n3574)
         );
  AOI22XL U896 ( .A0(n4103), .A1(n1222), .B0(n3963), .B1(n2946), .Y(n4251) );
  NAND2XL U897 ( .A(N886), .B(n807), .Y(n572) );
  OAI211X1 U898 ( .A0(n332), .A1(n689), .B0(n580), .C0(n579), .Y(n4401) );
  OAI211X1 U899 ( .A0(n332), .A1(n690), .B0(n583), .C0(n582), .Y(n4402) );
  NAND2XL U900 ( .A(SHA256_result[1]), .B(n323), .Y(n523) );
  NAND2XL U901 ( .A(N842), .B(n807), .Y(n522) );
  NAND2XL U902 ( .A(N849), .B(n807), .Y(n505) );
  NAND2XL U903 ( .A(N845), .B(n807), .Y(n515) );
  AOI21XL U904 ( .A0(SHA256_result[4]), .A1(n341), .B0(n326), .Y(n514) );
  NAND2XL U905 ( .A(N844), .B(n807), .Y(n517) );
  AOI21XL U906 ( .A0(SHA256_result[3]), .A1(n341), .B0(n326), .Y(n516) );
  NAND2XL U907 ( .A(N841), .B(n807), .Y(n525) );
  AOI21XL U908 ( .A0(n344), .A1(SHA256_result[14]), .B0(n329), .Y(n492) );
  NAND2XL U909 ( .A(n322), .B(SHA256_result[13]), .Y(n495) );
  NAND2XL U910 ( .A(n322), .B(SHA256_result[12]), .Y(n497) );
  NAND2XL U911 ( .A(N852), .B(n807), .Y(n499) );
  AOI21XL U912 ( .A0(n345), .A1(SHA256_result[11]), .B0(n328), .Y(n498) );
  NAND2XL U913 ( .A(N851), .B(n807), .Y(n501) );
  AOI21XL U914 ( .A0(n344), .A1(SHA256_result[10]), .B0(n328), .Y(n500) );
  NAND2XL U915 ( .A(N850), .B(n807), .Y(n502) );
  NAND2XL U916 ( .A(n322), .B(SHA256_result[9]), .Y(n503) );
  NAND2XL U917 ( .A(N848), .B(n807), .Y(n506) );
  NAND2XL U918 ( .A(n322), .B(SHA256_result[7]), .Y(n507) );
  NAND2XL U919 ( .A(N847), .B(n807), .Y(n509) );
  NAND2XL U920 ( .A(SHA256_result[5]), .B(n323), .Y(n513) );
  NAND2XL U921 ( .A(N846), .B(n807), .Y(n512) );
  NAND2XL U922 ( .A(N843), .B(n807), .Y(n519) );
  NAND2XL U923 ( .A(SHA256_result[2]), .B(n323), .Y(n520) );
  OAI21X4 U924 ( .A0(output_enable), .A1(inner_busy), .B0(n3114), .Y(n3577) );
  OAI211X1 U925 ( .A0(n333), .A1(n681), .B0(n570), .C0(n569), .Y(n4397) );
  OAI211X1 U926 ( .A0(n334), .A1(n687), .B0(n577), .C0(n576), .Y(n4400) );
  OAI211X1 U927 ( .A0(n332), .A1(n691), .B0(n585), .C0(n584), .Y(n4403) );
  NAND2XL U928 ( .A(N932), .B(n807), .Y(n615) );
  AOI21XL U929 ( .A0(n343), .A1(SHA256_result[91]), .B0(n328), .Y(n614) );
  OAI211XL U930 ( .A0(n332), .A1(n243), .B0(n619), .C0(n618), .Y(n4418) );
  NAND2XL U931 ( .A(N930), .B(n807), .Y(n619) );
  AOI21XL U932 ( .A0(n343), .A1(SHA256_result[89]), .B0(n328), .Y(n618) );
  OAI211XL U933 ( .A0(n334), .A1(n715), .B0(n621), .C0(n620), .Y(n4419) );
  NAND2XL U934 ( .A(N929), .B(n807), .Y(n621) );
  AOI21XL U935 ( .A0(n343), .A1(n31), .B0(n328), .Y(n620) );
  OAI211XL U936 ( .A0(n333), .A1(n705), .B0(n613), .C0(n612), .Y(n4415) );
  NAND2XL U937 ( .A(N933), .B(n807), .Y(n613) );
  AOI21XL U938 ( .A0(n343), .A1(SHA256_result[92]), .B0(n327), .Y(n612) );
  NAND2XL U939 ( .A(H7[6]), .B(n205), .Y(n508) );
  NAND2XL U940 ( .A(H7[5]), .B(n205), .Y(n511) );
  NAND2XL U941 ( .A(H7[2]), .B(n205), .Y(n518) );
  NAND2XL U942 ( .A(n103), .B(n345), .Y(n716) );
  OAI21X4 U943 ( .A0(SHA256_result[196]), .A1(SHA256_result[228]), .B0(
        SHA256_result[164]), .Y(n1079) );
  OAI21X4 U944 ( .A0(n315), .A1(SHA256_result[194]), .B0(SHA256_result[162]), 
        .Y(n1081) );
  NAND2XL U945 ( .A(n337), .B(n291), .Y(n634) );
  NAND2XL U946 ( .A(N896), .B(n807), .Y(n548) );
  NAND2XL U947 ( .A(N890), .B(n807), .Y(n561) );
  NAND2XL U948 ( .A(N889), .B(n807), .Y(n564) );
  NAND2XL U949 ( .A(N888), .B(n807), .Y(n567) );
  NAND2XL U950 ( .A(N936), .B(n807), .Y(n606) );
  AOI21XL U951 ( .A0(n343), .A1(SHA256_result[95]), .B0(n327), .Y(n605) );
  NAND2XL U952 ( .A(N901), .B(n807), .Y(n533) );
  AOI21XL U953 ( .A0(n344), .A1(SHA256_result[60]), .B0(n326), .Y(n532) );
  NAND2XL U954 ( .A(n338), .B(SHA256_result[91]), .Y(n537) );
  NAND2XL U955 ( .A(N900), .B(n807), .Y(n536) );
  NAND2XL U956 ( .A(n339), .B(SHA256_result[90]), .Y(n540) );
  NAND2XL U957 ( .A(N899), .B(n807), .Y(n539) );
  AOI21XL U958 ( .A0(n344), .A1(SHA256_result[58]), .B0(n326), .Y(n538) );
  NAND2XL U959 ( .A(n338), .B(SHA256_result[89]), .Y(n543) );
  NAND2XL U960 ( .A(N898), .B(n807), .Y(n542) );
  NAND2XL U961 ( .A(n338), .B(n31), .Y(n546) );
  NAND2XL U962 ( .A(N897), .B(n807), .Y(n545) );
  AOI21XL U963 ( .A0(n344), .A1(n119), .B0(n326), .Y(n544) );
  OAI2BB1XL U964 ( .A0N(n115), .A1N(n345), .B0(n802), .Y(n700) );
  CLKBUFX8 U965 ( .A(SHA256_result[246]), .Y(n302) );
  CLKBUFX8 U966 ( .A(SHA256_result[247]), .Y(n301) );
  NAND2XL U967 ( .A(N1040), .B(n356), .Y(n1032) );
  NAND2XL U968 ( .A(N1035), .B(n124), .Y(n1043) );
  OAI211XL U969 ( .A0(n26), .A1(n1090), .B0(n983), .C0(n982), .Y(n4669) );
  NAND2XL U970 ( .A(N1062), .B(n355), .Y(n983) );
  OAI211XL U971 ( .A0(n27), .A1(n1095), .B0(n985), .C0(n984), .Y(n4670) );
  NAND2XL U972 ( .A(N1061), .B(n355), .Y(n985) );
  OAI211XL U973 ( .A0(n26), .A1(n1098), .B0(n987), .C0(n986), .Y(n4671) );
  NAND2XL U974 ( .A(N1060), .B(n355), .Y(n987) );
  AOI21XL U975 ( .A0(n399), .A1(SHA256_result[219]), .B0(n389), .Y(n986) );
  MX2X4 U976 ( .A(n119), .B(n31), .S0(n102), .Y(f1_EFG_32[24]) );
  NAND2XL U977 ( .A(N1033), .B(n356), .Y(n1049) );
  NAND2XL U978 ( .A(N1010), .B(n355), .Y(n946) );
  NAND2XL U979 ( .A(N1005), .B(n355), .Y(n962) );
  AOI21XL U980 ( .A0(SHA256_result[164]), .A1(n399), .B0(n389), .Y(n961) );
  NAND2XL U981 ( .A(N1046), .B(n356), .Y(n1018) );
  NAND2XL U982 ( .A(N1050), .B(n356), .Y(n1010) );
  AOI21XL U983 ( .A0(SHA256_result[209]), .A1(n399), .B0(n390), .Y(n1009) );
  NAND2XL U984 ( .A(N1048), .B(n356), .Y(n1014) );
  NAND2XL U985 ( .A(N1013), .B(n355), .Y(n935) );
  NAND2XL U986 ( .A(N1009), .B(n355), .Y(n949) );
  NAND2XL U987 ( .A(N1007), .B(n355), .Y(n956) );
  NAND2XL U988 ( .A(N1006), .B(n355), .Y(n959) );
  AOI21XL U989 ( .A0(n399), .A1(SHA256_result[175]), .B0(n387), .Y(n927) );
  NAND2XL U990 ( .A(N1014), .B(n355), .Y(n932) );
  NAND2XL U991 ( .A(N1002), .B(n355), .Y(n971) );
  AOI21XL U992 ( .A0(SHA256_result[161]), .A1(n399), .B0(n389), .Y(n970) );
  OAI211XL U993 ( .A0(n332), .A1(n113), .B0(n609), .C0(n608), .Y(n4413) );
  NAND2XL U994 ( .A(n321), .B(SHA256_result[94]), .Y(n609) );
  NAND2XL U995 ( .A(n321), .B(SHA256_result[93]), .Y(n611) );
  OAI211XL U996 ( .A0(n332), .A1(n116), .B0(n617), .C0(n616), .Y(n4417) );
  NAND2XL U997 ( .A(N931), .B(n807), .Y(n616) );
  NAND2XL U998 ( .A(n321), .B(SHA256_result[90]), .Y(n617) );
  NAND2XL U999 ( .A(N995), .B(n355), .Y(n824) );
  OAI211XL U1000 ( .A0(n1329), .A1(n21), .B0(n850), .C0(n849), .Y(n4621) );
  NAND2XL U1001 ( .A(N982), .B(n354), .Y(n850) );
  AOI21XL U1002 ( .A0(n399), .A1(SHA256_result[141]), .B0(n390), .Y(n849) );
  OAI211XL U1003 ( .A0(n1328), .A1(n27), .B0(n895), .C0(n894), .Y(n4603) );
  OAI211XL U1004 ( .A0(n1237), .A1(n25), .B0(n899), .C0(n898), .Y(n4637) );
  OAI211XL U1005 ( .A0(n1236), .A1(n27), .B0(n901), .C0(n900), .Y(n4638) );
  NAND2XL U1006 ( .A(N1028), .B(n369), .Y(n903) );
  AOI21XL U1007 ( .A0(n399), .A1(SHA256_result[187]), .B0(n387), .Y(n902) );
  NAND2XL U1008 ( .A(N1027), .B(n370), .Y(n905) );
  AOI21XL U1009 ( .A0(n399), .A1(SHA256_result[186]), .B0(n387), .Y(n904) );
  NAND2XL U1010 ( .A(N1054), .B(n356), .Y(n1002) );
  NAND2XL U1011 ( .A(N1051), .B(n356), .Y(n1008) );
  AOI21XL U1012 ( .A0(SHA256_result[210]), .A1(n399), .B0(n390), .Y(n1007) );
  NAND2XL U1013 ( .A(N1049), .B(n356), .Y(n1012) );
  AOI21XL U1014 ( .A0(SHA256_result[208]), .A1(n399), .B0(n390), .Y(n1011) );
  NAND2XL U1015 ( .A(N1020), .B(n371), .Y(n919) );
  AOI21XL U1016 ( .A0(n399), .A1(SHA256_result[179]), .B0(n388), .Y(n918) );
  OAI211XL U1017 ( .A0(n1319), .A1(n26), .B0(n921), .C0(n920), .Y(n4648) );
  NAND2XL U1018 ( .A(N1019), .B(n372), .Y(n921) );
  AOI21XL U1019 ( .A0(n399), .A1(n32), .B0(n388), .Y(n920) );
  OAI21X4 U1020 ( .A0(SHA256_result[205]), .A1(SHA256_result[237]), .B0(
        SHA256_result[173]), .Y(n1070) );
  NAND2XL U1021 ( .A(SHA256_result[133]), .B(n399), .Y(n874) );
  NAND2XL U1022 ( .A(N974), .B(n354), .Y(n873) );
  NAND3BXL U1023 ( .AN(n883), .B(n376), .C(n882), .Y(n4631) );
  NAND2XL U1024 ( .A(SHA256_result[131]), .B(n399), .Y(n882) );
  NAND3BXL U1025 ( .AN(n879), .B(n375), .C(n878), .Y(n4630) );
  NAND2XL U1026 ( .A(SHA256_result[132]), .B(n399), .Y(n878) );
  NAND2XL U1027 ( .A(N973), .B(n353), .Y(n877) );
  NAND3BXL U1028 ( .AN(n890), .B(n375), .C(n889), .Y(n4633) );
  NAND2XL U1029 ( .A(SHA256_result[129]), .B(n399), .Y(n889) );
  NAND2XL U1030 ( .A(N970), .B(n369), .Y(n888) );
  NAND2XL U1031 ( .A(SHA256_result[223]), .B(n399), .Y(n978) );
  NAND2XL U1032 ( .A(SHA256_result[217]), .B(n399), .Y(n991) );
  NAND2XL U1033 ( .A(N1058), .B(n370), .Y(n990) );
  NAND3BXL U1034 ( .AN(n995), .B(n375), .C(n994), .Y(n4674) );
  NAND2XL U1035 ( .A(SHA256_result[216]), .B(n399), .Y(n994) );
  NAND2XL U1036 ( .A(N1057), .B(n356), .Y(n993) );
  NAND3BXL U1037 ( .AN(n1000), .B(n376), .C(n999), .Y(n4676) );
  NAND2XL U1038 ( .A(SHA256_result[214]), .B(n399), .Y(n999) );
  NAND2XL U1039 ( .A(N1055), .B(n356), .Y(n998) );
  NAND2XL U1040 ( .A(SHA256_result[138]), .B(n399), .Y(n857) );
  NAND2XL U1041 ( .A(N979), .B(n354), .Y(n856) );
  NAND3BXL U1042 ( .AN(n865), .B(n382), .C(n864), .Y(n4626) );
  NAND2XL U1043 ( .A(SHA256_result[136]), .B(n399), .Y(n864) );
  NAND2XL U1044 ( .A(N977), .B(n354), .Y(n863) );
  NAND2XL U1045 ( .A(N871), .B(n807), .Y(n452) );
  AOI21XL U1046 ( .A0(n344), .A1(SHA256_result[21]), .B0(n328), .Y(n476) );
  AOI21XL U1047 ( .A0(n345), .A1(SHA256_result[27]), .B0(n328), .Y(n459) );
  NAND2XL U1048 ( .A(n340), .B(SHA256_result[57]), .Y(n466) );
  AOI21XL U1049 ( .A0(n345), .A1(SHA256_result[25]), .B0(n328), .Y(n464) );
  NAND2XL U1050 ( .A(n340), .B(n119), .Y(n469) );
  AOI21XL U1051 ( .A0(n345), .A1(SHA256_result[24]), .B0(n328), .Y(n467) );
  AOI21XL U1052 ( .A0(n345), .A1(SHA256_result[23]), .B0(n328), .Y(n470) );
  AOI21XL U1053 ( .A0(n345), .A1(SHA256_result[22]), .B0(n328), .Y(n473) );
  AOI21XL U1054 ( .A0(n345), .A1(SHA256_result[15]), .B0(n328), .Y(n489) );
  INVXL U1055 ( .A(SHA256_result[161]), .Y(n969) );
  NAND3BX2 U1056 ( .AN(n442), .B(n2878), .C(n1221), .Y(n448) );
  NAND2XL U1057 ( .A(n442), .B(n2878), .Y(n440) );
  AOI31XL U1058 ( .A0(n3963), .A1(n2878), .A2(n425), .B0(n1261), .Y(n3502) );
  INVXL U1059 ( .A(n3378), .Y(n1261) );
  MX2XL U1060 ( .A(SHA256_result[149]), .B(SHA256_result[181]), .S0(n438), .Y(
        mux1[21]) );
  MX2XL U1061 ( .A(SHA256_result[145]), .B(SHA256_result[177]), .S0(n438), .Y(
        mux1[17]) );
  MX2XL U1062 ( .A(SHA256_result[147]), .B(SHA256_result[179]), .S0(n438), .Y(
        mux1[19]) );
  NOR2XL U1063 ( .A(round[6]), .B(n423), .Y(n4249) );
  MX2XL U1064 ( .A(SHA256_result[144]), .B(SHA256_result[176]), .S0(n438), .Y(
        mux1[16]) );
  MX2XL U1065 ( .A(SHA256_result[150]), .B(SHA256_result[182]), .S0(n438), .Y(
        mux1[22]) );
  MX2XL U1066 ( .A(SHA256_result[146]), .B(n32), .S0(n438), .Y(mux1[18]) );
  MX2XL U1067 ( .A(SHA256_result[148]), .B(SHA256_result[180]), .S0(n438), .Y(
        mux1[20]) );
  MX2XL U1068 ( .A(SHA256_result[152]), .B(SHA256_result[184]), .S0(n438), .Y(
        mux1[24]) );
  MX2XL U1069 ( .A(SHA256_result[153]), .B(n86), .S0(n438), .Y(mux1[25]) );
  MX2XL U1070 ( .A(SHA256_result[151]), .B(SHA256_result[183]), .S0(n438), .Y(
        mux1[23]) );
  AND2X1 U1071 ( .A(n1221), .B(n4247), .Y(n256) );
  AOI211XL U1072 ( .A0(n1264), .A1(n2906), .B0(n4237), .C0(n4238), .Y(n4236)
         );
  AOI21XL U1073 ( .A0(n4000), .A1(n258), .B0(n1250), .Y(n4234) );
  AOI21XL U1074 ( .A0(n258), .A1(n1224), .B0(n3949), .Y(n4228) );
  AOI211XL U1075 ( .A0(n4231), .A1(n427), .B0(n4232), .C0(n4017), .Y(n4230) );
  AOI32XL U1076 ( .A0(n422), .A1(n427), .A2(n249), .B0(n4103), .B1(n1223), .Y(
        n4220) );
  AOI211XL U1077 ( .A0(n4012), .A1(n253), .B0(n1252), .C0(n4223), .Y(n4222) );
  AOI31XL U1078 ( .A0(n1224), .A1(n2906), .A2(n4016), .B0(n4226), .Y(n4221) );
  AOI222XL U1079 ( .A0(n4193), .A1(n432), .B0(n4071), .B1(n4042), .C0(n4194), 
        .C1(n2906), .Y(n4186) );
  NOR3XL U1080 ( .A(n3955), .B(n4058), .C(n1262), .Y(n4187) );
  AOI211XL U1081 ( .A0(n3962), .A1(n429), .B0(n4189), .C0(n4190), .Y(n4188) );
  AOI2BB2XL U1082 ( .B0(n3947), .B1(n2925), .A0N(n290), .A1N(n3948), .Y(n3940)
         );
  AOI22XL U1083 ( .A0(n3964), .A1(n259), .B0(n3965), .B1(n286), .Y(n3951) );
  NOR3XL U1084 ( .A(n3961), .B(n3962), .C(n3963), .Y(n3952) );
  AOI221XL U1085 ( .A0(n3954), .A1(n320), .B0(n3955), .B1(n2925), .C0(n3956), 
        .Y(n3953) );
  AOI2BB1XL U1086 ( .A0N(n3955), .A1N(n3973), .B0(n2925), .Y(n4171) );
  NOR2BX1 U1087 ( .AN(round[4]), .B(n319), .Y(n257) );
  NOR2XL U1088 ( .A(n2938), .B(n431), .Y(n4016) );
  NOR2XL U1089 ( .A(n2938), .B(n424), .Y(n4027) );
  NOR2XL U1090 ( .A(n2906), .B(n808), .Y(n4029) );
  NOR3XL U1091 ( .A(n2925), .B(n427), .C(n1275), .Y(n4149) );
  OAI31XL U1092 ( .A0(n2938), .A1(n255), .A2(n1305), .B0(n3972), .Y(n3983) );
  NOR3XL U1093 ( .A(n2925), .B(n431), .C(n1267), .Y(n4074) );
  NOR2XL U1094 ( .A(n2925), .B(n2906), .Y(n4051) );
  NOR2XL U1095 ( .A(n3985), .B(n2925), .Y(n4193) );
  AOI211XL U1096 ( .A0(n320), .A1(n2925), .B0(n4012), .C0(n4192), .Y(n4191) );
  AOI21XL U1097 ( .A0(n1302), .A1(n1303), .B0(n429), .Y(n4192) );
  AOI22XL U1098 ( .A0(n318), .A1(n4053), .B0(n286), .B1(n422), .Y(n4050) );
  NAND2XL U1099 ( .A(n4042), .B(n2925), .Y(n4124) );
  MX2XL U1100 ( .A(SHA256_result[25]), .B(SHA256_result[57]), .S0(
        mux_control_0_), .Y(mux2[25]) );
  MX2XL U1101 ( .A(SHA256_result[26]), .B(SHA256_result[58]), .S0(
        mux_control_0_), .Y(mux2[26]) );
  AOI31XL U1102 ( .A0(n1271), .A1(n1253), .A2(n4087), .B0(n2906), .Y(n4223) );
  AOI222XL U1103 ( .A0(n253), .A1(n4014), .B0(n4013), .B1(n2925), .C0(n3973), 
        .C1(n318), .Y(n4209) );
  AOI221XL U1104 ( .A0(n4012), .A1(n4055), .B0(n3963), .B1(n320), .C0(n4214), 
        .Y(n4208) );
  AOI22XL U1105 ( .A0(n3973), .A1(n2925), .B0(n257), .B1(n286), .Y(n4141) );
  AOI211XL U1106 ( .A0(n3954), .A1(n4042), .B0(n4112), .C0(n3984), .Y(n4111)
         );
  AOI22XL U1107 ( .A0(n4114), .A1(n426), .B0(n4066), .B1(n2925), .Y(n4109) );
  AOI22XL U1108 ( .A0(n431), .A1(n4097), .B0(n4063), .B1(n2906), .Y(n4089) );
  NOR2XL U1109 ( .A(n2938), .B(n320), .Y(n3946) );
  NOR3XL U1110 ( .A(n430), .B(n255), .C(n2906), .Y(n4158) );
  NAND2XL U1111 ( .A(output_enable), .B(n3114), .Y(n3677) );
  NOR2XL U1112 ( .A(n2925), .B(n2947), .Y(n4225) );
  OAI33XL U1113 ( .A0(n290), .A1(n422), .A2(n1306), .B0(n1256), .B1(n2906), 
        .B2(n289), .Y(n4238) );
  MX2XL U1114 ( .A(SHA256_result[24]), .B(n119), .S0(mux_control_0_), .Y(
        mux2[24]) );
  AOI22XL U1115 ( .A0(n3708), .A1(SHA256_result[91]), .B0(n3709), .B1(
        SHA256_result[95]), .Y(n3698) );
  AOI22XL U1116 ( .A0(n3708), .A1(n31), .B0(n3709), .B1(SHA256_result[92]), 
        .Y(n3885) );
  AOI22XL U1117 ( .A0(n3708), .A1(SHA256_result[89]), .B0(n3709), .B1(
        SHA256_result[93]), .Y(n3837) );
  AOI22XL U1118 ( .A0(n3708), .A1(SHA256_result[90]), .B0(n3709), .B1(
        SHA256_result[94]), .Y(n3795) );
  MX2XL U1119 ( .A(SHA256_result[27]), .B(SHA256_result[59]), .S0(
        mux_control_0_), .Y(mux2[27]) );
  AOI22XL U1120 ( .A0(n3759), .A1(SHA256_result[218]), .B0(n3760), .B1(
        SHA256_result[222]), .Y(n3815) );
  AOI22XL U1121 ( .A0(n3757), .A1(SHA256_result[210]), .B0(n3758), .B1(
        SHA256_result[214]), .Y(n3816) );
  AOI21XL U1122 ( .A0(n1259), .A1(n4107), .B0(n2925), .Y(n4130) );
  AOI2BB1XL U1123 ( .A0N(n4000), .A1N(n4147), .B0(n2906), .Y(n4146) );
  AOI22XL U1124 ( .A0(n3720), .A1(SHA256_result[57]), .B0(n3721), .B1(
        SHA256_result[61]), .Y(n3841) );
  AOI22XL U1125 ( .A0(n3720), .A1(SHA256_result[58]), .B0(n3721), .B1(
        SHA256_result[62]), .Y(n3799) );
  AOI22XL U1126 ( .A0(n3720), .A1(SHA256_result[59]), .B0(n3721), .B1(
        SHA256_result[63]), .Y(n3710) );
  AOI22XL U1127 ( .A0(n3720), .A1(n119), .B0(n3721), .B1(SHA256_result[60]), 
        .Y(n3895) );
  AOI22XL U1128 ( .A0(n3771), .A1(SHA256_result[184]), .B0(n3772), .B1(
        SHA256_result[188]), .Y(n3927) );
  AOI22XL U1129 ( .A0(n3769), .A1(SHA256_result[176]), .B0(n3770), .B1(
        SHA256_result[180]), .Y(n3928) );
  AOI22XL U1130 ( .A0(n3771), .A1(SHA256_result[186]), .B0(n3772), .B1(
        SHA256_result[190]), .Y(n3819) );
  AOI22XL U1131 ( .A0(n3769), .A1(n32), .B0(n3770), .B1(SHA256_result[182]), 
        .Y(n3820) );
  AOI22XL U1132 ( .A0(n3771), .A1(n86), .B0(n3772), .B1(SHA256_result[189]), 
        .Y(n3861) );
  AOI22XL U1133 ( .A0(n3769), .A1(SHA256_result[177]), .B0(n3770), .B1(
        SHA256_result[181]), .Y(n3862) );
  AOI22XL U1134 ( .A0(n3771), .A1(SHA256_result[187]), .B0(n3772), .B1(
        SHA256_result[191]), .Y(n3761) );
  AOI22XL U1135 ( .A0(n3769), .A1(SHA256_result[179]), .B0(n3770), .B1(
        SHA256_result[183]), .Y(n3762) );
  AOI22XL U1136 ( .A0(n3759), .A1(SHA256_result[219]), .B0(n3760), .B1(
        SHA256_result[223]), .Y(n3749) );
  AOI22XL U1137 ( .A0(n3757), .A1(SHA256_result[211]), .B0(n3758), .B1(
        SHA256_result[215]), .Y(n3750) );
  AOI22XL U1138 ( .A0(n3759), .A1(SHA256_result[217]), .B0(n3760), .B1(
        SHA256_result[221]), .Y(n3857) );
  AOI22XL U1139 ( .A0(n3757), .A1(SHA256_result[209]), .B0(n3758), .B1(
        SHA256_result[213]), .Y(n3858) );
  AOI22XL U1140 ( .A0(n3759), .A1(SHA256_result[216]), .B0(n3760), .B1(
        SHA256_result[220]), .Y(n3921) );
  AOI22XL U1141 ( .A0(n3757), .A1(SHA256_result[208]), .B0(n3758), .B1(
        SHA256_result[212]), .Y(n3922) );
  AOI22XL U1142 ( .A0(n3679), .A1(SHA256_result[3]), .B0(n3726), .B1(
        SHA256_result[7]), .Y(n3725) );
  AOI22XL U1143 ( .A0(n3679), .A1(SHA256_result[0]), .B0(n3726), .B1(
        SHA256_result[4]), .Y(n3906) );
  AOI22XL U1144 ( .A0(n3679), .A1(SHA256_result[1]), .B0(n3726), .B1(
        SHA256_result[5]), .Y(n3848) );
  AOI22XL U1145 ( .A0(n3679), .A1(SHA256_result[2]), .B0(n3726), .B1(
        SHA256_result[6]), .Y(n3806) );
  AOI22XL U1146 ( .A0(n3747), .A1(n300), .B0(n3748), .B1(n296), .Y(n3913) );
  AOI22XL U1147 ( .A0(n3745), .A1(n308), .B0(n3746), .B1(n304), .Y(n3914) );
  AND3X1 U1148 ( .A(n3114), .B(n2878), .C(inner_busy), .Y(n266) );
  INVXL U1149 ( .A(n2947), .Y(n424) );
  NOR3XL U1150 ( .A(n1280), .B(n432), .C(n2906), .Y(n4178) );
  AOI22XL U1151 ( .A0(n3727), .A1(SHA256_result[8]), .B0(n3728), .B1(
        SHA256_result[12]), .Y(n3905) );
  AOI22XL U1152 ( .A0(n3727), .A1(SHA256_result[10]), .B0(n3728), .B1(
        SHA256_result[14]), .Y(n3805) );
  AOI22XL U1153 ( .A0(n3727), .A1(SHA256_result[11]), .B0(n3728), .B1(
        SHA256_result[15]), .Y(n3724) );
  AOI22XL U1154 ( .A0(n3727), .A1(SHA256_result[9]), .B0(n3728), .B1(
        SHA256_result[13]), .Y(n3847) );
  AOI22XL U1155 ( .A0(n3779), .A1(SHA256_result[139]), .B0(n3780), .B1(
        SHA256_result[143]), .Y(n3775) );
  AOI22XL U1156 ( .A0(n3779), .A1(SHA256_result[136]), .B0(n3780), .B1(
        SHA256_result[140]), .Y(n3937) );
  AOI22XL U1157 ( .A0(n3779), .A1(SHA256_result[137]), .B0(n3780), .B1(
        SHA256_result[141]), .Y(n3867) );
  AOI22XL U1158 ( .A0(n3779), .A1(SHA256_result[138]), .B0(n3780), .B1(
        SHA256_result[142]), .Y(n3825) );
  AOI22XL U1159 ( .A0(n3777), .A1(SHA256_result[128]), .B0(n3778), .B1(
        SHA256_result[132]), .Y(n3938) );
  AOI22XL U1160 ( .A0(n3777), .A1(SHA256_result[129]), .B0(n3778), .B1(
        SHA256_result[133]), .Y(n3868) );
  AOI22XL U1161 ( .A0(n3777), .A1(SHA256_result[131]), .B0(n3778), .B1(
        SHA256_result[135]), .Y(n3776) );
  AOI31XL U1162 ( .A0(n432), .A1(n2906), .A2(n4027), .B0(n4028), .Y(n4023) );
  AOI22XL U1163 ( .A0(n3777), .A1(SHA256_result[130]), .B0(n3778), .B1(
        SHA256_result[134]), .Y(n3826) );
  INVXL U1164 ( .A(n103), .Y(n715) );
  INVXL U1165 ( .A(SHA256_result[211]), .Y(n1320) );
  INVXL U1166 ( .A(n110), .Y(n703) );
  INVXL U1167 ( .A(SHA256_result[179]), .Y(n1335) );
  INVXL U1168 ( .A(SHA256_result[186]), .Y(n1341) );
  INVXL U1169 ( .A(n32), .Y(n1334) );
  INVXL U1170 ( .A(SHA256_result[182]), .Y(n1338) );
  INVXL U1171 ( .A(SHA256_result[219]), .Y(n1235) );
  INVXL U1172 ( .A(SHA256_result[210]), .Y(n1319) );
  INVXL U1173 ( .A(SHA256_result[213]), .Y(n1322) );
  INVXL U1174 ( .A(SHA256_result[184]), .Y(n1340) );
  INVXL U1175 ( .A(SHA256_result[176]), .Y(n1332) );
  INVXL U1176 ( .A(SHA256_result[214]), .Y(n1323) );
  INVXL U1177 ( .A(SHA256_result[218]), .Y(n1234) );
  INVXL U1178 ( .A(SHA256_result[187]), .Y(n1342) );
  INVXL U1179 ( .A(SHA256_result[58]), .Y(n1398) );
  INVXL U1180 ( .A(SHA256_result[181]), .Y(n1337) );
  INVXL U1181 ( .A(SHA256_result[183]), .Y(n1339) );
  INVXL U1182 ( .A(SHA256_result[180]), .Y(n1336) );
  INVXL U1183 ( .A(SHA256_result[215]), .Y(n1324) );
  INVXL U1184 ( .A(SHA256_result[212]), .Y(n1321) );
  INVXL U1185 ( .A(SHA256_result[209]), .Y(n1318) );
  INVXL U1186 ( .A(SHA256_result[177]), .Y(n1333) );
  NAND3XL U1187 ( .A(n434), .B(n2938), .C(n253), .Y(n3985) );
  NAND2XL U1188 ( .A(n257), .B(n434), .Y(n4086) );
  INVX1 U1189 ( .A(n359), .Y(n355) );
  INVX1 U1190 ( .A(n386), .Y(n381) );
  INVX1 U1191 ( .A(n385), .Y(n383) );
  INVX1 U1192 ( .A(n385), .Y(n384) );
  INVX1 U1193 ( .A(n388), .Y(n375) );
  INVX1 U1194 ( .A(n387), .Y(n376) );
  INVX1 U1195 ( .A(n387), .Y(n377) );
  INVX1 U1196 ( .A(n442), .Y(n1219) );
  OAI21XL U1197 ( .A0(n808), .A1(n1298), .B0(n1277), .Y(n4207) );
  INVX1 U1198 ( .A(n358), .Y(n356) );
  INVX1 U1199 ( .A(n347), .Y(n341) );
  INVX1 U1200 ( .A(n800), .Y(n347) );
  INVX1 U1201 ( .A(n1198), .Y(n385) );
  INVX1 U1202 ( .A(n373), .Y(n360) );
  INVX1 U1203 ( .A(n800), .Y(n346) );
  INVX1 U1204 ( .A(n751), .Y(n325) );
  INVX1 U1205 ( .A(n1198), .Y(n388) );
  INVX1 U1206 ( .A(n1198), .Y(n387) );
  INVX1 U1207 ( .A(n370), .Y(n366) );
  INVX1 U1208 ( .A(n369), .Y(n365) );
  INVX1 U1209 ( .A(n124), .Y(n364) );
  INVX1 U1210 ( .A(n371), .Y(n363) );
  INVX1 U1211 ( .A(n372), .Y(n362) );
  INVX1 U1212 ( .A(n372), .Y(n361) );
  INVX1 U1213 ( .A(n369), .Y(n368) );
  INVX1 U1214 ( .A(n370), .Y(n367) );
  INVX1 U1215 ( .A(n247), .Y(n348) );
  INVX1 U1216 ( .A(n247), .Y(n349) );
  INVX1 U1217 ( .A(n247), .Y(n350) );
  INVX1 U1218 ( .A(n247), .Y(n351) );
  INVX1 U1219 ( .A(n4012), .Y(n1301) );
  NOR2X1 U1220 ( .A(n808), .B(n1305), .Y(n4017) );
  INVX1 U1221 ( .A(n4015), .Y(n1276) );
  INVX1 U1222 ( .A(n4044), .Y(n1291) );
  INVX1 U1223 ( .A(n4063), .Y(n1253) );
  INVX1 U1224 ( .A(n4041), .Y(n1270) );
  INVX1 U1225 ( .A(n4137), .Y(n1260) );
  NAND2BX1 U1226 ( .AN(n4081), .B(n1291), .Y(n4165) );
  OAI21XL U1227 ( .A0(n1305), .A1(n1251), .B0(n1255), .Y(n4114) );
  INVX1 U1228 ( .A(n4036), .Y(n1255) );
  INVX1 U1229 ( .A(n4057), .Y(n1278) );
  INVX1 U1230 ( .A(n4164), .Y(n1277) );
  INVX1 U1231 ( .A(n4030), .Y(n1299) );
  INVX1 U1232 ( .A(n4104), .Y(n1266) );
  INVX1 U1233 ( .A(n4096), .Y(n1290) );
  INVX1 U1234 ( .A(n4040), .Y(n1264) );
  NAND2X1 U1235 ( .A(n812), .B(n450), .Y(n751) );
  NAND2XL U1236 ( .A(next_E[7]), .B(n338), .Y(n772) );
  NAND2X1 U1237 ( .A(N944), .B(n807), .Y(n773) );
  INVX1 U1238 ( .A(n1186), .Y(n374) );
  OAI221XL U1239 ( .A0(n362), .A1(n1004), .B0(n1232), .B1(n24), .C0(n1003), 
        .Y(n4678) );
  INVX1 U1240 ( .A(N1053), .Y(n1004) );
  OAI221XL U1241 ( .A0(n362), .A1(n1020), .B0(n27), .B1(n1146), .C0(n1019), 
        .Y(n4686) );
  INVX1 U1242 ( .A(N1045), .Y(n1020) );
  NAND2X1 U1243 ( .A(n247), .B(SHA256_result[204]), .Y(n1019) );
  OAI221XL U1244 ( .A0(n363), .A1(n997), .B0(n22), .B1(n1115), .C0(n996), .Y(
        n4675) );
  INVX1 U1245 ( .A(N1056), .Y(n997) );
  OAI221XL U1246 ( .A0(n361), .A1(n1036), .B0(n22), .B1(n1170), .C0(n1035), 
        .Y(n4692) );
  INVX1 U1247 ( .A(N1039), .Y(n1036) );
  NAND2X1 U1248 ( .A(n247), .B(SHA256_result[198]), .Y(n1035) );
  OAI221XL U1249 ( .A0(n361), .A1(n1038), .B0(n27), .B1(n1175), .C0(n1037), 
        .Y(n4693) );
  INVX1 U1250 ( .A(N1038), .Y(n1038) );
  NAND2X1 U1251 ( .A(n247), .B(SHA256_result[197]), .Y(n1037) );
  OAI221XL U1252 ( .A0(n362), .A1(n1047), .B0(n23), .B1(n1193), .C0(n1046), 
        .Y(n4697) );
  INVX1 U1253 ( .A(N1034), .Y(n1047) );
  NAND2X1 U1254 ( .A(n247), .B(SHA256_result[193]), .Y(n1046) );
  OAI221XL U1255 ( .A0(n362), .A1(n1006), .B0(n1231), .B1(n25), .C0(n1005), 
        .Y(n4679) );
  INVX1 U1256 ( .A(N1052), .Y(n1006) );
  NAND2X1 U1257 ( .A(n247), .B(SHA256_result[211]), .Y(n1005) );
  OAI221XL U1258 ( .A0(n362), .A1(n1016), .B0(n1226), .B1(n28), .C0(n1015), 
        .Y(n4684) );
  INVX1 U1259 ( .A(N1047), .Y(n1016) );
  NAND2X1 U1260 ( .A(n247), .B(SHA256_result[206]), .Y(n1015) );
  INVX1 U1261 ( .A(n809), .Y(n1222) );
  INVX1 U1262 ( .A(n405), .Y(n401) );
  INVX1 U1263 ( .A(n405), .Y(n403) );
  INVX1 U1264 ( .A(n1186), .Y(n371) );
  INVX1 U1265 ( .A(n1186), .Y(n372) );
  INVX1 U1266 ( .A(n1186), .Y(n369) );
  INVX1 U1267 ( .A(n1186), .Y(n370) );
  NOR2X1 U1268 ( .A(n1279), .B(n431), .Y(n4057) );
  INVX1 U1269 ( .A(n4004), .Y(n1279) );
  OAI21XL U1270 ( .A0(n1306), .A1(n289), .B0(n1296), .Y(n4032) );
  NOR2X1 U1271 ( .A(n1301), .B(n426), .Y(n4227) );
  AOI31X1 U1272 ( .A0(n3993), .A1(n3994), .A2(n3995), .B0(n418), .Y(N3160) );
  NOR3X1 U1273 ( .A(n3996), .B(n3997), .C(n3998), .Y(n3995) );
  AOI22X1 U1274 ( .A0(n1269), .A1(n431), .B0(n4004), .B1(n429), .Y(n3993) );
  AOI211X1 U1275 ( .A0(n4000), .A1(n3954), .B0(n4001), .C0(n4002), .Y(n3994)
         );
  BUFX3 U1276 ( .A(n1220), .Y(n286) );
  INVX1 U1277 ( .A(n255), .Y(n1220) );
  INVX1 U1278 ( .A(n808), .Y(n1224) );
  NOR2X1 U1279 ( .A(n1292), .B(n1305), .Y(n4044) );
  OAI222XL U1280 ( .A0(n425), .A1(n1301), .B0(n427), .B1(n1271), .C0(n255), 
        .C1(n1276), .Y(n4136) );
  NOR2X1 U1281 ( .A(n1295), .B(n425), .Y(n4024) );
  NOR2X1 U1282 ( .A(n1304), .B(n423), .Y(n4015) );
  NOR2X1 U1283 ( .A(n1254), .B(n290), .Y(n4063) );
  INVX1 U1284 ( .A(n4000), .Y(n1271) );
  NOR2X1 U1285 ( .A(n1291), .B(n430), .Y(n4137) );
  NOR2X1 U1286 ( .A(n1258), .B(n434), .Y(n4043) );
  NOR2X1 U1287 ( .A(n1295), .B(n429), .Y(n4081) );
  NOR2X1 U1288 ( .A(n1271), .B(n431), .Y(n4041) );
  INVX1 U1289 ( .A(n253), .Y(n1251) );
  OAI21XL U1290 ( .A0(n2947), .A1(n1306), .B0(n1276), .Y(n3989) );
  INVX1 U1291 ( .A(n4093), .Y(n1269) );
  NOR2X1 U1292 ( .A(n1303), .B(n2947), .Y(n4088) );
  NOR2X1 U1293 ( .A(n3955), .B(n4009), .Y(n4108) );
  OAI21XL U1294 ( .A0(n426), .A1(n1271), .B0(n4087), .Y(n4084) );
  NAND3X1 U1295 ( .A(n1270), .B(n1281), .C(n4010), .Y(n4008) );
  INVX1 U1296 ( .A(n4240), .Y(n1250) );
  INVX1 U1297 ( .A(n4233), .Y(n1258) );
  NAND3X1 U1298 ( .A(n1270), .B(n1246), .C(n4040), .Y(n4037) );
  AOI2BB1X1 U1299 ( .A0N(n3955), .A1N(n4039), .B0(n431), .Y(n4038) );
  BUFX3 U1300 ( .A(n1288), .Y(n289) );
  INVX1 U1301 ( .A(n4055), .Y(n1288) );
  NOR2X1 U1302 ( .A(n1306), .B(n431), .Y(n3954) );
  NOR2X1 U1303 ( .A(n289), .B(n429), .Y(n3973) );
  INVX1 U1304 ( .A(n3960), .Y(n1256) );
  OAI211X1 U1305 ( .A0(n434), .A1(n4067), .B0(n1276), .C0(n1305), .Y(n4097) );
  NOR2X1 U1306 ( .A(n4151), .B(n431), .Y(n3962) );
  NOR2X1 U1307 ( .A(n1292), .B(n808), .Y(n4066) );
  NOR2X1 U1308 ( .A(n4086), .B(n422), .Y(n4056) );
  NOR2X1 U1309 ( .A(n1275), .B(n255), .Y(n3947) );
  NOR2X1 U1310 ( .A(n289), .B(n1275), .Y(n4147) );
  OAI21XL U1311 ( .A0(n1298), .A1(n1256), .B0(n1273), .Y(n4190) );
  NOR2X1 U1312 ( .A(n1306), .B(n426), .Y(n4071) );
  OAI2BB2X1 U1313 ( .B0(n255), .B1(n1304), .A0N(n249), .A1N(n4059), .Y(n3984)
         );
  NOR2X1 U1314 ( .A(n289), .B(n422), .Y(n4013) );
  NOR2X1 U1315 ( .A(n1306), .B(n255), .Y(n4096) );
  AOI31X1 U1316 ( .A0(n1286), .A1(n1273), .A2(n1272), .B0(n434), .Y(n4065) );
  INVX1 U1317 ( .A(n4003), .Y(n1286) );
  INVX1 U1318 ( .A(n4066), .Y(n1272) );
  INVX1 U1319 ( .A(n4150), .Y(n1274) );
  NAND2X1 U1320 ( .A(n4055), .B(n4042), .Y(n4040) );
  NOR2X1 U1321 ( .A(n1299), .B(n422), .Y(n3991) );
  NOR2X1 U1322 ( .A(n3960), .B(n4083), .Y(n4067) );
  NOR2X1 U1323 ( .A(n3992), .B(n426), .Y(n4164) );
  INVX1 U1324 ( .A(n4083), .Y(n1280) );
  NOR2X1 U1325 ( .A(n1256), .B(n434), .Y(n4036) );
  NAND2X1 U1326 ( .A(n429), .B(n425), .Y(n4026) );
  NOR2X1 U1327 ( .A(n289), .B(n1304), .Y(n4075) );
  NAND3BX1 U1328 ( .AN(n4058), .B(n4019), .C(n1295), .Y(n4198) );
  AOI21X1 U1329 ( .A0(n3999), .A1(n1290), .B0(n429), .Y(n4245) );
  OAI21XL U1330 ( .A0(n431), .A1(n1256), .B0(n1287), .Y(n4095) );
  NAND3X1 U1331 ( .A(n1295), .B(n4094), .C(n1246), .Y(n4092) );
  OAI21XL U1332 ( .A0(n1303), .A1(n290), .B0(n1279), .Y(n3986) );
  AOI21X1 U1333 ( .A0(n3992), .A1(n1267), .B0(n290), .Y(n4172) );
  NAND3X1 U1334 ( .A(n1253), .B(n1259), .C(n3999), .Y(n3996) );
  INVX1 U1335 ( .A(n4151), .Y(n1289) );
  INVX1 U1336 ( .A(n4105), .Y(n1283) );
  AOI21X1 U1337 ( .A0(n1255), .A1(n1257), .B0(n431), .Y(n3976) );
  INVX1 U1338 ( .A(n4122), .Y(n1282) );
  OAI21XL U1339 ( .A0(n1294), .A1(n3950), .B0(n429), .Y(n4183) );
  INVX1 U1340 ( .A(n3999), .Y(n1294) );
  NAND2X1 U1341 ( .A(n4017), .B(n431), .Y(n4184) );
  AOI21X1 U1342 ( .A0(n4086), .A1(n1254), .B0(n255), .Y(n4085) );
  AOI2BB1X1 U1343 ( .A0N(n4025), .A1N(n4132), .B0(n429), .Y(n4131) );
  AOI2BB1X1 U1344 ( .A0N(n3947), .A1N(n4003), .B0(n434), .Y(n4002) );
  INVX1 U1345 ( .A(next_A[0]), .Y(n1199) );
  NOR2X1 U1346 ( .A(n426), .B(n429), .Y(n4059) );
  INVXL U1347 ( .A(next_E[18]), .Y(n734) );
  NOR2X1 U1348 ( .A(n180), .B(n104), .Y(n805) );
  NAND2BXL U1349 ( .AN(n795), .B(next_E[15]), .Y(n744) );
  NAND2BX1 U1350 ( .AN(n26), .B(next_A[31]), .Y(n1084) );
  OAI221XL U1351 ( .A0(n360), .A1(n1149), .B0(n28), .B1(n1148), .C0(n1147), 
        .Y(n4752) );
  INVXL U1352 ( .A(next_A[12]), .Y(n1148) );
  NAND2X1 U1353 ( .A(SHA256_result[236]), .B(n247), .Y(n1147) );
  INVX1 U1354 ( .A(N1077), .Y(n1149) );
  NAND2X1 U1355 ( .A(n440), .B(n423), .Y(n441) );
  XOR3X2 U1356 ( .A(n312), .B(n304), .C(n295), .Y(f3_A_32[7]) );
  NAND2BX1 U1357 ( .AN(first_block_core), .B(n107), .Y(n3115) );
  INVX1 U1358 ( .A(n448), .Y(n815) );
  OAI211X1 U1359 ( .A0(n330), .A1(n787), .B0(n786), .C0(n785), .Y(n4567) );
  NAND2X1 U1360 ( .A(N940), .B(n807), .Y(n786) );
  OAI211X1 U1361 ( .A0(n335), .A1(n791), .B0(n790), .C0(n789), .Y(n4568) );
  INVX1 U1362 ( .A(next_E[2]), .Y(n791) );
  OAI211X1 U1363 ( .A0(n1157), .A1(n21), .B0(n1156), .C0(n1155), .Y(n4754) );
  INVXL U1364 ( .A(next_A[10]), .Y(n1157) );
  NAND2X1 U1365 ( .A(N1075), .B(n357), .Y(n1156) );
  AOI21X1 U1366 ( .A0(n311), .A1(n399), .B0(n390), .Y(n1155) );
  OAI211X1 U1367 ( .A0(n334), .A1(n794), .B0(n793), .C0(n792), .Y(n4569) );
  NAND2X1 U1368 ( .A(N938), .B(n807), .Y(n793) );
  XOR3X2 U1369 ( .A(n316), .B(SHA256_result[236]), .C(n303), .Y(f3_A_32[31])
         );
  XOR3X2 U1370 ( .A(n315), .B(SHA256_result[237]), .C(n302), .Y(f3_A_32[0]) );
  NAND2XL U1371 ( .A(next_E[9]), .B(n339), .Y(n766) );
  NAND2X1 U1372 ( .A(N946), .B(n807), .Y(n765) );
  NAND4X1 U1373 ( .A(n1109), .B(n1108), .C(n382), .D(n1107), .Y(n4739) );
  NAND2XL U1374 ( .A(next_A[25]), .B(n29), .Y(n1109) );
  NAND2X1 U1375 ( .A(N1090), .B(n357), .Y(n1108) );
  NAND2XL U1376 ( .A(next_A[19]), .B(n29), .Y(n1128) );
  NAND2XL U1377 ( .A(next_A[15]), .B(n30), .Y(n1138) );
  NAND2XL U1378 ( .A(next_A[16]), .B(n29), .Y(n1135) );
  NAND4X1 U1379 ( .A(n1141), .B(n1140), .C(n384), .D(n1139), .Y(n4750) );
  NAND2XL U1380 ( .A(next_A[14]), .B(n29), .Y(n1141) );
  NAND2X1 U1381 ( .A(N1079), .B(n357), .Y(n1140) );
  NAND4X1 U1382 ( .A(n1144), .B(n1143), .C(n383), .D(n1142), .Y(n4751) );
  NAND2X1 U1383 ( .A(N1078), .B(n357), .Y(n1143) );
  NAND3X1 U1384 ( .A(n776), .B(n775), .C(n774), .Y(n4564) );
  NAND2XL U1385 ( .A(next_E[6]), .B(n339), .Y(n776) );
  NAND2X1 U1386 ( .A(N943), .B(n807), .Y(n775) );
  XOR3X2 U1387 ( .A(n16), .B(n302), .C(n293), .Y(f3_A_32[9]) );
  XOR3X2 U1388 ( .A(n313), .B(n307), .C(n298), .Y(f3_A_32[4]) );
  XOR3X2 U1389 ( .A(n317), .B(SHA256_result[236]), .C(n301), .Y(f3_A_32[10])
         );
  XOR3X2 U1390 ( .A(n311), .B(n303), .C(n294), .Y(f3_A_32[8]) );
  XOR3X2 U1391 ( .A(n314), .B(n308), .C(n299), .Y(f3_A_32[3]) );
  BUFX3 U1392 ( .A(n798), .Y(n287) );
  NAND3BX1 U1393 ( .AN(n1204), .B(n1203), .C(n1202), .Y(n4764) );
  OAI211X1 U1394 ( .A0(n332), .A1(n779), .B0(n778), .C0(n777), .Y(n4565) );
  INVXL U1395 ( .A(next_E[5]), .Y(n779) );
  NAND2X1 U1396 ( .A(N942), .B(n807), .Y(n778) );
  OAI211X1 U1397 ( .A0(n335), .A1(n783), .B0(n782), .C0(n781), .Y(n4566) );
  INVX1 U1398 ( .A(next_E[4]), .Y(n783) );
  NAND2XL U1399 ( .A(next_E[8]), .B(n338), .Y(n769) );
  NAND2X1 U1400 ( .A(N945), .B(n807), .Y(n770) );
  NAND3BX1 U1401 ( .AN(n1162), .B(n379), .C(n1161), .Y(n4755) );
  INVXL U1402 ( .A(next_A[9]), .Y(n1160) );
  NAND3BX1 U1403 ( .AN(n1174), .B(n379), .C(n1173), .Y(n4758) );
  INVXL U1404 ( .A(next_A[5]), .Y(n1177) );
  NAND3BX1 U1405 ( .AN(n1192), .B(n378), .C(n1191), .Y(n4762) );
  INVX1 U1406 ( .A(next_A[2]), .Y(n1190) );
  NAND3BX1 U1407 ( .AN(n1197), .B(n382), .C(n1196), .Y(n4763) );
  NAND2XL U1408 ( .A(next_E[11]), .B(n337), .Y(n758) );
  NAND2XL U1411 ( .A(n186), .B(n337), .Y(n761) );
  NAND2X1 U1414 ( .A(N947), .B(n807), .Y(n762) );
  NAND2XL U1417 ( .A(next_E[13]), .B(n339), .Y(n752) );
  NAND2X1 U1420 ( .A(N950), .B(n807), .Y(n753) );
  NAND2X1 U1421 ( .A(N1070), .B(n353), .Y(n1176) );
  NAND2X1 U1424 ( .A(N1074), .B(n357), .Y(n1159) );
  NAND2X1 U1427 ( .A(N1071), .B(n357), .Y(n1171) );
  NAND2X1 U1432 ( .A(N1067), .B(n357), .Y(n1189) );
  NAND2X1 U1437 ( .A(N1066), .B(n357), .Y(n1194) );
  NAND2X1 U1438 ( .A(n1113), .B(n1112), .Y(n4740) );
  NAND2BXL U1441 ( .AN(n22), .B(next_A[26]), .Y(n1104) );
  NAND2X1 U1444 ( .A(n1121), .B(n1120), .Y(n4742) );
  NAND2BXL U1447 ( .AN(n25), .B(next_A[22]), .Y(n1120) );
  NAND2BXL U1450 ( .AN(n21), .B(next_A[11]), .Y(n1152) );
  NAND2X1 U1451 ( .A(n1130), .B(n1129), .Y(n4746) );
  NAND2BXL U1454 ( .AN(n25), .B(next_A[18]), .Y(n1129) );
  AOI22X1 U1457 ( .A0(N1083), .A1(n353), .B0(n247), .B1(n306), .Y(n1130) );
  NAND2BXL U1462 ( .AN(n26), .B(next_A[23]), .Y(n1116) );
  NAND2X1 U1468 ( .A(n1123), .B(n1122), .Y(n4743) );
  NAND2BXL U1469 ( .AN(n26), .B(next_A[21]), .Y(n1122) );
  AOI22X1 U1470 ( .A0(N1086), .A1(n353), .B0(n247), .B1(n303), .Y(n1123) );
  NAND2X1 U1471 ( .A(n1125), .B(n1124), .Y(n4744) );
  NAND2X1 U1474 ( .A(n1132), .B(n1131), .Y(n4747) );
  AOI22X1 U1477 ( .A0(N1082), .A1(n353), .B0(n247), .B1(n307), .Y(n1132) );
  OAI222XL U1480 ( .A0(n21), .A1(n944), .B0(n368), .B1(n861), .C0(n351), .C1(
        n860), .Y(n4625) );
  INVX1 U1483 ( .A(N978), .Y(n861) );
  OAI222XL U1484 ( .A0(n25), .A1(n951), .B0(n368), .B1(n868), .C0(n350), .C1(
        n867), .Y(n4627) );
  INVX1 U1487 ( .A(N976), .Y(n868) );
  OAI222XL U1490 ( .A0(n22), .A1(n954), .B0(n366), .B1(n871), .C0(n349), .C1(
        n870), .Y(n4628) );
  INVX1 U1496 ( .A(N975), .Y(n871) );
  OAI222XL U1502 ( .A0(n25), .A1(n967), .B0(n367), .B1(n886), .C0(n349), .C1(
        n885), .Y(n4632) );
  INVX1 U1503 ( .A(N971), .Y(n886) );
  OAI222XL U1506 ( .A0(n26), .A1(n973), .B0(n368), .B1(n893), .C0(n348), .C1(
        n892), .Y(n4634) );
  INVX1 U1509 ( .A(N969), .Y(n893) );
  OAI222XL U1510 ( .A0(n24), .A1(n1166), .B0(n368), .B1(n1165), .C0(n348), 
        .C1(n1164), .Y(n4756) );
  INVXL U1513 ( .A(next_A[8]), .Y(n1166) );
  INVX1 U1516 ( .A(N1073), .Y(n1165) );
  OAI222XL U1517 ( .A0(n27), .A1(n1169), .B0(n365), .B1(n1168), .C0(n350), 
        .C1(n217), .Y(n4757) );
  INVXL U1518 ( .A(next_A[7]), .Y(n1169) );
  INVX1 U1521 ( .A(N1072), .Y(n1168) );
  OAI222XL U1524 ( .A0(n24), .A1(n1183), .B0(n368), .B1(n1182), .C0(n352), 
        .C1(n1181), .Y(n4760) );
  INVX1 U1525 ( .A(next_A[4]), .Y(n1183) );
  INVX1 U1530 ( .A(N1069), .Y(n1182) );
  OAI222XL U1531 ( .A0(n27), .A1(n1187), .B0(n367), .B1(n1185), .C0(n204), 
        .C1(n220), .Y(n4761) );
  INVX1 U1536 ( .A(N1068), .Y(n1185) );
  OAI221XL U1538 ( .A0(n361), .A1(n1042), .B0(n23), .B1(n220), .C0(n1041), .Y(
        n4695) );
  INVX1 U1539 ( .A(N1036), .Y(n1042) );
  NAND2X1 U1540 ( .A(n247), .B(n100), .Y(n1041) );
  OAI221XL U1541 ( .A0(n361), .A1(n1031), .B0(n28), .B1(n1164), .C0(n1030), 
        .Y(n4690) );
  INVX1 U1542 ( .A(N1041), .Y(n1031) );
  NAND2X1 U1543 ( .A(n247), .B(SHA256_result[200]), .Y(n1030) );
  OAI221XL U1544 ( .A0(n361), .A1(n1040), .B0(n21), .B1(n1181), .C0(n1039), 
        .Y(n4694) );
  INVX1 U1545 ( .A(N1037), .Y(n1040) );
  NAND2X1 U1546 ( .A(n247), .B(SHA256_result[196]), .Y(n1039) );
  XOR3X2 U1547 ( .A(n316), .B(SHA256_result[237]), .C(n300), .Y(f3_A_32[11])
         );
  CLKINVX3 U1548 ( .A(n430), .Y(n429) );
  XOR3X2 U1549 ( .A(n317), .B(n312), .C(n303), .Y(f3_A_32[19]) );
  XOR3X2 U1550 ( .A(n313), .B(n306), .C(n295), .Y(f3_A_32[16]) );
  XOR3X2 U1551 ( .A(n314), .B(n307), .C(n296), .Y(f3_A_32[15]) );
  XOR3X2 U1552 ( .A(n315), .B(n310), .C(n299), .Y(f3_A_32[12]) );
  INVX1 U1553 ( .A(n256), .Y(n405) );
  INVX1 U1554 ( .A(n3574), .Y(n1245) );
  NOR2X1 U1555 ( .A(n3677), .B(n3679), .Y(n3678) );
  INVX1 U1556 ( .A(n257), .Y(n1302) );
  AOI31X1 U1557 ( .A0(n4152), .A1(n4153), .A2(n4154), .B0(n417), .Y(N3146) );
  NOR3X1 U1558 ( .A(n4056), .B(n1266), .C(n3955), .Y(n4152) );
  MXI2XL U1559 ( .A(n1209), .B(n1208), .S0(mux_control_0_), .Y(mux2[5]) );
  MXI2XL U1560 ( .A(n1211), .B(n1210), .S0(mux_control_0_), .Y(mux2[4]) );
  MXI2XL U1561 ( .A(n1207), .B(n1206), .S0(mux_control_0_), .Y(mux2[6]) );
  MXI2XL U1562 ( .A(n1216), .B(n162), .S0(mux_control_0_), .Y(mux2[1]) );
  MXI2XL U1563 ( .A(n1213), .B(n1212), .S0(mux_control_0_), .Y(mux2[3]) );
  NAND2BX1 U1564 ( .AN(n3503), .B(n3502), .Y(n3501) );
  AOI31X1 U1565 ( .A0(n4167), .A1(n4168), .A2(n4169), .B0(n417), .Y(N3144) );
  NOR3X1 U1566 ( .A(n4171), .B(n1249), .C(n4172), .Y(n4167) );
  AOI31X1 U1567 ( .A0(n4133), .A1(n4134), .A2(n4135), .B0(n417), .Y(N3148) );
  AOI211X1 U1568 ( .A0(n4013), .A1(n257), .B0(n4081), .C0(n4138), .Y(n4134) );
  AOI31X1 U1569 ( .A0(n4160), .A1(n4161), .A2(n4162), .B0(n417), .Y(N3145) );
  AOI211X1 U1570 ( .A0(n4165), .A1(n425), .B0(n4166), .C0(n3969), .Y(n4160) );
  AOI31X1 U1571 ( .A0(n4060), .A1(n4061), .A2(n4062), .B0(n418), .Y(N3155) );
  NOR3X1 U1572 ( .A(n4072), .B(n4011), .C(n4058), .Y(n4061) );
  AOI31X1 U1573 ( .A0(n4115), .A1(n4116), .A2(n4117), .B0(n418), .Y(N3150) );
  NOR2BX1 U1574 ( .AN(n4052), .B(n4043), .Y(n4116) );
  AOI31X1 U1575 ( .A0(n4033), .A1(n4034), .A2(n4035), .B0(n418), .Y(N3157) );
  AOI31X1 U1576 ( .A0(n4125), .A1(n4126), .A2(n4127), .B0(n418), .Y(N3149) );
  NOR3X1 U1577 ( .A(n4130), .B(n3990), .C(n4131), .Y(n4125) );
  NOR3X1 U1578 ( .A(n1266), .B(n3963), .C(n4024), .Y(n4126) );
  AOI211X1 U1579 ( .A0(n95), .A1(n425), .B0(n4128), .C0(n4129), .Y(n4127) );
  AOI31X1 U1580 ( .A0(n4195), .A1(n4196), .A2(n4197), .B0(n417), .Y(N3140) );
  AOI221X1 U1581 ( .A0(n4015), .A1(n4055), .B0(n3965), .B1(n289), .C0(n4200), 
        .Y(n4196) );
  NOR4BX1 U1582 ( .AN(n1255), .B(n4198), .C(n4199), .D(n4017), .Y(n4197) );
  AOI31X1 U1583 ( .A0(n3979), .A1(n3980), .A2(n3981), .B0(n418), .Y(N3161) );
  AOI2BB2X1 U1584 ( .B0(n3991), .B1(n434), .A0N(n3992), .A1N(n290), .Y(n3979)
         );
  NOR3X1 U1585 ( .A(n3982), .B(n3983), .C(n3984), .Y(n3981) );
  AOI31X1 U1586 ( .A0(n4201), .A1(n4202), .A2(n4203), .B0(n417), .Y(N3139) );
  AOI21X1 U1587 ( .A0(n4158), .A1(n319), .B0(n4207), .Y(n4201) );
  NOR3X1 U1588 ( .A(n4204), .B(n3955), .C(n4041), .Y(n4203) );
  AOI31X1 U1589 ( .A0(n4174), .A1(n4175), .A2(n4176), .B0(n417), .Y(N3143) );
  NOR4BX1 U1590 ( .AN(n3985), .B(n4177), .C(n4178), .D(n1219), .Y(n4176) );
  AOI31X1 U1591 ( .A0(n4241), .A1(n4242), .A2(n4243), .B0(n417), .Y(N3133) );
  AOI222X1 U1592 ( .A0(n4225), .A1(n3946), .B0(n4071), .B1(n4027), .C0(n3960), 
        .C1(n3944), .Y(n4242) );
  AOI31X1 U1593 ( .A0(n4020), .A1(n4021), .A2(n4022), .B0(n418), .Y(N3158) );
  NOR4BX1 U1594 ( .AN(n4023), .B(n4024), .C(n4025), .D(n3998), .Y(n4022) );
  AOI221X1 U1595 ( .A0(n4029), .A1(n257), .B0(n4030), .B1(n1224), .C0(n4031), 
        .Y(n4021) );
  AOI31X1 U1596 ( .A0(n4045), .A1(n4046), .A2(n4047), .B0(n418), .Y(N3156) );
  NOR2BX1 U1597 ( .AN(n4048), .B(n4049), .Y(n4047) );
  AOI31X1 U1598 ( .A0(n1248), .A1(n4098), .A2(n4099), .B0(n418), .Y(N3152) );
  AOI222X1 U1599 ( .A0(n4003), .A1(n434), .B0(n4105), .B1(n4014), .C0(n4029), 
        .C1(n318), .Y(n4098) );
  INVX1 U1600 ( .A(n4106), .Y(n1248) );
  NOR2X1 U1601 ( .A(n4100), .B(n4101), .Y(n4099) );
  AOI31X1 U1602 ( .A0(n4005), .A1(n4006), .A2(n4007), .B0(n418), .Y(N3159) );
  AOI21X1 U1603 ( .A0(n4015), .A1(n4016), .B0(n3978), .Y(n4005) );
  NOR3X1 U1604 ( .A(n4008), .B(n4009), .C(n3991), .Y(n4007) );
  AOI31X1 U1605 ( .A0(n3966), .A1(n3967), .A2(n1263), .B0(n418), .Y(N3162) );
  INVX1 U1606 ( .A(n3968), .Y(n1263) );
  AOI31X1 U1607 ( .A0(n4180), .A1(n4181), .A2(n4182), .B0(n417), .Y(N3142) );
  AOI22X1 U1608 ( .A0(n4029), .A1(n257), .B0(n1265), .B1(n2946), .Y(n4181) );
  AOI2BB1X1 U1609 ( .A0N(n1306), .A1N(n4185), .B0(n4129), .Y(n4180) );
  XOR3X2 U1610 ( .A(n313), .B(n309), .C(n297), .Y(f3_A_32[25]) );
  XOR3X2 U1611 ( .A(n314), .B(n310), .C(n298), .Y(f3_A_32[24]) );
  XOR3X2 U1612 ( .A(n315), .B(n15), .C(n301), .Y(f3_A_32[21]) );
  XOR3X2 U1613 ( .A(n316), .B(n311), .C(n302), .Y(f3_A_32[20]) );
  AOI21X1 U1614 ( .A0(n4215), .A1(n4216), .B0(n417), .Y(N3137) );
  NOR3X1 U1615 ( .A(n4219), .B(n4190), .C(n4207), .Y(n4215) );
  AOI211X1 U1616 ( .A0(n4070), .A1(n258), .B0(n4217), .C0(n4218), .Y(n4216) );
  OAI222XL U1617 ( .A0(n318), .A1(n4185), .B0(n434), .B1(n1274), .C0(n320), 
        .C1(n1300), .Y(n4219) );
  INVX1 U1618 ( .A(n428), .Y(n427) );
  OAI222XL U1619 ( .A0(n1306), .A1(n1258), .B0(n4108), .B1(n427), .C0(n319), 
        .C1(n1290), .Y(n4128) );
  NOR2X1 U1620 ( .A(n808), .B(n319), .Y(n4000) );
  INVX1 U1621 ( .A(n4014), .Y(n1292) );
  INVX1 U1622 ( .A(n4051), .Y(n1304) );
  INVX1 U1623 ( .A(n260), .Y(n1303) );
  OAI21XL U1624 ( .A0(n320), .A1(n1253), .B0(n4151), .Y(n4214) );
  NOR2X1 U1625 ( .A(n290), .B(n425), .Y(n4069) );
  INVX1 U1626 ( .A(n4194), .Y(n1287) );
  NAND2X1 U1627 ( .A(n4017), .B(n319), .Y(n4093) );
  NOR2X1 U1628 ( .A(n1287), .B(n2947), .Y(n4233) );
  INVX1 U1629 ( .A(n4029), .Y(n1267) );
  OAI21XL U1630 ( .A0(n320), .A1(n1256), .B0(n1271), .Y(n4211) );
  AOI21X1 U1631 ( .A0(n3869), .A1(n3870), .B0(n3677), .Y(N3575) );
  NOR4X1 U1632 ( .A(n3909), .B(n3910), .C(n3911), .D(n3912), .Y(n3869) );
  NOR4X1 U1633 ( .A(n3871), .B(n3872), .C(n3873), .D(n3874), .Y(n3870) );
  NAND4X1 U1634 ( .A(n3935), .B(n3936), .C(n3937), .D(n3938), .Y(n3909) );
  AOI21X1 U1635 ( .A0(n3827), .A1(n3828), .B0(n3677), .Y(N3576) );
  NOR4X1 U1636 ( .A(n3849), .B(n3850), .C(n3851), .D(n3852), .Y(n3827) );
  NOR4X1 U1637 ( .A(n3829), .B(n3830), .C(n3831), .D(n3832), .Y(n3828) );
  NAND4X1 U1638 ( .A(n3865), .B(n3866), .C(n3867), .D(n3868), .Y(n3849) );
  AOI21X1 U1639 ( .A0(n3785), .A1(n3786), .B0(n3677), .Y(N3577) );
  NOR4X1 U1640 ( .A(n3807), .B(n3808), .C(n3809), .D(n3810), .Y(n3785) );
  NOR4X1 U1641 ( .A(n3787), .B(n3788), .C(n3789), .D(n3790), .Y(n3786) );
  NAND4X1 U1642 ( .A(n3823), .B(n3824), .C(n3825), .D(n3826), .Y(n3807) );
  AOI21X1 U1643 ( .A0(n3680), .A1(n3681), .B0(n3677), .Y(N3578) );
  NOR4X1 U1644 ( .A(n3733), .B(n3734), .C(n3735), .D(n3736), .Y(n3680) );
  NOR4X1 U1645 ( .A(n3682), .B(n3683), .C(n3684), .D(n3685), .Y(n3681) );
  NAND4X1 U1646 ( .A(n3773), .B(n3774), .C(n3775), .D(n3776), .Y(n3733) );
  NAND2X1 U1647 ( .A(n4069), .B(n260), .Y(n3972) );
  XOR3X2 U1648 ( .A(n312), .B(n306), .C(n294), .Y(f3_A_32[28]) );
  XOR3X2 U1649 ( .A(n311), .B(n305), .C(n293), .Y(f3_A_32[29]) );
  XOR3X2 U1650 ( .A(n317), .B(n16), .C(n304), .Y(f3_A_32[30]) );
  OR3XL U1651 ( .A(n3983), .B(n4063), .C(n3962), .Y(n4129) );
  AOI2BB1X1 U1652 ( .A0N(n4032), .A1N(n3983), .B0(n422), .Y(n4031) );
  NAND3BX1 U1653 ( .AN(n3963), .B(n1284), .C(n3985), .Y(n4079) );
  INVX1 U1654 ( .A(n4024), .Y(n1284) );
  BUFX3 U1655 ( .A(n1297), .Y(n290) );
  INVX1 U1656 ( .A(n4016), .Y(n1297) );
  OR3XL U1657 ( .A(n4044), .B(n3962), .C(n3990), .Y(n4232) );
  OR3XL U1658 ( .A(n4193), .B(n3988), .C(n4147), .Y(n4217) );
  INVX1 U1659 ( .A(n4224), .Y(n1252) );
  AOI21X1 U1660 ( .A0(n2946), .A1(n4137), .B0(n4214), .Y(n4224) );
  OAI222XL U1661 ( .A0(n427), .A1(n4173), .B0(n4179), .B1(n422), .C0(n290), 
        .C1(n1283), .Y(n4177) );
  OAI222XL U1662 ( .A0(n318), .A1(n3985), .B0(n1292), .B1(n1306), .C0(n320), 
        .C1(n1246), .Y(n3982) );
  OAI222XL U1663 ( .A0(n3957), .A1(n289), .B0(n1305), .B1(n1274), .C0(n3958), 
        .C1(n1251), .Y(n3956) );
  OAI222XL U1664 ( .A0(n1306), .A1(n1280), .B0(n318), .B1(n1274), .C0(n422), 
        .C1(n3958), .Y(n4170) );
  INVX1 U1665 ( .A(n4027), .Y(n1275) );
  OAI221XL U1666 ( .A0(n4107), .A1(n320), .B0(n4094), .B1(n429), .C0(n4108), 
        .Y(n4106) );
  OAI221XL U1667 ( .A0(n4051), .A1(n290), .B0(n434), .B1(n255), .C0(n4151), 
        .Y(n4148) );
  NOR2X1 U1668 ( .A(n289), .B(n319), .Y(n4003) );
  NAND2X1 U1669 ( .A(n3946), .B(n4051), .Y(n4151) );
  NOR2X1 U1670 ( .A(n425), .B(n319), .Y(n4083) );
  OAI211X1 U1671 ( .A0(n434), .A1(n429), .B0(n1256), .C0(n318), .Y(n4118) );
  NOR2X1 U1672 ( .A(n2946), .B(n434), .Y(n4105) );
  NOR2X1 U1673 ( .A(n426), .B(n2946), .Y(n4122) );
  INVX1 U1674 ( .A(n4158), .Y(n1259) );
  NOR2X1 U1675 ( .A(n290), .B(n318), .Y(n4132) );
  NAND4X1 U1676 ( .A(n3853), .B(n3854), .C(n3855), .D(n3856), .Y(n3852) );
  AOI22X1 U1677 ( .A0(n3747), .A1(n299), .B0(n3748), .B1(n295), .Y(n3853) );
  NAND4X1 U1678 ( .A(n3811), .B(n3812), .C(n3813), .D(n3814), .Y(n3810) );
  AOI22X1 U1679 ( .A0(n3747), .A1(n298), .B0(n3748), .B1(n294), .Y(n3811) );
  NAND4X1 U1680 ( .A(n3737), .B(n3738), .C(n3739), .D(n3740), .Y(n3736) );
  AOI22X1 U1681 ( .A0(n3747), .A1(n297), .B0(n3748), .B1(n293), .Y(n3737) );
  AOI21X1 U1682 ( .A0(n2946), .A1(n3960), .B0(n4147), .Y(n4087) );
  INVX1 U1683 ( .A(n4124), .Y(n1265) );
  OAI2BB1X1 U1684 ( .A0N(n3946), .A1N(n259), .B0(n4094), .Y(n3950) );
  OAI21XL U1685 ( .A0(n318), .A1(n1292), .B0(n1299), .Y(n4140) );
  AOI21X1 U1686 ( .A0(n1224), .A1(n4016), .B0(n4003), .Y(n4185) );
  AOI22X1 U1687 ( .A0(n3944), .A1(n1224), .B0(n260), .B1(n3946), .Y(n3943) );
  INVX1 U1688 ( .A(n4149), .Y(n1273) );
  OAI21XL U1689 ( .A0(n4067), .A1(n1293), .B0(n4068), .Y(n4064) );
  INVX1 U1690 ( .A(n4071), .Y(n1293) );
  OAI21XL U1691 ( .A0(n4069), .A1(n4070), .B0(n434), .Y(n4068) );
  INVX1 U1692 ( .A(n4011), .Y(n1281) );
  INVX1 U1693 ( .A(n4225), .Y(n1254) );
  OR2X2 U1694 ( .A(n4094), .B(n319), .Y(n3971) );
  NAND4BXL U1695 ( .AN(n3969), .B(n3970), .C(n3971), .D(n3972), .Y(n3968) );
  AOI21X1 U1696 ( .A0(n4082), .A1(n4010), .B0(n318), .Y(n4200) );
  AOI21X1 U1697 ( .A0(n4019), .A1(n4010), .B0(n318), .Y(n4166) );
  INVX1 U1698 ( .A(n4173), .Y(n1249) );
  INVX1 U1699 ( .A(n259), .Y(n1306) );
  OR2X2 U1700 ( .A(n4028), .B(n4193), .Y(n4213) );
  NOR2X1 U1701 ( .A(n319), .B(n434), .Y(n3965) );
  NOR2X1 U1702 ( .A(n426), .B(n318), .Y(n3944) );
  INVX1 U1703 ( .A(n302), .Y(n1119) );
  INVX1 U1704 ( .A(n300), .Y(n1111) );
  INVX1 U1705 ( .A(n293), .Y(n1051) );
  INVXL U1706 ( .A(n185), .Y(n788) );
  INVXL U1707 ( .A(n285), .Y(n796) );
  INVX1 U1708 ( .A(n306), .Y(n1230) );
  INVX1 U1709 ( .A(n307), .Y(n1229) );
  INVX1 U1710 ( .A(n303), .Y(n1233) );
  INVX1 U1711 ( .A(n304), .Y(n1232) );
  INVXL U1712 ( .A(n280), .Y(n743) );
  INVX1 U1713 ( .A(n298), .Y(n1103) );
  INVX1 U1714 ( .A(n301), .Y(n1115) );
  INVX1 U1715 ( .A(n296), .Y(n1095) );
  INVX1 U1716 ( .A(n299), .Y(n1106) );
  INVX1 U1717 ( .A(n308), .Y(n1228) );
  INVX1 U1718 ( .A(n305), .Y(n1231) );
  INVX1 U1719 ( .A(n294), .Y(n1086) );
  INVX1 U1720 ( .A(n297), .Y(n1098) );
  INVX1 U1721 ( .A(n295), .Y(n1090) );
  INVXL U1722 ( .A(next_E[19]), .Y(n731) );
  INVXL U1723 ( .A(next_E[17]), .Y(n737) );
  MX2X1 U1724 ( .A(SHA256_result[159]), .B(SHA256_result[191]), .S0(n438), .Y(
        mux1[31]) );
  NAND2XL U1725 ( .A(next_E[28]), .B(n339), .Y(n708) );
  NAND2XL U1726 ( .A(next_E[24]), .B(n339), .Y(n718) );
  NAND2BXL U1727 ( .AN(n330), .B(n70), .Y(n710) );
  NAND2BXL U1728 ( .AN(n334), .B(n198), .Y(n723) );
  NAND2BXL U1729 ( .AN(n330), .B(next_E[23]), .Y(n720) );
  NAND2X1 U1730 ( .A(H4[29]), .B(n205), .Y(n702) );
  NAND2X1 U1731 ( .A(N934), .B(n807), .Y(n610) );
  OAI221XL U1732 ( .A0(n287), .A1(n631), .B0(n112), .B1(n795), .C0(n630), .Y(
        n4424) );
  INVX1 U1733 ( .A(N924), .Y(n631) );
  NAND2XL U1734 ( .A(n321), .B(SHA256_result[83]), .Y(n630) );
  INVX1 U1735 ( .A(N926), .Y(n627) );
  NAND2XL U1736 ( .A(n321), .B(SHA256_result[85]), .Y(n626) );
  OAI221XL U1737 ( .A0(n287), .A1(n629), .B0(n1369), .B1(n334), .C0(n628), .Y(
        n4423) );
  INVX1 U1738 ( .A(N925), .Y(n629) );
  NAND2XL U1739 ( .A(n321), .B(SHA256_result[84]), .Y(n628) );
  OAI221XL U1740 ( .A0(n287), .A1(n636), .B0(n1367), .B1(n333), .C0(n635), .Y(
        n4426) );
  INVX1 U1741 ( .A(N922), .Y(n636) );
  NAND2XL U1742 ( .A(n321), .B(SHA256_result[81]), .Y(n635) );
  OAI221XL U1743 ( .A0(n798), .A1(n482), .B0(n1392), .B1(n332), .C0(n481), .Y(
        n4295) );
  INVX1 U1744 ( .A(N860), .Y(n482) );
  OAI221XL U1745 ( .A0(n287), .A1(n484), .B0(n1391), .B1(n335), .C0(n483), .Y(
        n4296) );
  INVX1 U1746 ( .A(N859), .Y(n484) );
  INVX1 U1747 ( .A(N861), .Y(n480) );
  OAI221XL U1748 ( .A0(n287), .A1(n455), .B0(n1401), .B1(n335), .C0(n454), .Y(
        n4285) );
  INVX1 U1749 ( .A(N870), .Y(n455) );
  OAI221XL U1750 ( .A0(n287), .A1(n557), .B0(n1375), .B1(n333), .C0(n556), .Y(
        n4392) );
  INVX1 U1751 ( .A(N892), .Y(n557) );
  NAND2XL U1752 ( .A(n321), .B(SHA256_result[51]), .Y(n556) );
  OAI221XL U1753 ( .A0(n798), .A1(n529), .B0(n1386), .B1(n331), .C0(n528), .Y(
        n4381) );
  INVX1 U1754 ( .A(N903), .Y(n529) );
  INVX1 U1755 ( .A(N895), .Y(n551) );
  NAND2XL U1756 ( .A(n322), .B(SHA256_result[54]), .Y(n550) );
  OAI221XL U1757 ( .A0(n287), .A1(n553), .B0(n1377), .B1(n333), .C0(n552), .Y(
        n4390) );
  INVX1 U1758 ( .A(N894), .Y(n553) );
  NAND2XL U1759 ( .A(n322), .B(SHA256_result[53]), .Y(n552) );
  OAI221XL U1760 ( .A0(n287), .A1(n555), .B0(n1376), .B1(n335), .C0(n554), .Y(
        n4391) );
  INVX1 U1761 ( .A(N893), .Y(n555) );
  NAND2XL U1762 ( .A(n322), .B(SHA256_result[52]), .Y(n554) );
  OAI221XL U1763 ( .A0(n798), .A1(n531), .B0(n1385), .B1(n332), .C0(n530), .Y(
        n4382) );
  INVX1 U1764 ( .A(N902), .Y(n531) );
  OAI221XL U1765 ( .A0(n798), .A1(n463), .B0(n1398), .B1(n333), .C0(n462), .Y(
        n4288) );
  INVX1 U1766 ( .A(N867), .Y(n463) );
  OAI221XL U1767 ( .A0(n798), .A1(n486), .B0(n1390), .B1(n335), .C0(n485), .Y(
        n4297) );
  INVX1 U1768 ( .A(N858), .Y(n486) );
  OAI221XL U1769 ( .A0(n798), .A1(n488), .B0(n1389), .B1(n335), .C0(n487), .Y(
        n4298) );
  INVX1 U1770 ( .A(N857), .Y(n488) );
  OAI221XL U1771 ( .A0(n287), .A1(n559), .B0(n1374), .B1(n333), .C0(n558), .Y(
        n4393) );
  INVX1 U1772 ( .A(N891), .Y(n559) );
  NAND2XL U1773 ( .A(n321), .B(SHA256_result[50]), .Y(n558) );
  OAI221XL U1774 ( .A0(n798), .A1(n527), .B0(n1387), .B1(n335), .C0(n526), .Y(
        n4380) );
  INVX1 U1775 ( .A(N904), .Y(n527) );
  NAND2X1 U1776 ( .A(n322), .B(SHA256_result[63]), .Y(n526) );
  XOR3X2 U1777 ( .A(n222), .B(n309), .C(n298), .Y(f3_A_32[13]) );
  XOR3X2 U1778 ( .A(n292), .B(SHA256_result[113]), .C(SHA256_result[118]), .Y(
        f4_E_32[11]) );
  OAI211X1 U1779 ( .A0(n331), .A1(n137), .B0(n649), .C0(n648), .Y(n4432) );
  NAND2X1 U1780 ( .A(N916), .B(n807), .Y(n649) );
  NAND2XL U1781 ( .A(SHA256_result[74]), .B(n323), .Y(n652) );
  NAND2X1 U1782 ( .A(N915), .B(n807), .Y(n651) );
  NAND2X1 U1783 ( .A(N913), .B(n807), .Y(n657) );
  OAI211X1 U1784 ( .A0(n407), .A1(n112), .B0(n419), .C0(n3309), .Y(n4519) );
  NAND2X1 U1785 ( .A(H4[19]), .B(n205), .Y(n3309) );
  OAI211X1 U1786 ( .A0(n335), .A1(n746), .B0(n642), .C0(n641), .Y(n4429) );
  NAND2X1 U1787 ( .A(N919), .B(n807), .Y(n642) );
  NAND2X1 U1788 ( .A(H4[14]), .B(n205), .Y(n3312) );
  NAND2X1 U1789 ( .A(N908), .B(n807), .Y(n672) );
  OAI211X1 U1790 ( .A0(n795), .A1(n763), .B0(n655), .C0(n654), .Y(n4434) );
  NAND2X1 U1791 ( .A(N914), .B(n807), .Y(n654) );
  NAND2X1 U1792 ( .A(H4[9]), .B(n205), .Y(n3314) );
  OAI211X1 U1793 ( .A0(n410), .A1(n784), .B0(n3318), .C0(n419), .Y(n4535) );
  NAND2X1 U1794 ( .A(H4[3]), .B(n205), .Y(n3318) );
  NAND2X1 U1795 ( .A(N918), .B(n807), .Y(n644) );
  OAI211X1 U1796 ( .A0(n1312), .A1(n24), .B0(n949), .C0(n948), .Y(n4658) );
  AOI21XL U1797 ( .A0(SHA256_result[168]), .A1(n399), .B0(n389), .Y(n948) );
  OAI211X1 U1798 ( .A0(n1316), .A1(n27), .B0(n930), .C0(n929), .Y(n4652) );
  OAI211X1 U1799 ( .A0(n1314), .A1(n22), .B0(n935), .C0(n934), .Y(n4654) );
  AOI21XL U1800 ( .A0(SHA256_result[172]), .A1(n399), .B0(n389), .Y(n934) );
  AOI21XL U1801 ( .A0(SHA256_result[166]), .A1(n399), .B0(n389), .Y(n955) );
  AOI21XL U1802 ( .A0(SHA256_result[165]), .A1(n399), .B0(n389), .Y(n958) );
  OAI211XL U1803 ( .A0(n795), .A1(n684), .B0(n495), .C0(n494), .Y(n4301) );
  NAND2X1 U1804 ( .A(N854), .B(n807), .Y(n494) );
  OAI211XL U1805 ( .A0(n331), .A1(n686), .B0(n497), .C0(n496), .Y(n4302) );
  NAND2X1 U1806 ( .A(N853), .B(n807), .Y(n496) );
  OAI211XL U1807 ( .A0(n406), .A1(n686), .B0(n3197), .C0(n419), .Y(n4367) );
  NAND2XL U1808 ( .A(SHA256_result[45]), .B(n323), .Y(n573) );
  OAI211XL U1809 ( .A0(n406), .A1(n683), .B0(n3182), .C0(n419), .Y(n4334) );
  NAND2X1 U1810 ( .A(N921), .B(n807), .Y(n638) );
  AOI21XL U1811 ( .A0(n343), .A1(SHA256_result[80]), .B0(n328), .Y(n637) );
  NAND2X1 U1812 ( .A(N927), .B(n807), .Y(n624) );
  NAND2XL U1813 ( .A(n321), .B(SHA256_result[86]), .Y(n625) );
  NAND2X1 U1814 ( .A(N928), .B(n807), .Y(n622) );
  NAND2XL U1815 ( .A(n321), .B(SHA256_result[87]), .Y(n623) );
  OAI211X1 U1816 ( .A0(n1340), .A1(n24), .B0(n828), .C0(n827), .Y(n4610) );
  AOI21X1 U1817 ( .A0(n399), .A1(SHA256_result[152]), .B0(n390), .Y(n827) );
  OAI211X1 U1818 ( .A0(n1332), .A1(n21), .B0(n844), .C0(n843), .Y(n4618) );
  AOI21X1 U1819 ( .A0(n399), .A1(SHA256_result[144]), .B0(n390), .Y(n843) );
  NAND2X1 U1820 ( .A(N1000), .B(n124), .Y(n895) );
  AOI21X1 U1821 ( .A0(n399), .A1(SHA256_result[159]), .B0(n387), .Y(n894) );
  OAI211X1 U1822 ( .A0(n409), .A1(n1367), .B0(n419), .C0(n3311), .Y(n4521) );
  NAND2X1 U1823 ( .A(H4[17]), .B(n205), .Y(n3311) );
  OAI211X1 U1824 ( .A0(n332), .A1(n145), .B0(n647), .C0(n646), .Y(n4431) );
  NAND2XL U1825 ( .A(SHA256_result[76]), .B(n323), .Y(n647) );
  NAND2X1 U1826 ( .A(N917), .B(n807), .Y(n646) );
  NAND2X1 U1827 ( .A(H4[12]), .B(n205), .Y(n3313) );
  OAI211X1 U1828 ( .A0(n335), .A1(n82), .B0(n590), .C0(n589), .Y(n4405) );
  NAND2X1 U1829 ( .A(N879), .B(n807), .Y(n589) );
  OAI211X1 U1830 ( .A0(n332), .A1(n668), .B0(n595), .C0(n594), .Y(n4407) );
  NAND2X1 U1831 ( .A(N877), .B(n807), .Y(n594) );
  NAND2X1 U1832 ( .A(H4[24]), .B(n205), .Y(n3308) );
  NAND2X1 U1833 ( .A(H4[28]), .B(n205), .Y(n3307) );
  NAND2X1 U1834 ( .A(N935), .B(n807), .Y(n608) );
  NAND2X1 U1835 ( .A(H4[30]), .B(n205), .Y(n3306) );
  NAND2X1 U1836 ( .A(N1018), .B(n370), .Y(n923) );
  AOI21X1 U1837 ( .A0(n399), .A1(SHA256_result[177]), .B0(n385), .Y(n922) );
  NAND2X1 U1838 ( .A(N1022), .B(n124), .Y(n915) );
  AOI21X1 U1839 ( .A0(n399), .A1(SHA256_result[181]), .B0(n388), .Y(n914) );
  NAND2X1 U1840 ( .A(N1016), .B(n372), .Y(n928) );
  AOI21X1 U1841 ( .A0(n399), .A1(SHA256_result[173]), .B0(n389), .Y(n931) );
  OAI211X1 U1842 ( .A0(n1341), .A1(n25), .B0(n824), .C0(n823), .Y(n4608) );
  AOI21X1 U1843 ( .A0(n399), .A1(SHA256_result[154]), .B0(n390), .Y(n823) );
  OAI211X1 U1844 ( .A0(n1335), .A1(n22), .B0(n838), .C0(n837), .Y(n4615) );
  AOI21X1 U1845 ( .A0(n399), .A1(SHA256_result[147]), .B0(n390), .Y(n837) );
  OAI211X1 U1846 ( .A0(n1334), .A1(n22), .B0(n840), .C0(n839), .Y(n4616) );
  AOI21X1 U1847 ( .A0(n399), .A1(SHA256_result[146]), .B0(n390), .Y(n839) );
  OAI211X1 U1848 ( .A0(n1333), .A1(n25), .B0(n842), .C0(n841), .Y(n4617) );
  AOI21X1 U1849 ( .A0(n399), .A1(SHA256_result[145]), .B0(n390), .Y(n841) );
  NAND2X1 U1850 ( .A(N1030), .B(n371), .Y(n899) );
  AOI21X1 U1851 ( .A0(n399), .A1(SHA256_result[189]), .B0(n388), .Y(n898) );
  NAND2X1 U1852 ( .A(N1029), .B(n372), .Y(n901) );
  AOI21X1 U1853 ( .A0(n399), .A1(SHA256_result[188]), .B0(n385), .Y(n900) );
  OAI211X1 U1854 ( .A0(n1313), .A1(n28), .B0(n946), .C0(n945), .Y(n4657) );
  AOI21XL U1855 ( .A0(SHA256_result[169]), .A1(n399), .B0(n389), .Y(n945) );
  NAND2X1 U1856 ( .A(N1023), .B(n369), .Y(n913) );
  AOI21X1 U1857 ( .A0(n399), .A1(SHA256_result[182]), .B0(n387), .Y(n912) );
  OAI211X1 U1858 ( .A0(n1344), .A1(n24), .B0(n818), .C0(n817), .Y(n4605) );
  NAND2X1 U1859 ( .A(N998), .B(n124), .Y(n818) );
  OAI211X1 U1860 ( .A0(n1338), .A1(n28), .B0(n832), .C0(n831), .Y(n4612) );
  AOI21X1 U1861 ( .A0(n399), .A1(SHA256_result[150]), .B0(n388), .Y(n831) );
  OAI211X1 U1862 ( .A0(n1331), .A1(n26), .B0(n846), .C0(n845), .Y(n4619) );
  AOI21X1 U1863 ( .A0(n399), .A1(SHA256_result[143]), .B0(n390), .Y(n845) );
  OAI211X1 U1864 ( .A0(n1330), .A1(n23), .B0(n848), .C0(n847), .Y(n4620) );
  AOI21X1 U1865 ( .A0(n399), .A1(SHA256_result[142]), .B0(n390), .Y(n847) );
  OAI211X1 U1866 ( .A0(n406), .A1(n1319), .B0(n419), .C0(n3277), .Y(n4457) );
  NAND2X1 U1867 ( .A(H1[18]), .B(n205), .Y(n3277) );
  OAI211X1 U1868 ( .A0(n410), .A1(n1318), .B0(n419), .C0(n3278), .Y(n4458) );
  NAND2X1 U1869 ( .A(H1[17]), .B(n205), .Y(n3278) );
  OAI211X1 U1870 ( .A0(n408), .A1(n1322), .B0(n419), .C0(n3276), .Y(n4454) );
  NAND2X1 U1871 ( .A(H1[21]), .B(n205), .Y(n3276) );
  OAI211X1 U1872 ( .A0(n412), .A1(n1235), .B0(n419), .C0(n3272), .Y(n4448) );
  NAND2X1 U1873 ( .A(H1[27]), .B(n205), .Y(n3272) );
  OAI211X1 U1874 ( .A0(n412), .A1(n1341), .B0(n419), .C0(n3290), .Y(n4480) );
  NAND2X1 U1875 ( .A(H2[26]), .B(n205), .Y(n3290) );
  OAI211X1 U1876 ( .A0(n1244), .A1(n1335), .B0(n419), .C0(n3293), .Y(n4487) );
  NAND2X1 U1877 ( .A(H2[19]), .B(n205), .Y(n3293) );
  OAI211X1 U1878 ( .A0(n408), .A1(n1334), .B0(n419), .C0(n3294), .Y(n4488) );
  NAND2X1 U1879 ( .A(H2[18]), .B(n205), .Y(n3294) );
  OAI211X1 U1880 ( .A0(n412), .A1(n1333), .B0(n419), .C0(n3295), .Y(n4489) );
  NAND2X1 U1881 ( .A(H2[17]), .B(n205), .Y(n3295) );
  OAI211X1 U1882 ( .A0(n406), .A1(n1237), .B0(n419), .C0(n3270), .Y(n4446) );
  NAND2X1 U1883 ( .A(H1[29]), .B(n205), .Y(n3270) );
  OAI211X1 U1884 ( .A0(n412), .A1(n1236), .B0(n419), .C0(n3271), .Y(n4447) );
  NAND2X1 U1885 ( .A(H1[28]), .B(n205), .Y(n3271) );
  OAI211X1 U1886 ( .A0(n408), .A1(n1323), .B0(n419), .C0(n3275), .Y(n4453) );
  NAND2X1 U1887 ( .A(H1[22]), .B(n205), .Y(n3275) );
  OAI211X1 U1888 ( .A0(n406), .A1(n1344), .B0(n419), .C0(n3287), .Y(n4477) );
  NAND2X1 U1889 ( .A(H2[29]), .B(n205), .Y(n3287) );
  OAI211X1 U1890 ( .A0(n409), .A1(n1338), .B0(n419), .C0(n3291), .Y(n4484) );
  NAND2X1 U1891 ( .A(H2[22]), .B(n205), .Y(n3291) );
  OAI211X1 U1892 ( .A0(n408), .A1(n1342), .B0(n419), .C0(n3289), .Y(n4479) );
  NAND2X1 U1893 ( .A(H2[27]), .B(n205), .Y(n3289) );
  OAI211X1 U1894 ( .A0(n1244), .A1(n1343), .B0(n419), .C0(n3288), .Y(n4478) );
  NAND2X1 U1895 ( .A(H2[28]), .B(n205), .Y(n3288) );
  OAI211X1 U1896 ( .A0(n408), .A1(n1337), .B0(n419), .C0(n3292), .Y(n4485) );
  NAND2X1 U1897 ( .A(H2[21]), .B(n205), .Y(n3292) );
  OAI211X1 U1898 ( .A0(n25), .A1(n933), .B0(n852), .C0(n851), .Y(n4622) );
  AOI21X1 U1899 ( .A0(n399), .A1(SHA256_result[140]), .B0(n390), .Y(n851) );
  OAI211X1 U1900 ( .A0(n409), .A1(n1398), .B0(n419), .C0(n3189), .Y(n4353) );
  NAND2X1 U1901 ( .A(H6[26]), .B(n205), .Y(n3189) );
  OAI211X1 U1902 ( .A0(n408), .A1(n1390), .B0(n419), .C0(n3193), .Y(n4362) );
  NAND2X1 U1903 ( .A(H6[17]), .B(n205), .Y(n3193) );
  OAI211X1 U1904 ( .A0(n412), .A1(n1389), .B0(n419), .C0(n3194), .Y(n4363) );
  NAND2X1 U1905 ( .A(H6[16]), .B(n205), .Y(n3194) );
  NAND2X1 U1906 ( .A(N912), .B(n807), .Y(n660) );
  OAI211X1 U1907 ( .A0(n408), .A1(n1374), .B0(n419), .C0(n3179), .Y(n4329) );
  NAND2X1 U1908 ( .A(H5[18]), .B(n205), .Y(n3179) );
  OAI211X1 U1909 ( .A0(n1244), .A1(n1387), .B0(n419), .C0(n3174), .Y(n4316) );
  NAND2X1 U1910 ( .A(H5[31]), .B(n205), .Y(n3174) );
  AOI21X1 U1911 ( .A0(SHA256_result[213]), .A1(n399), .B0(n389), .Y(n1001) );
  OAI211X1 U1912 ( .A0(n334), .A1(n743), .B0(n640), .C0(n639), .Y(n4428) );
  NAND2X1 U1913 ( .A(N920), .B(n807), .Y(n639) );
  NAND2XL U1914 ( .A(n323), .B(SHA256_result[79]), .Y(n640) );
  OAI211X1 U1915 ( .A0(n407), .A1(n1154), .B0(n3513), .C0(n419), .Y(n4723) );
  NAND2X1 U1916 ( .A(H0[10]), .B(n205), .Y(n3513) );
  OAI211X1 U1917 ( .A0(n410), .A1(n1158), .B0(n3514), .C0(n419), .Y(n4724) );
  NAND2X1 U1918 ( .A(H0[9]), .B(n205), .Y(n3514) );
  AOI21X1 U1919 ( .A0(n399), .A1(SHA256_result[220]), .B0(n389), .Y(n984) );
  OAI211X1 U1920 ( .A0(n411), .A1(n1106), .B0(n3507), .C0(n419), .Y(n4708) );
  NAND2X1 U1921 ( .A(H0[25]), .B(n205), .Y(n3507) );
  OAI211X1 U1922 ( .A0(n406), .A1(n1188), .B0(n3518), .C0(n419), .Y(n4731) );
  NAND2X1 U1923 ( .A(H0[2]), .B(n205), .Y(n3518) );
  AOI21X1 U1924 ( .A0(n399), .A1(SHA256_result[221]), .B0(n389), .Y(n982) );
  NAND2X1 U1925 ( .A(N907), .B(n807), .Y(n674) );
  NAND2XL U1926 ( .A(n83), .B(n322), .Y(n663) );
  NAND2X1 U1927 ( .A(N911), .B(n807), .Y(n662) );
  NAND2XL U1928 ( .A(n129), .B(n323), .Y(n666) );
  NAND2X1 U1929 ( .A(N910), .B(n807), .Y(n665) );
  NAND2XL U1930 ( .A(SHA256_result[68]), .B(n323), .Y(n670) );
  NAND2X1 U1931 ( .A(N909), .B(n807), .Y(n669) );
  NAND2X1 U1932 ( .A(N906), .B(n807), .Y(n676) );
  NAND2X1 U1933 ( .A(N905), .B(n807), .Y(n679) );
  AOI21XL U1934 ( .A0(n96), .A1(n399), .B0(n390), .Y(n1048) );
  NAND2X1 U1935 ( .A(N880), .B(n807), .Y(n587) );
  OAI211XL U1936 ( .A0(n332), .A1(n206), .B0(n597), .C0(n596), .Y(n4408) );
  NAND2X1 U1937 ( .A(N876), .B(n807), .Y(n597) );
  NAND2X1 U1938 ( .A(N887), .B(n807), .Y(n570) );
  NAND2X1 U1939 ( .A(N884), .B(n807), .Y(n577) );
  NAND2X1 U1940 ( .A(N881), .B(n807), .Y(n585) );
  NAND2X1 U1941 ( .A(N874), .B(n807), .Y(n602) );
  OAI211XL U1942 ( .A0(n331), .A1(n699), .B0(n604), .C0(n603), .Y(n4411) );
  NAND2X1 U1943 ( .A(N873), .B(n807), .Y(n604) );
  OAI211XL U1944 ( .A0(n334), .A1(n162), .B0(n523), .C0(n522), .Y(n4313) );
  NAND2X1 U1945 ( .A(N883), .B(n807), .Y(n579) );
  NAND2X1 U1946 ( .A(N882), .B(n807), .Y(n582) );
  NAND2X1 U1947 ( .A(N875), .B(n807), .Y(n599) );
  AOI21X1 U1948 ( .A0(SHA256_result[207]), .A1(n399), .B0(n390), .Y(n1013) );
  OAI211X1 U1949 ( .A0(n1225), .A1(n23), .B0(n1018), .C0(n1017), .Y(n4685) );
  AOI21XL U1950 ( .A0(SHA256_result[205]), .A1(n399), .B0(n390), .Y(n1017) );
  OAI211XL U1951 ( .A0(n332), .A1(n682), .B0(n493), .C0(n492), .Y(n4300) );
  NAND2X1 U1952 ( .A(N855), .B(n807), .Y(n493) );
  OAI211XL U1953 ( .A0(n333), .A1(n688), .B0(n499), .C0(n498), .Y(n4303) );
  OAI211XL U1954 ( .A0(n335), .A1(n160), .B0(n501), .C0(n500), .Y(n4304) );
  OAI211XL U1955 ( .A0(n332), .A1(n166), .B0(n503), .C0(n502), .Y(n4305) );
  OAI211XL U1956 ( .A0(n330), .A1(n183), .B0(n505), .C0(n504), .Y(n4306) );
  OAI211XL U1957 ( .A0(n335), .A1(n692), .B0(n507), .C0(n506), .Y(n4307) );
  OAI211XL U1958 ( .A0(n333), .A1(n1206), .B0(n510), .C0(n509), .Y(n4308) );
  OAI211XL U1959 ( .A0(n335), .A1(n1208), .B0(n513), .C0(n512), .Y(n4309) );
  OAI211XL U1960 ( .A0(n795), .A1(n89), .B0(n517), .C0(n516), .Y(n4311) );
  OAI211X1 U1961 ( .A0(n408), .A1(n1427), .B0(n419), .C0(n3118), .Y(n4253) );
  INVX1 U1962 ( .A(SHA256_result[30]), .Y(n1427) );
  NAND2X1 U1963 ( .A(H7[30]), .B(n205), .Y(n3118) );
  OAI211X1 U1964 ( .A0(n409), .A1(n1425), .B0(n419), .C0(n3119), .Y(n4255) );
  INVX1 U1965 ( .A(SHA256_result[28]), .Y(n1425) );
  NAND2X1 U1966 ( .A(H7[28]), .B(n205), .Y(n3119) );
  OAI211X1 U1967 ( .A0(n406), .A1(n1424), .B0(n419), .C0(n3120), .Y(n4256) );
  INVX1 U1968 ( .A(SHA256_result[27]), .Y(n1424) );
  NAND2X1 U1969 ( .A(H7[27]), .B(n205), .Y(n3120) );
  OAI211X1 U1970 ( .A0(n411), .A1(n1422), .B0(n419), .C0(n3121), .Y(n4258) );
  INVX1 U1971 ( .A(SHA256_result[25]), .Y(n1422) );
  NAND2X1 U1972 ( .A(H7[25]), .B(n205), .Y(n3121) );
  OAI211X1 U1973 ( .A0(n412), .A1(n1421), .B0(n419), .C0(n3122), .Y(n4259) );
  INVX1 U1974 ( .A(SHA256_result[24]), .Y(n1421) );
  NAND2X1 U1975 ( .A(H7[24]), .B(n205), .Y(n3122) );
  OAI211X1 U1976 ( .A0(n406), .A1(n1420), .B0(n419), .C0(n3123), .Y(n4260) );
  INVX1 U1977 ( .A(SHA256_result[23]), .Y(n1420) );
  NAND2X1 U1978 ( .A(H7[23]), .B(n205), .Y(n3123) );
  OAI211X1 U1979 ( .A0(n409), .A1(n1419), .B0(n419), .C0(n3124), .Y(n4261) );
  INVX1 U1980 ( .A(SHA256_result[22]), .Y(n1419) );
  NAND2X1 U1981 ( .A(H7[22]), .B(n205), .Y(n3124) );
  OAI211X1 U1982 ( .A0(n408), .A1(n1418), .B0(n419), .C0(n3125), .Y(n4262) );
  INVX1 U1983 ( .A(SHA256_result[21]), .Y(n1418) );
  NAND2X1 U1984 ( .A(H7[21]), .B(n205), .Y(n3125) );
  INVX1 U1985 ( .A(SHA256_result[15]), .Y(n1412) );
  INVX1 U1986 ( .A(SHA256_result[14]), .Y(n1411) );
  OAI211X1 U1987 ( .A0(n408), .A1(n1400), .B0(n419), .C0(n3187), .Y(n4351) );
  OAI211X1 U1988 ( .A0(n407), .A1(n1399), .B0(n419), .C0(n3188), .Y(n4352) );
  OAI211X1 U1989 ( .A0(n410), .A1(n1397), .B0(n419), .C0(n3190), .Y(n4354) );
  OAI211X1 U1990 ( .A0(n406), .A1(n120), .B0(n419), .C0(n3191), .Y(n4355) );
  NAND2X1 U1991 ( .A(H6[24]), .B(n205), .Y(n3191) );
  OAI211X1 U1992 ( .A0(n407), .A1(n1396), .B0(n419), .C0(n3192), .Y(n4356) );
  INVXL U1993 ( .A(SHA256_result[55]), .Y(n1396) );
  NAND2X1 U1994 ( .A(H6[23]), .B(n205), .Y(n3192) );
  INVXL U1995 ( .A(SHA256_result[47]), .Y(n1388) );
  OAI211XL U1996 ( .A0(n412), .A1(n682), .B0(n3196), .C0(n419), .Y(n4365) );
  OAI211XL U1997 ( .A0(n407), .A1(n688), .B0(n3198), .C0(n419), .Y(n4368) );
  OAI211XL U1998 ( .A0(n412), .A1(n183), .B0(n3199), .C0(n419), .Y(n4371) );
  OAI211XL U1999 ( .A0(n409), .A1(n692), .B0(n3200), .C0(n419), .Y(n4372) );
  OAI211XL U2000 ( .A0(n412), .A1(n1208), .B0(n3201), .C0(n419), .Y(n4374) );
  OAI211XL U2001 ( .A0(n409), .A1(n89), .B0(n3202), .C0(n419), .Y(n4376) );
  OAI211X1 U2002 ( .A0(n409), .A1(n1384), .B0(n419), .C0(n3175), .Y(n4319) );
  OAI211X1 U2003 ( .A0(n1244), .A1(n1383), .B0(n419), .C0(n3176), .Y(n4320) );
  OAI211X1 U2004 ( .A0(n411), .A1(n1381), .B0(n419), .C0(n3177), .Y(n4322) );
  OAI211X1 U2005 ( .A0(n407), .A1(n1380), .B0(n419), .C0(n3178), .Y(n4323) );
  INVX1 U2006 ( .A(n31), .Y(n1380) );
  NAND2X1 U2007 ( .A(H5[24]), .B(n205), .Y(n3178) );
  OAI211X1 U2008 ( .A0(n412), .A1(n1372), .B0(n419), .C0(n3180), .Y(n4331) );
  INVXL U2009 ( .A(SHA256_result[80]), .Y(n1372) );
  NAND2X1 U2010 ( .A(H5[16]), .B(n205), .Y(n3180) );
  OAI211XL U2011 ( .A0(n411), .A1(n681), .B0(n3181), .C0(n419), .Y(n4333) );
  OAI211XL U2012 ( .A0(n412), .A1(n687), .B0(n3183), .C0(n419), .Y(n4336) );
  OAI211XL U2013 ( .A0(n407), .A1(n206), .B0(n3185), .C0(n419), .Y(n4344) );
  OAI211X1 U2014 ( .A0(n408), .A1(n1368), .B0(n419), .C0(n3310), .Y(n4520) );
  OAI211X1 U2015 ( .A0(n412), .A1(n135), .B0(n3315), .C0(n419), .Y(n4532) );
  NAND2X1 U2016 ( .A(H4[6]), .B(n205), .Y(n3315) );
  OAI211X1 U2017 ( .A0(n408), .A1(n148), .B0(n3316), .C0(n419), .Y(n4533) );
  NAND2X1 U2018 ( .A(H4[5]), .B(n205), .Y(n3316) );
  OAI211X1 U2019 ( .A0(n407), .A1(n780), .B0(n3317), .C0(n419), .Y(n4534) );
  NAND2X1 U2020 ( .A(H4[4]), .B(n205), .Y(n3317) );
  OAI211X1 U2021 ( .A0(n407), .A1(n788), .B0(n3319), .C0(n419), .Y(n4536) );
  NAND2X1 U2022 ( .A(H4[2]), .B(n205), .Y(n3319) );
  OAI211X1 U2023 ( .A0(n412), .A1(n156), .B0(n3320), .C0(n419), .Y(n4537) );
  NAND2X1 U2024 ( .A(H4[1]), .B(n205), .Y(n3320) );
  OAI211X1 U2025 ( .A0(n411), .A1(n796), .B0(n3321), .C0(n419), .Y(n4538) );
  NAND2X1 U2026 ( .A(H4[0]), .B(n205), .Y(n3321) );
  OAI211X1 U2027 ( .A0(n410), .A1(n1365), .B0(n419), .C0(n3381), .Y(n4573) );
  INVX1 U2028 ( .A(SHA256_result[157]), .Y(n1365) );
  NAND2X1 U2029 ( .A(H3[29]), .B(n205), .Y(n3381) );
  OAI211X1 U2030 ( .A0(n410), .A1(n1362), .B0(n419), .C0(n3382), .Y(n4576) );
  INVX1 U2031 ( .A(SHA256_result[154]), .Y(n1362) );
  NAND2X1 U2032 ( .A(H3[26]), .B(n205), .Y(n3382) );
  OAI211X1 U2033 ( .A0(n407), .A1(n1360), .B0(n419), .C0(n3383), .Y(n4578) );
  INVX1 U2034 ( .A(SHA256_result[152]), .Y(n1360) );
  NAND2X1 U2035 ( .A(H3[24]), .B(n205), .Y(n3383) );
  OAI211X1 U2036 ( .A0(n408), .A1(n1358), .B0(n419), .C0(n3384), .Y(n4580) );
  INVX1 U2037 ( .A(SHA256_result[150]), .Y(n1358) );
  NAND2X1 U2038 ( .A(H3[22]), .B(n205), .Y(n3384) );
  OAI211X1 U2039 ( .A0(n408), .A1(n1355), .B0(n419), .C0(n3385), .Y(n4583) );
  INVX1 U2040 ( .A(SHA256_result[147]), .Y(n1355) );
  NAND2X1 U2041 ( .A(H3[19]), .B(n205), .Y(n3385) );
  OAI211X1 U2042 ( .A0(n408), .A1(n1354), .B0(n419), .C0(n3386), .Y(n4584) );
  INVX1 U2043 ( .A(SHA256_result[146]), .Y(n1354) );
  NAND2X1 U2044 ( .A(H3[18]), .B(n205), .Y(n3386) );
  OAI211X1 U2045 ( .A0(n406), .A1(n1353), .B0(n419), .C0(n3387), .Y(n4585) );
  INVX1 U2046 ( .A(SHA256_result[145]), .Y(n1353) );
  NAND2X1 U2047 ( .A(H3[17]), .B(n205), .Y(n3387) );
  OAI211X1 U2048 ( .A0(n406), .A1(n1352), .B0(n419), .C0(n3388), .Y(n4586) );
  INVX1 U2049 ( .A(SHA256_result[144]), .Y(n1352) );
  NAND2X1 U2050 ( .A(H3[16]), .B(n205), .Y(n3388) );
  INVX1 U2051 ( .A(SHA256_result[143]), .Y(n1351) );
  INVX1 U2052 ( .A(SHA256_result[142]), .Y(n1350) );
  INVX1 U2053 ( .A(SHA256_result[140]), .Y(n1348) );
  OAI211X1 U2054 ( .A0(n407), .A1(n1346), .B0(n419), .C0(n3380), .Y(n4571) );
  INVX1 U2055 ( .A(SHA256_result[159]), .Y(n1346) );
  NAND2X1 U2056 ( .A(H3[31]), .B(n205), .Y(n3380) );
  OAI211X1 U2057 ( .A0(n406), .A1(n1327), .B0(n419), .C0(n3269), .Y(n4444) );
  INVX1 U2058 ( .A(SHA256_result[223]), .Y(n1327) );
  NAND2X1 U2059 ( .A(H1[31]), .B(n205), .Y(n3269) );
  OAI211X1 U2060 ( .A0(n406), .A1(n1326), .B0(n419), .C0(n3273), .Y(n4450) );
  OAI211X1 U2061 ( .A0(n407), .A1(n1325), .B0(n419), .C0(n3274), .Y(n4451) );
  OAI211X1 U2062 ( .A0(n408), .A1(n925), .B0(n419), .C0(n3279), .Y(n4459) );
  NAND2X1 U2063 ( .A(H1[16]), .B(n205), .Y(n3279) );
  OAI211X1 U2064 ( .A0(n412), .A1(n1086), .B0(n3504), .C0(n419), .Y(n4703) );
  NAND2X1 U2065 ( .A(H0[30]), .B(n205), .Y(n3504) );
  OAI211X1 U2066 ( .A0(n412), .A1(n1090), .B0(n3505), .C0(n419), .Y(n4704) );
  NAND2X1 U2067 ( .A(H0[29]), .B(n205), .Y(n3505) );
  OAI211X1 U2068 ( .A0(n407), .A1(n1098), .B0(n3506), .C0(n419), .Y(n4706) );
  NAND2X1 U2069 ( .A(H0[27]), .B(n205), .Y(n3506) );
  OAI211X1 U2070 ( .A0(n410), .A1(n1231), .B0(n419), .C0(n3508), .Y(n4714) );
  NAND2X1 U2071 ( .A(H0[19]), .B(n205), .Y(n3508) );
  OAI211X1 U2072 ( .A0(n409), .A1(n1228), .B0(n419), .C0(n3509), .Y(n4717) );
  NAND2X1 U2073 ( .A(H0[16]), .B(n205), .Y(n3509) );
  OAI211X1 U2074 ( .A0(n407), .A1(n1227), .B0(n419), .C0(n3510), .Y(n4718) );
  NAND2X1 U2075 ( .A(H0[15]), .B(n205), .Y(n3510) );
  OAI211X1 U2076 ( .A0(n411), .A1(n1226), .B0(n419), .C0(n3511), .Y(n4719) );
  NAND2X1 U2077 ( .A(H0[14]), .B(n205), .Y(n3511) );
  OAI211X1 U2078 ( .A0(n1244), .A1(n1225), .B0(n419), .C0(n3512), .Y(n4720) );
  NAND2X1 U2079 ( .A(H0[13]), .B(n205), .Y(n3512) );
  OAI211X1 U2080 ( .A0(n407), .A1(n1170), .B0(n3515), .C0(n419), .Y(n4727) );
  NAND2X1 U2081 ( .A(H0[6]), .B(n205), .Y(n3515) );
  OAI211X1 U2082 ( .A0(n410), .A1(n1175), .B0(n3516), .C0(n419), .Y(n4728) );
  NAND2X1 U2083 ( .A(H0[5]), .B(n205), .Y(n3516) );
  XOR3X2 U2084 ( .A(n219), .B(n306), .C(n297), .Y(f3_A_32[5]) );
  XOR3X2 U2085 ( .A(SHA256_result[228]), .B(n309), .C(n300), .Y(f3_A_32[2]) );
  XOR3X2 U2086 ( .A(n150), .B(n291), .C(n90), .Y(f4_E_32[12]) );
  NAND2XL U2087 ( .A(next_E[14]), .B(n337), .Y(n749) );
  NAND4X1 U2088 ( .A(n756), .B(n755), .C(n802), .D(n754), .Y(n4558) );
  NAND2XL U2089 ( .A(n146), .B(n345), .Y(n754) );
  NAND2XL U2090 ( .A(next_E[12]), .B(n339), .Y(n756) );
  NAND2X1 U2091 ( .A(N949), .B(n807), .Y(n755) );
  OAI21XL U2092 ( .A0(n420), .A1(n137), .B0(n757), .Y(n4527) );
  NAND2X1 U2093 ( .A(H4[11]), .B(n205), .Y(n757) );
  NAND2X1 U2094 ( .A(H4[10]), .B(n205), .Y(n760) );
  NAND2X1 U2095 ( .A(H4[8]), .B(n205), .Y(n767) );
  OAI2BB1X2 U2096 ( .A0N(SHA256_result[207]), .A1N(n309), .B0(n1068), .Y(
        f2_ABC_32[15]) );
  OAI21X1 U2097 ( .A0(SHA256_result[207]), .A1(n309), .B0(SHA256_result[175]), 
        .Y(n1068) );
  XOR3X2 U2098 ( .A(n147), .B(n105), .C(SHA256_result[113]), .Y(f4_E_32[6]) );
  XOR3X2 U2099 ( .A(n171), .B(n106), .C(n118), .Y(f4_E_32[20]) );
  XOR3X2 U2100 ( .A(n146), .B(n244), .C(n115), .Y(f4_E_32[19]) );
  MX2X1 U2101 ( .A(SHA256_result[58]), .B(SHA256_result[90]), .S0(n117), .Y(
        f1_EFG_32[26]) );
  XOR3X2 U2102 ( .A(n222), .B(n310), .C(n301), .Y(f3_A_32[1]) );
  XOR3X2 U2103 ( .A(n18), .B(n305), .C(n296), .Y(f3_A_32[6]) );
  OAI2BB2X1 U2104 ( .B0(n420), .B1(n1320), .A0N(H1[19]), .A1N(n205), .Y(n4456)
         );
  OAI2BB2X1 U2105 ( .B0(n420), .B1(n1403), .A0N(H6[31]), .A1N(n205), .Y(n4348)
         );
  OAI2BB2X1 U2106 ( .B0(n420), .B1(n1370), .A0N(H4[21]), .A1N(n205), .Y(n4517)
         );
  OAI2BB2X1 U2107 ( .B0(n420), .B1(n1369), .A0N(H4[20]), .A1N(n205), .Y(n4518)
         );
  OAI2BB2X1 U2108 ( .B0(n420), .B1(n1321), .A0N(H1[20]), .A1N(n205), .Y(n4455)
         );
  OAI2BB2X1 U2109 ( .B0(n420), .B1(n1324), .A0N(H1[23]), .A1N(n205), .Y(n4452)
         );
  OAI2BB2X1 U2110 ( .B0(n420), .B1(n1234), .A0N(H1[26]), .A1N(n205), .Y(n4449)
         );
  OAI2BB2X1 U2111 ( .B0(n420), .B1(n1340), .A0N(H2[24]), .A1N(n205), .Y(n4482)
         );
  OAI2BB2X1 U2112 ( .B0(n420), .B1(n1332), .A0N(H2[16]), .A1N(n205), .Y(n4490)
         );
  OAI2BB2X1 U2113 ( .B0(n420), .B1(n1238), .A0N(H1[30]), .A1N(n205), .Y(n4445)
         );
  OAI2BB2X1 U2114 ( .B0(n420), .B1(n87), .A0N(H2[25]), .A1N(n205), .Y(n4481)
         );
  OAI2BB2X1 U2115 ( .B0(n420), .B1(n1345), .A0N(H2[30]), .A1N(n205), .Y(n4476)
         );
  OAI2BB2X1 U2116 ( .B0(n420), .B1(n1339), .A0N(H2[23]), .A1N(n205), .Y(n4483)
         );
  OAI2BB2X1 U2117 ( .B0(n420), .B1(n1336), .A0N(H2[20]), .A1N(n205), .Y(n4486)
         );
  OAI2BB2X1 U2118 ( .B0(n420), .B1(n1328), .A0N(H2[31]), .A1N(n205), .Y(n4475)
         );
  OAI2BB2X1 U2119 ( .B0(n420), .B1(n1392), .A0N(H6[19]), .A1N(n205), .Y(n4360)
         );
  OAI2BB2X1 U2120 ( .B0(n420), .B1(n1391), .A0N(H6[18]), .A1N(n205), .Y(n4361)
         );
  OAI2BB2X1 U2121 ( .B0(n420), .B1(n1393), .A0N(H6[20]), .A1N(n205), .Y(n4359)
         );
  OAI2BB2X1 U2122 ( .B0(n420), .B1(n1401), .A0N(H6[29]), .A1N(n205), .Y(n4350)
         );
  OAI2BB2X1 U2123 ( .B0(n420), .B1(n1375), .A0N(H5[19]), .A1N(n205), .Y(n4328)
         );
  OAI2BB2X1 U2124 ( .B0(n420), .B1(n1386), .A0N(H5[30]), .A1N(n205), .Y(n4317)
         );
  OAI2BB2X1 U2125 ( .B0(n420), .B1(n1378), .A0N(H5[22]), .A1N(n205), .Y(n4325)
         );
  OAI2BB2X1 U2126 ( .B0(n420), .B1(n1377), .A0N(H5[21]), .A1N(n205), .Y(n4326)
         );
  OAI2BB2X1 U2127 ( .B0(n420), .B1(n1376), .A0N(H5[20]), .A1N(n205), .Y(n4327)
         );
  OAI2BB2X1 U2128 ( .B0(n420), .B1(n1385), .A0N(H5[29]), .A1N(n205), .Y(n4318)
         );
  OAI21XL U2129 ( .A0(n420), .A1(n967), .B0(n966), .Y(n4504) );
  OAI21XL U2130 ( .A0(n420), .A1(n973), .B0(n972), .Y(n4506) );
  OAI21XL U2131 ( .A0(n420), .A1(n217), .B0(n1167), .Y(n4726) );
  NAND2X1 U2132 ( .A(H0[7]), .B(n205), .Y(n1167) );
  OAI211XL U2133 ( .A0(n334), .A1(n1210), .B0(n515), .C0(n514), .Y(n4310) );
  OAI211XL U2134 ( .A0(n335), .A1(n685), .B0(n575), .C0(n574), .Y(n4399) );
  NAND2X1 U2135 ( .A(N885), .B(n807), .Y(n575) );
  NAND2X1 U2136 ( .A(N878), .B(n807), .Y(n592) );
  AOI21XL U2137 ( .A0(n174), .A1(n342), .B0(n327), .Y(n591) );
  OAI21XL U2138 ( .A0(n420), .A1(n170), .B0(n750), .Y(n4525) );
  NAND2X1 U2139 ( .A(H4[13]), .B(n205), .Y(n750) );
  NAND2X1 U2140 ( .A(H0[3]), .B(n205), .Y(n1184) );
  OAI2BB2X1 U2141 ( .B0(n420), .B1(n1428), .A0N(H7[31]), .A1N(n205), .Y(n4252)
         );
  INVX1 U2142 ( .A(SHA256_result[31]), .Y(n1428) );
  OAI2BB2X1 U2143 ( .B0(n420), .B1(n1426), .A0N(H7[29]), .A1N(n205), .Y(n4254)
         );
  INVX1 U2144 ( .A(SHA256_result[29]), .Y(n1426) );
  OAI2BB2X1 U2145 ( .B0(n420), .B1(n1423), .A0N(H7[26]), .A1N(n205), .Y(n4257)
         );
  INVX1 U2146 ( .A(SHA256_result[26]), .Y(n1423) );
  OAI2BB2X1 U2147 ( .B0(n420), .B1(n1417), .A0N(H7[20]), .A1N(n205), .Y(n4263)
         );
  INVX1 U2148 ( .A(SHA256_result[20]), .Y(n1417) );
  OAI2BB2X1 U2149 ( .B0(n420), .B1(n1416), .A0N(H7[19]), .A1N(n205), .Y(n4264)
         );
  INVX1 U2150 ( .A(SHA256_result[19]), .Y(n1416) );
  INVX1 U2151 ( .A(SHA256_result[18]), .Y(n1415) );
  INVX1 U2152 ( .A(SHA256_result[17]), .Y(n1414) );
  INVX1 U2153 ( .A(SHA256_result[16]), .Y(n1413) );
  INVX1 U2154 ( .A(SHA256_result[13]), .Y(n1410) );
  INVX1 U2155 ( .A(SHA256_result[12]), .Y(n1409) );
  OAI2BB2X1 U2156 ( .B0(n420), .B1(n1402), .A0N(H6[30]), .A1N(n205), .Y(n4349)
         );
  INVX1 U2157 ( .A(SHA256_result[62]), .Y(n1402) );
  OAI2BB2X1 U2158 ( .B0(n420), .B1(n1395), .A0N(H6[22]), .A1N(n205), .Y(n4357)
         );
  INVXL U2159 ( .A(SHA256_result[54]), .Y(n1395) );
  OAI2BB2X1 U2160 ( .B0(n420), .B1(n1394), .A0N(H6[21]), .A1N(n205), .Y(n4358)
         );
  INVXL U2161 ( .A(SHA256_result[53]), .Y(n1394) );
  OAI2BB2X1 U2162 ( .B0(n420), .B1(n1382), .A0N(H5[26]), .A1N(n205), .Y(n4321)
         );
  OAI2BB2X1 U2163 ( .B0(n420), .B1(n1379), .A0N(H5[23]), .A1N(n205), .Y(n4324)
         );
  INVXL U2164 ( .A(SHA256_result[87]), .Y(n1379) );
  OAI2BB2X1 U2165 ( .B0(n420), .B1(n1373), .A0N(H5[17]), .A1N(n205), .Y(n4330)
         );
  INVXL U2166 ( .A(SHA256_result[81]), .Y(n1373) );
  INVXL U2167 ( .A(SHA256_result[79]), .Y(n1371) );
  OAI21XL U2168 ( .A0(n420), .A1(n1164), .B0(n1163), .Y(n4725) );
  NAND2X1 U2169 ( .A(H0[8]), .B(n205), .Y(n1163) );
  INVX1 U2170 ( .A(SHA256_result[158]), .Y(n1366) );
  INVX1 U2171 ( .A(SHA256_result[156]), .Y(n1364) );
  INVX1 U2172 ( .A(SHA256_result[155]), .Y(n1363) );
  INVX1 U2173 ( .A(SHA256_result[153]), .Y(n1361) );
  INVX1 U2174 ( .A(SHA256_result[151]), .Y(n1359) );
  INVX1 U2175 ( .A(SHA256_result[149]), .Y(n1357) );
  INVX1 U2176 ( .A(SHA256_result[148]), .Y(n1356) );
  INVX1 U2177 ( .A(SHA256_result[139]), .Y(n1347) );
  OAI21XL U2178 ( .A0(n420), .A1(n1181), .B0(n1180), .Y(n4729) );
  NAND2X1 U2179 ( .A(H0[4]), .B(n205), .Y(n1180) );
  NAND2X1 U2180 ( .A(H4[31]), .B(n205), .Y(n804) );
  OAI21XL U2181 ( .A0(n420), .A1(n684), .B0(n571), .Y(n4366) );
  OAI21XL U2182 ( .A0(n420), .A1(n685), .B0(n645), .Y(n4335) );
  OAI21XL U2183 ( .A0(n420), .A1(n739), .B0(n738), .Y(n4522) );
  NAND2X1 U2184 ( .A(H4[16]), .B(n205), .Y(n738) );
  OAI21XL U2185 ( .A0(n420), .A1(n722), .B0(n721), .Y(n4516) );
  NAND2X1 U2186 ( .A(H4[22]), .B(n205), .Y(n721) );
  OAI21XL U2187 ( .A0(n420), .A1(n116), .B0(n711), .Y(n4512) );
  NAND2X1 U2188 ( .A(H4[26]), .B(n205), .Y(n711) );
  OAI21XL U2189 ( .A0(n420), .A1(n243), .B0(n713), .Y(n4513) );
  NAND2X1 U2190 ( .A(H4[25]), .B(n205), .Y(n713) );
  OAI21XL U2191 ( .A0(n420), .A1(n121), .B0(n709), .Y(n4511) );
  NAND2X1 U2192 ( .A(H4[27]), .B(n205), .Y(n709) );
  OAI21XL U2193 ( .A0(n420), .A1(n91), .B0(n719), .Y(n4515) );
  NAND2X1 U2194 ( .A(H4[23]), .B(n205), .Y(n719) );
  OAI21XL U2195 ( .A0(n420), .A1(n128), .B0(n664), .Y(n4342) );
  OAI21XL U2196 ( .A0(n420), .A1(n1216), .B0(n521), .Y(n4282) );
  OAI21XL U2197 ( .A0(n420), .A1(n1207), .B0(n508), .Y(n4277) );
  OAI21XL U2198 ( .A0(n420), .A1(n1209), .B0(n511), .Y(n4278) );
  OAI21XL U2199 ( .A0(n420), .A1(n1151), .B0(n1150), .Y(n4722) );
  NAND2X1 U2200 ( .A(H0[11]), .B(n205), .Y(n1150) );
  OAI21XL U2201 ( .A0(n420), .A1(n1119), .B0(n1118), .Y(n4711) );
  NAND2X1 U2202 ( .A(H0[22]), .B(n205), .Y(n1118) );
  OAI21XL U2203 ( .A0(n420), .A1(n1111), .B0(n1110), .Y(n4709) );
  NAND2X1 U2204 ( .A(H0[24]), .B(n205), .Y(n1110) );
  OAI21XL U2205 ( .A0(n420), .A1(n1051), .B0(n1050), .Y(n4702) );
  NAND2X1 U2206 ( .A(H0[31]), .B(n205), .Y(n1050) );
  NAND2X1 U2207 ( .A(H4[7]), .B(n205), .Y(n771) );
  OAI21XL U2208 ( .A0(n420), .A1(n743), .B0(n742), .Y(n4523) );
  NAND2X1 U2209 ( .A(H4[15]), .B(n205), .Y(n742) );
  OAI21XL U2210 ( .A0(n420), .A1(n1146), .B0(n1145), .Y(n4721) );
  NAND2X1 U2211 ( .A(H0[12]), .B(n205), .Y(n1145) );
  OAI21XL U2212 ( .A0(n420), .A1(n1095), .B0(n1094), .Y(n4705) );
  NAND2X1 U2213 ( .A(H0[28]), .B(n205), .Y(n1094) );
  OAI21XL U2214 ( .A0(n420), .A1(n1103), .B0(n1102), .Y(n4707) );
  NAND2X1 U2215 ( .A(H0[26]), .B(n205), .Y(n1102) );
  OAI21XL U2216 ( .A0(n420), .A1(n1115), .B0(n1114), .Y(n4710) );
  NAND2X1 U2217 ( .A(H0[23]), .B(n205), .Y(n1114) );
  OAI21XL U2218 ( .A0(n420), .A1(n160), .B0(n578), .Y(n4369) );
  OAI21XL U2219 ( .A0(n420), .A1(n166), .B0(n581), .Y(n4370) );
  OAI21XL U2220 ( .A0(n420), .A1(n1206), .B0(n588), .Y(n4373) );
  OAI21XL U2221 ( .A0(n420), .A1(n1210), .B0(n593), .Y(n4375) );
  OAI21XL U2222 ( .A0(n420), .A1(n689), .B0(n650), .Y(n4337) );
  OAI21XL U2223 ( .A0(n420), .A1(n690), .B0(n653), .Y(n4338) );
  OAI21XL U2224 ( .A0(n420), .A1(n691), .B0(n656), .Y(n4339) );
  OAI21XL U2225 ( .A0(n420), .A1(n699), .B0(n678), .Y(n4347) );
  OAI21XL U2226 ( .A0(n420), .A1(n1215), .B0(n518), .Y(n4281) );
  OAI211XL U2227 ( .A0(n332), .A1(n1217), .B0(n525), .C0(n524), .Y(n4314) );
  NAND3BX1 U2228 ( .AN(n992), .B(n379), .C(n991), .Y(n4673) );
  NAND3BX1 U2230 ( .AN(n1023), .B(n376), .C(n1022), .Y(n4687) );
  NAND2XL U2231 ( .A(SHA256_result[203]), .B(n399), .Y(n1022) );
  NAND2X1 U2232 ( .A(N1044), .B(n356), .Y(n1021) );
  NAND3BX1 U2233 ( .AN(n1026), .B(n377), .C(n1025), .Y(n4688) );
  NAND2XL U2234 ( .A(SHA256_result[202]), .B(n399), .Y(n1025) );
  NAND2X1 U2235 ( .A(N1043), .B(n356), .Y(n1024) );
  NAND3BX1 U2236 ( .AN(n1045), .B(n378), .C(n1044), .Y(n4696) );
  NAND2XL U2237 ( .A(SHA256_result[194]), .B(n399), .Y(n1044) );
  OAI21XL U2238 ( .A0(n21), .A1(n1188), .B0(n1043), .Y(n1045) );
  NAND3BX1 U2239 ( .AN(n1034), .B(n377), .C(n1033), .Y(n4691) );
  NAND2XL U2240 ( .A(SHA256_result[199]), .B(n399), .Y(n1033) );
  NAND3BX1 U2241 ( .AN(n979), .B(n375), .C(n978), .Y(n4667) );
  NAND2X1 U2242 ( .A(N1064), .B(n355), .Y(n977) );
  NAND3BX1 U2243 ( .AN(n858), .B(n382), .C(n857), .Y(n4624) );
  OAI21XL U2244 ( .A0(n28), .A1(n941), .B0(n856), .Y(n858) );
  NAND3BX1 U2245 ( .AN(n875), .B(n375), .C(n874), .Y(n4629) );
  NAND3BX1 U2246 ( .AN(n1029), .B(n377), .C(n1028), .Y(n4689) );
  NAND2XL U2247 ( .A(SHA256_result[201]), .B(n399), .Y(n1028) );
  NAND2X1 U2248 ( .A(N1042), .B(n356), .Y(n1027) );
  NAND3X1 U2249 ( .A(n537), .B(n536), .C(n535), .Y(n4384) );
  NAND3X1 U2250 ( .A(n543), .B(n542), .C(n541), .Y(n4386) );
  NAND3X1 U2251 ( .A(n546), .B(n545), .C(n544), .Y(n4387) );
  NAND3X1 U2252 ( .A(n534), .B(n533), .C(n532), .Y(n4383) );
  NAND3X1 U2253 ( .A(n549), .B(n548), .C(n547), .Y(n4388) );
  NAND2XL U2254 ( .A(n337), .B(SHA256_result[87]), .Y(n549) );
  NAND3X1 U2255 ( .A(n568), .B(n567), .C(n566), .Y(n4396) );
  NAND2XL U2256 ( .A(n337), .B(SHA256_result[79]), .Y(n568) );
  AOI21XL U2257 ( .A0(n344), .A1(SHA256_result[47]), .B0(n327), .Y(n566) );
  NAND3X1 U2258 ( .A(n540), .B(n539), .C(n538), .Y(n4385) );
  NAND3X1 U2259 ( .A(n562), .B(n561), .C(n560), .Y(n4394) );
  NAND2XL U2260 ( .A(n338), .B(SHA256_result[81]), .Y(n562) );
  AOI21XL U2261 ( .A0(n344), .A1(SHA256_result[49]), .B0(n326), .Y(n560) );
  NAND3X1 U2262 ( .A(n565), .B(n564), .C(n563), .Y(n4395) );
  NAND2XL U2263 ( .A(n339), .B(SHA256_result[80]), .Y(n565) );
  AOI21XL U2264 ( .A0(n344), .A1(SHA256_result[48]), .B0(n326), .Y(n563) );
  NAND3X1 U2265 ( .A(n453), .B(n452), .C(n451), .Y(n4284) );
  NAND2X1 U2266 ( .A(n336), .B(SHA256_result[62]), .Y(n453) );
  NAND3X1 U2267 ( .A(n458), .B(n457), .C(n456), .Y(n4286) );
  NAND2X1 U2268 ( .A(n336), .B(SHA256_result[60]), .Y(n458) );
  NAND2X1 U2269 ( .A(N869), .B(n807), .Y(n457) );
  NAND3X1 U2270 ( .A(n461), .B(n460), .C(n459), .Y(n4287) );
  NAND2X1 U2271 ( .A(N868), .B(n807), .Y(n460) );
  NAND2X1 U2272 ( .A(n336), .B(SHA256_result[59]), .Y(n461) );
  NAND3X1 U2273 ( .A(n466), .B(n465), .C(n464), .Y(n4289) );
  NAND2X1 U2274 ( .A(N866), .B(n807), .Y(n465) );
  NAND3X1 U2275 ( .A(n469), .B(n468), .C(n467), .Y(n4290) );
  NAND2X1 U2276 ( .A(N865), .B(n807), .Y(n468) );
  NAND3X1 U2277 ( .A(n472), .B(n471), .C(n470), .Y(n4291) );
  NAND2X1 U2278 ( .A(N864), .B(n807), .Y(n471) );
  NAND2XL U2279 ( .A(n340), .B(SHA256_result[55]), .Y(n472) );
  NAND3X1 U2280 ( .A(n475), .B(n474), .C(n473), .Y(n4292) );
  NAND2X1 U2281 ( .A(N863), .B(n807), .Y(n474) );
  NAND2XL U2282 ( .A(n336), .B(SHA256_result[54]), .Y(n475) );
  NAND3X1 U2283 ( .A(n478), .B(n477), .C(n476), .Y(n4293) );
  NAND2X1 U2284 ( .A(N862), .B(n807), .Y(n477) );
  NAND2XL U2285 ( .A(n338), .B(SHA256_result[53]), .Y(n478) );
  NAND3X1 U2286 ( .A(n491), .B(n490), .C(n489), .Y(n4299) );
  NAND2X1 U2287 ( .A(N856), .B(n807), .Y(n490) );
  NAND2XL U2288 ( .A(n340), .B(SHA256_result[47]), .Y(n491) );
  NAND3X1 U2289 ( .A(n607), .B(n606), .C(n605), .Y(n4412) );
  NAND2XL U2290 ( .A(n339), .B(n106), .Y(n607) );
  NAND3X1 U2291 ( .A(n634), .B(n633), .C(n632), .Y(n4425) );
  NAND2X1 U2292 ( .A(N923), .B(n807), .Y(n633) );
  AOI21XL U2293 ( .A0(n343), .A1(SHA256_result[82]), .B0(n328), .Y(n632) );
  BUFX12 U2294 ( .A(SHA256_result[239]), .Y(n309) );
  BUFX12 U2295 ( .A(SHA256_result[234]), .Y(n311) );
  BUFX12 U2296 ( .A(SHA256_result[233]), .Y(n312) );
  BUFX12 U2297 ( .A(SHA256_result[226]), .Y(n315) );
  BUFX12 U2298 ( .A(SHA256_result[230]), .Y(n313) );
  BUFX12 U2299 ( .A(SHA256_result[229]), .Y(n314) );
  MX2X1 U2300 ( .A(SHA256_result[31]), .B(SHA256_result[63]), .S0(
        mux_control_0_), .Y(mux2[31]) );
  NAND2BXL U2301 ( .AN(n334), .B(next_E[16]), .Y(n740) );
  NAND2BXL U2302 ( .AN(n333), .B(next_E[20]), .Y(n727) );
  OAI211XL U2303 ( .A0(n408), .A1(n1217), .B0(n3204), .C0(n419), .Y(n4379) );
  NAND4X1 U2304 ( .A(n1262), .B(n2946), .C(n2925), .D(n2878), .Y(n3578) );
  NAND3X1 U2305 ( .A(n427), .B(n2906), .C(n4042), .Y(n4107) );
  INVXL U2306 ( .A(SHA256_result[203]), .Y(n939) );
  INVX1 U2307 ( .A(N1012), .Y(n938) );
  OAI222XL U2308 ( .A0(n26), .A1(n943), .B0(n365), .B1(n942), .C0(n351), .C1(
        n941), .Y(n4656) );
  INVXL U2309 ( .A(SHA256_result[202]), .Y(n943) );
  INVX1 U2310 ( .A(N1011), .Y(n942) );
  OAI222XL U2311 ( .A0(n23), .A1(n953), .B0(n366), .B1(n952), .C0(n350), .C1(
        n951), .Y(n4659) );
  INVXL U2312 ( .A(SHA256_result[199]), .Y(n953) );
  INVX1 U2313 ( .A(N1008), .Y(n952) );
  OAI222XL U2314 ( .A0(n26), .A1(n98), .B0(n366), .B1(n965), .C0(n349), .C1(
        n964), .Y(n4663) );
  INVX1 U2315 ( .A(N1004), .Y(n965) );
  OAI222XL U2316 ( .A0(n23), .A1(n1308), .B0(n367), .B1(n968), .C0(n352), .C1(
        n967), .Y(n4664) );
  INVX1 U2317 ( .A(N1003), .Y(n968) );
  OAI222XL U2318 ( .A0(n25), .A1(n97), .B0(n365), .B1(n974), .C0(n204), .C1(
        n973), .Y(n4666) );
  INVX1 U2319 ( .A(N1001), .Y(n974) );
  OAI221XL U2320 ( .A0(n366), .A1(n854), .B0(n27), .B1(n937), .C0(n853), .Y(
        n4623) );
  INVX1 U2321 ( .A(N980), .Y(n854) );
  OAI221XL U2322 ( .A0(n364), .A1(n826), .B0(n87), .B1(n25), .C0(n825), .Y(
        n4609) );
  INVX1 U2323 ( .A(N994), .Y(n826) );
  NAND2X1 U2324 ( .A(n247), .B(SHA256_result[153]), .Y(n825) );
  OAI221XL U2325 ( .A0(n364), .A1(n897), .B0(n1238), .B1(n22), .C0(n896), .Y(
        n4636) );
  INVX1 U2326 ( .A(N1031), .Y(n897) );
  NAND2X1 U2327 ( .A(n247), .B(SHA256_result[190]), .Y(n896) );
  OAI221XL U2328 ( .A0(n360), .A1(n814), .B0(n1345), .B1(n26), .C0(n813), .Y(
        n4604) );
  INVX1 U2329 ( .A(N999), .Y(n814) );
  NAND2X1 U2330 ( .A(n247), .B(SHA256_result[158]), .Y(n813) );
  OAI221XL U2331 ( .A0(n365), .A1(n830), .B0(n1339), .B1(n21), .C0(n829), .Y(
        n4611) );
  INVX1 U2332 ( .A(N992), .Y(n830) );
  NAND2X1 U2333 ( .A(n247), .B(SHA256_result[151]), .Y(n829) );
  OAI221XL U2334 ( .A0(n365), .A1(n836), .B0(n1336), .B1(n22), .C0(n835), .Y(
        n4614) );
  INVX1 U2335 ( .A(N989), .Y(n836) );
  NAND2X1 U2336 ( .A(n247), .B(SHA256_result[148]), .Y(n835) );
  OAI221XL U2337 ( .A0(n366), .A1(n822), .B0(n1342), .B1(n26), .C0(n821), .Y(
        n4607) );
  INVX1 U2338 ( .A(N996), .Y(n822) );
  NAND2X1 U2339 ( .A(n247), .B(SHA256_result[155]), .Y(n821) );
  OAI221XL U2340 ( .A0(n362), .A1(n820), .B0(n1343), .B1(n23), .C0(n819), .Y(
        n4606) );
  INVX1 U2341 ( .A(N997), .Y(n820) );
  NAND2X1 U2342 ( .A(n247), .B(SHA256_result[156]), .Y(n819) );
  OAI221XL U2343 ( .A0(n366), .A1(n834), .B0(n1337), .B1(n21), .C0(n833), .Y(
        n4613) );
  INVX1 U2344 ( .A(N990), .Y(n834) );
  NAND2X1 U2345 ( .A(n247), .B(SHA256_result[149]), .Y(n833) );
  OAI221XL U2346 ( .A0(n363), .A1(n989), .B0(n22), .B1(n1103), .C0(n988), .Y(
        n4672) );
  INVX1 U2347 ( .A(N1059), .Y(n989) );
  OAI221XL U2348 ( .A0(n365), .A1(n907), .B0(n28), .B1(n1326), .C0(n906), .Y(
        n4641) );
  INVX1 U2349 ( .A(N1026), .Y(n907) );
  OAI221XL U2350 ( .A0(n364), .A1(n909), .B0(n23), .B1(n1325), .C0(n908), .Y(
        n4642) );
  INVX1 U2351 ( .A(N1025), .Y(n909) );
  OAI221XL U2352 ( .A0(n363), .A1(n911), .B0(n25), .B1(n1324), .C0(n910), .Y(
        n4643) );
  INVX1 U2353 ( .A(N1024), .Y(n911) );
  OAI221XL U2354 ( .A0(n363), .A1(n917), .B0(n27), .B1(n1321), .C0(n916), .Y(
        n4646) );
  INVX1 U2355 ( .A(N1021), .Y(n917) );
  OAI221XL U2356 ( .A0(n363), .A1(n926), .B0(n28), .B1(n925), .C0(n924), .Y(
        n4650) );
  INVX1 U2357 ( .A(N1017), .Y(n926) );
  OAI221XL U2358 ( .A0(n363), .A1(n976), .B0(n28), .B1(n1327), .C0(n975), .Y(
        n4635) );
  INVX1 U2359 ( .A(N1032), .Y(n976) );
  NAND2X1 U2360 ( .A(n247), .B(SHA256_result[191]), .Y(n975) );
  OAI221XL U2361 ( .A0(n363), .A1(n981), .B0(n27), .B1(n1086), .C0(n980), .Y(
        n4668) );
  INVX1 U2362 ( .A(N1063), .Y(n981) );
  NAND2X1 U2363 ( .A(n247), .B(SHA256_result[222]), .Y(n980) );
  INVXL U2364 ( .A(SHA256_result[170]), .Y(n941) );
  INVXL U2365 ( .A(SHA256_result[163]), .Y(n964) );
  INVXL U2366 ( .A(SHA256_result[162]), .Y(n967) );
  INVXL U2367 ( .A(SHA256_result[160]), .Y(n973) );
  INVXL U2368 ( .A(SHA256_result[167]), .Y(n951) );
  MX2XL U2369 ( .A(SHA256_result[141]), .B(SHA256_result[173]), .S0(n438), .Y(
        mux1[13]) );
  INVXL U2370 ( .A(SHA256_result[168]), .Y(n947) );
  INVXL U2371 ( .A(SHA256_result[164]), .Y(n960) );
  INVXL U2372 ( .A(SHA256_result[165]), .Y(n957) );
  INVXL U2373 ( .A(SHA256_result[169]), .Y(n944) );
  INVXL U2374 ( .A(SHA256_result[166]), .Y(n954) );
  INVX1 U2375 ( .A(SHA256_result[137]), .Y(n860) );
  INVX1 U2376 ( .A(SHA256_result[134]), .Y(n870) );
  INVX1 U2377 ( .A(SHA256_result[135]), .Y(n867) );
  OAI2BB1X1 U2378 ( .A0N(SHA256_result[216]), .A1N(n300), .B0(n1059), .Y(
        f2_ABC_32[24]) );
  OAI2BB1X1 U2379 ( .A0N(SHA256_result[217]), .A1N(n299), .B0(n1058), .Y(
        f2_ABC_32[25]) );
  OAI2BB1X1 U2380 ( .A0N(n298), .A1N(SHA256_result[218]), .B0(n1057), .Y(
        f2_ABC_32[26]) );
  OAI21XL U2381 ( .A0(n298), .A1(SHA256_result[218]), .B0(SHA256_result[186]), 
        .Y(n1057) );
  XOR3X2 U2382 ( .A(n292), .B(n106), .C(n291), .Y(f4_E_32[25]) );
  OAI222XL U2383 ( .A0(round[6]), .A1(n4248), .B0(n4249), .B1(n1285), .C0(n809), .C1(n808), .Y(n4247) );
  INVX1 U2384 ( .A(n4248), .Y(n1285) );
  MX2X1 U2385 ( .A(SHA256_result[59]), .B(SHA256_result[91]), .S0(n123), .Y(
        f1_EFG_32[27]) );
  MX2X1 U2386 ( .A(SHA256_result[60]), .B(SHA256_result[92]), .S0(n94), .Y(
        f1_EFG_32[28]) );
  XOR3X2 U2387 ( .A(n219), .B(n305), .C(n294), .Y(f3_A_32[17]) );
  XOR3X2 U2388 ( .A(n222), .B(SHA256_result[236]), .C(n300), .Y(f3_A_32[22])
         );
  XOR3X2 U2389 ( .A(n18), .B(n304), .C(n293), .Y(f3_A_32[18]) );
  XOR3X2 U2390 ( .A(n88), .B(n308), .C(n297), .Y(f3_A_32[14]) );
  MX2XL U2391 ( .A(SHA256_result[143]), .B(SHA256_result[175]), .S0(n438), .Y(
        mux1[15]) );
  CLKINVX3 U2392 ( .A(n439), .Y(n438) );
  INVX1 U2393 ( .A(SHA256_result[129]), .Y(n887) );
  INVX1 U2394 ( .A(SHA256_result[138]), .Y(n855) );
  INVX1 U2395 ( .A(SHA256_result[136]), .Y(n862) );
  INVX1 U2396 ( .A(SHA256_result[131]), .Y(n880) );
  INVX1 U2397 ( .A(SHA256_result[132]), .Y(n876) );
  INVX1 U2398 ( .A(SHA256_result[133]), .Y(n872) );
  MX2XL U2399 ( .A(SHA256_result[142]), .B(SHA256_result[174]), .S0(n438), .Y(
        mux1[14]) );
  OAI2BB1X1 U2400 ( .A0N(SHA256_result[223]), .A1N(n293), .B0(n1052), .Y(
        f2_ABC_32[31]) );
  OAI21XL U2401 ( .A0(n293), .A1(SHA256_result[223]), .B0(SHA256_result[191]), 
        .Y(n1052) );
  OAI222XL U2402 ( .A0(n4156), .A1(n2938), .B0(n429), .B1(n4157), .C0(n432), 
        .C1(n1247), .Y(n4155) );
  INVX1 U2403 ( .A(n4009), .Y(n1247) );
  AOI31X1 U2404 ( .A0(n3951), .A1(n3952), .A2(n3953), .B0(n418), .Y(N3163) );
  AOI31X1 U2405 ( .A0(n4234), .A1(n4235), .A2(n4236), .B0(n417), .Y(N3134) );
  AOI31X1 U2406 ( .A0(n4220), .A1(n4221), .A2(n4222), .B0(n417), .Y(N3136) );
  AOI31X1 U2407 ( .A0(n4109), .A1(n4110), .A2(n4111), .B0(n418), .Y(N3151) );
  AOI211X1 U2408 ( .A0(n4113), .A1(n425), .B0(n3947), .C0(n4025), .Y(n4110) );
  AOI31X1 U2409 ( .A0(n4186), .A1(n4187), .A2(n4188), .B0(n417), .Y(N3141) );
  AOI31X1 U2410 ( .A0(n4228), .A1(n4229), .A2(n4230), .B0(n417), .Y(N3135) );
  AOI222XL U2411 ( .A0(n259), .A1(n4042), .B0(n4233), .B1(n2925), .C0(n4227), 
        .C1(n422), .Y(n4229) );
  AOI31X1 U2412 ( .A0(n4208), .A1(n4209), .A2(n4210), .B0(n417), .Y(N3138) );
  AOI211XL U2413 ( .A0(n259), .A1(n4211), .B0(n4212), .C0(n4213), .Y(n4210) );
  AOI31X1 U2414 ( .A0(n4076), .A1(n4077), .A2(n4078), .B0(n418), .Y(N3154) );
  AOI222XL U2415 ( .A0(n1269), .A1(n427), .B0(n4088), .B1(n432), .C0(n260), 
        .C1(n3946), .Y(n4076) );
  AOI221X1 U2416 ( .A0(n3954), .A1(n4083), .B0(n4084), .B1(n2906), .C0(n4085), 
        .Y(n4077) );
  NOR4BX1 U2417 ( .AN(n1296), .B(n4079), .C(n4080), .D(n4081), .Y(n4078) );
  AOI31X1 U2418 ( .A0(n4089), .A1(n4090), .A2(n4091), .B0(n418), .Y(N3153) );
  AOI211X1 U2419 ( .A0(n434), .A1(n4095), .B0(n4096), .C0(n1249), .Y(n4090) );
  NOR3X1 U2420 ( .A(n4092), .B(n1269), .C(n4075), .Y(n4091) );
  AOI31X1 U2421 ( .A0(n4141), .A1(n4142), .A2(n4143), .B0(n417), .Y(N3147) );
  AOI222XL U2422 ( .A0(n429), .A1(n4148), .B0(n4149), .B1(n4105), .C0(n4150), 
        .C1(n259), .Y(n4142) );
  NOR3X1 U2423 ( .A(n4144), .B(n4145), .C(n4146), .Y(n4143) );
  AOI31X1 U2424 ( .A0(n3939), .A1(n3940), .A2(n3941), .B0(n417), .Y(N3164) );
  NOR2X1 U2425 ( .A(n3949), .B(n3950), .Y(n3939) );
  OAI2BB1X1 U2426 ( .A0N(n297), .A1N(SHA256_result[219]), .B0(n1056), .Y(
        f2_ABC_32[27]) );
  OAI21XL U2427 ( .A0(n297), .A1(SHA256_result[219]), .B0(SHA256_result[187]), 
        .Y(n1056) );
  OAI2BB1X1 U2428 ( .A0N(n296), .A1N(SHA256_result[220]), .B0(n1055), .Y(
        f2_ABC_32[28]) );
  OAI21XL U2429 ( .A0(n296), .A1(SHA256_result[220]), .B0(SHA256_result[188]), 
        .Y(n1055) );
  BUFX3 U2430 ( .A(round[1]), .Y(n320) );
  MX2X1 U2431 ( .A(SHA256_result[62]), .B(SHA256_result[94]), .S0(n115), .Y(
        f1_EFG_32[30]) );
  INVX1 U2432 ( .A(SHA256_result[1]), .Y(n1216) );
  INVX1 U2433 ( .A(SHA256_result[5]), .Y(n1209) );
  INVX1 U2434 ( .A(SHA256_result[6]), .Y(n1207) );
  XOR3X2 U2435 ( .A(n219), .B(n308), .C(n296), .Y(f3_A_32[26]) );
  XOR3X2 U2436 ( .A(n88), .B(SHA256_result[237]), .C(n299), .Y(f3_A_32[23]) );
  XOR3X2 U2437 ( .A(n18), .B(n307), .C(n295), .Y(f3_A_32[27]) );
  MX2XL U2438 ( .A(SHA256_result[15]), .B(SHA256_result[47]), .S0(
        mux_control_0_), .Y(mux2[15]) );
  MX2X1 U2439 ( .A(SHA256_result[155]), .B(SHA256_result[187]), .S0(n438), .Y(
        mux1[27]) );
  MX2X1 U2440 ( .A(SHA256_result[154]), .B(SHA256_result[186]), .S0(n438), .Y(
        mux1[26]) );
  MX2XL U2441 ( .A(SHA256_result[17]), .B(SHA256_result[49]), .S0(
        mux_control_0_), .Y(mux2[17]) );
  INVX1 U2442 ( .A(SHA256_result[4]), .Y(n1211) );
  INVX1 U2443 ( .A(SHA256_result[2]), .Y(n1215) );
  INVX1 U2444 ( .A(SHA256_result[0]), .Y(n1218) );
  NAND2X1 U2445 ( .A(n264), .B(n3678), .Y(N3584) );
  XNOR2X1 U2446 ( .A(read_counter[5]), .B(n1242), .Y(n264) );
  NAND2X1 U2447 ( .A(n265), .B(n3678), .Y(N3583) );
  XOR2X1 U2448 ( .A(read_counter[4]), .B(n1241), .Y(n265) );
  NAND2BX1 U2449 ( .AN(N3566), .B(n3678), .Y(N3582) );
  NAND2BX1 U2450 ( .AN(N3565), .B(n3678), .Y(N3581) );
  NAND2BX1 U2451 ( .AN(N3564), .B(n3678), .Y(N3580) );
  NAND2X1 U2452 ( .A(read_counter[0]), .B(n3678), .Y(N3579) );
  INVX1 U2453 ( .A(n433), .Y(n432) );
  INVX1 U2454 ( .A(round[2]), .Y(n433) );
  INVX1 U2455 ( .A(n2947), .Y(n423) );
  OAI222XL U2456 ( .A0(n4102), .A1(n2938), .B0(n1305), .B1(n1282), .C0(n4103), 
        .C1(n1298), .Y(n4101) );
  AOI21XL U2457 ( .A0(n259), .A1(n289), .B0(n3989), .Y(n4102) );
  OAI222XL U2458 ( .A0(n432), .A1(n4191), .B0(n2938), .B1(n3992), .C0(n3948), 
        .C1(n808), .Y(n4189) );
  NOR2X1 U2459 ( .A(n1257), .B(n2938), .Y(n3990) );
  OAI221XL U2460 ( .A0(n422), .A1(n1301), .B0(n2925), .B1(n1275), .C0(n1276), 
        .Y(n4239) );
  NOR2X1 U2461 ( .A(n3958), .B(n2938), .Y(n4159) );
  NOR2X1 U2462 ( .A(n2938), .B(n808), .Y(n3964) );
  NOR2X1 U2463 ( .A(n1251), .B(n2938), .Y(n4070) );
  OAI2BB1X1 U2464 ( .A0N(n427), .A1N(n4017), .B0(n4018), .Y(n3978) );
  AOI31XL U2465 ( .A0(n425), .A1(n2938), .A2(n259), .B0(n1268), .Y(n4018) );
  INVX1 U2466 ( .A(n4019), .Y(n1268) );
  OAI21XL U2467 ( .A0(n2906), .A1(n1274), .B0(n1260), .Y(n4120) );
  NOR2X1 U2468 ( .A(n289), .B(n2938), .Y(n4194) );
  OAI2BB1X1 U2469 ( .A0N(n295), .A1N(SHA256_result[221]), .B0(n1054), .Y(
        f2_ABC_32[29]) );
  OAI21XL U2470 ( .A0(n295), .A1(SHA256_result[221]), .B0(SHA256_result[189]), 
        .Y(n1054) );
  OAI2BB1X1 U2471 ( .A0N(n294), .A1N(SHA256_result[222]), .B0(n1053), .Y(
        f2_ABC_32[30]) );
  OAI21XL U2472 ( .A0(n294), .A1(SHA256_result[222]), .B0(SHA256_result[190]), 
        .Y(n1053) );
  MX2XL U2473 ( .A(SHA256_result[23]), .B(SHA256_result[55]), .S0(
        mux_control_0_), .Y(mux2[23]) );
  MX2XL U2474 ( .A(SHA256_result[21]), .B(SHA256_result[53]), .S0(
        mux_control_0_), .Y(mux2[21]) );
  MX2XL U2475 ( .A(SHA256_result[22]), .B(SHA256_result[54]), .S0(
        mux_control_0_), .Y(mux2[22]) );
  MX2X1 U2476 ( .A(SHA256_result[156]), .B(SHA256_result[188]), .S0(n438), .Y(
        mux1[28]) );
  MX2X1 U2477 ( .A(SHA256_result[157]), .B(SHA256_result[189]), .S0(n438), .Y(
        mux1[29]) );
  MX2X1 U2478 ( .A(SHA256_result[158]), .B(SHA256_result[190]), .S0(n438), .Y(
        mux1[30]) );
  MX2XL U2479 ( .A(SHA256_result[16]), .B(SHA256_result[48]), .S0(
        mux_control_0_), .Y(mux2[16]) );
  MX2XL U2480 ( .A(SHA256_result[19]), .B(SHA256_result[51]), .S0(
        mux_control_0_), .Y(mux2[19]) );
  MX2XL U2481 ( .A(SHA256_result[18]), .B(SHA256_result[50]), .S0(
        mux_control_0_), .Y(mux2[18]) );
  MX2XL U2482 ( .A(SHA256_result[20]), .B(SHA256_result[52]), .S0(
        mux_control_0_), .Y(mux2[20]) );
  INVX1 U2483 ( .A(SHA256_result[3]), .Y(n1213) );
  MX2X1 U2484 ( .A(SHA256_result[63]), .B(SHA256_result[95]), .S0(n106), .Y(
        f1_EFG_32[31]) );
  NOR3X1 U2485 ( .A(n2938), .B(n425), .C(n1304), .Y(n4011) );
  OAI222XL U2486 ( .A0(n4050), .A1(n2906), .B0(n4051), .B1(n1287), .C0(n422), 
        .C1(n4052), .Y(n4049) );
  OAI21XL U2487 ( .A0(n431), .A1(n1251), .B0(n290), .Y(n4053) );
  OAI222XL U2488 ( .A0(n2938), .A1(n3992), .B0(n1306), .B1(n4040), .C0(n1275), 
        .C1(n4094), .Y(n4163) );
  OAI222XL U2489 ( .A0(n2906), .A1(n4010), .B0(n289), .B1(n1257), .C0(n425), 
        .C1(n3999), .Y(n4112) );
  OR2X2 U2490 ( .A(read_counter[1]), .B(read_counter[0]), .Y(n1239) );
  AOI22XL U2491 ( .A0(n3694), .A1(SHA256_result[113]), .B0(n3695), .B1(
        SHA256_result[117]), .Y(n3834) );
  MX2X1 U2492 ( .A(SHA256_result[30]), .B(SHA256_result[62]), .S0(
        mux_control_0_), .Y(mux2[30]) );
  NAND4X1 U2493 ( .A(n3686), .B(n3687), .C(n3688), .D(n3689), .Y(n3685) );
  AOI22XL U2494 ( .A0(n3696), .A1(n123), .B0(n3697), .B1(n106), .Y(n3686) );
  NAND4X1 U2495 ( .A(n3875), .B(n3876), .C(n3877), .D(n3878), .Y(n3874) );
  AOI22XL U2496 ( .A0(n3696), .A1(n103), .B0(n3697), .B1(n94), .Y(n3875) );
  AOI22XL U2497 ( .A0(n3694), .A1(SHA256_result[112]), .B0(n3695), .B1(
        SHA256_result[116]), .Y(n3876) );
  NAND4X1 U2498 ( .A(n3791), .B(n3792), .C(n3793), .D(n3794), .Y(n3790) );
  AOI22XL U2499 ( .A0(n3696), .A1(n118), .B0(n3697), .B1(n115), .Y(n3791) );
  AOI22XL U2500 ( .A0(n3694), .A1(n291), .B0(n3695), .B1(SHA256_result[118]), 
        .Y(n3792) );
  NAND4X1 U2501 ( .A(n3841), .B(n3842), .C(n3843), .D(n3844), .Y(n3830) );
  AOI22XL U2502 ( .A0(n3718), .A1(SHA256_result[49]), .B0(n3719), .B1(
        SHA256_result[53]), .Y(n3842) );
  NAND4X1 U2503 ( .A(n3895), .B(n3896), .C(n3897), .D(n3898), .Y(n3872) );
  AOI22XL U2504 ( .A0(n3718), .A1(SHA256_result[48]), .B0(n3719), .B1(
        SHA256_result[52]), .Y(n3896) );
  NAND4X1 U2505 ( .A(n3799), .B(n3800), .C(n3801), .D(n3802), .Y(n3788) );
  AOI22XL U2506 ( .A0(n3718), .A1(SHA256_result[50]), .B0(n3719), .B1(
        SHA256_result[54]), .Y(n3800) );
  NAND4X1 U2507 ( .A(n3710), .B(n3711), .C(n3712), .D(n3713), .Y(n3683) );
  AOI22XL U2508 ( .A0(n3718), .A1(SHA256_result[51]), .B0(n3719), .B1(
        SHA256_result[55]), .Y(n3711) );
  NAND4X1 U2509 ( .A(n3885), .B(n3886), .C(n3887), .D(n3888), .Y(n3873) );
  AOI22XL U2510 ( .A0(n3706), .A1(SHA256_result[80]), .B0(n3707), .B1(
        SHA256_result[84]), .Y(n3886) );
  NAND4X1 U2511 ( .A(n3837), .B(n3838), .C(n3839), .D(n3840), .Y(n3831) );
  AOI22XL U2512 ( .A0(n3706), .A1(SHA256_result[81]), .B0(n3707), .B1(
        SHA256_result[85]), .Y(n3838) );
  NAND4X1 U2513 ( .A(n3795), .B(n3796), .C(n3797), .D(n3798), .Y(n3789) );
  AOI22XL U2514 ( .A0(n3706), .A1(SHA256_result[82]), .B0(n3707), .B1(
        SHA256_result[86]), .Y(n3796) );
  NAND4X1 U2515 ( .A(n3698), .B(n3699), .C(n3700), .D(n3701), .Y(n3684) );
  AOI22XL U2516 ( .A0(n3706), .A1(SHA256_result[83]), .B0(n3707), .B1(
        SHA256_result[87]), .Y(n3699) );
  NAND4X1 U2517 ( .A(n3913), .B(n3914), .C(n3915), .D(n3916), .Y(n3912) );
  AOI22XL U2518 ( .A0(n3743), .A1(n18), .B0(n3744), .B1(SHA256_result[236]), 
        .Y(n3915) );
  NAND4X1 U2519 ( .A(n3927), .B(n3928), .C(n3929), .D(n3930), .Y(n3910) );
  AOI22XL U2520 ( .A0(n3767), .A1(SHA256_result[168]), .B0(n3768), .B1(
        SHA256_result[172]), .Y(n3929) );
  NAND4X1 U2521 ( .A(n3861), .B(n3862), .C(n3863), .D(n3864), .Y(n3850) );
  AOI22XL U2522 ( .A0(n3767), .A1(SHA256_result[169]), .B0(n3768), .B1(
        SHA256_result[173]), .Y(n3863) );
  NAND4X1 U2523 ( .A(n3819), .B(n3820), .C(n3821), .D(n3822), .Y(n3808) );
  AOI22XL U2524 ( .A0(n3767), .A1(SHA256_result[170]), .B0(n3768), .B1(
        SHA256_result[174]), .Y(n3821) );
  NAND4X1 U2525 ( .A(n3761), .B(n3762), .C(n3763), .D(n3764), .Y(n3734) );
  AOI22XL U2526 ( .A0(n3767), .A1(SHA256_result[171]), .B0(n3768), .B1(
        SHA256_result[175]), .Y(n3763) );
  NAND4X1 U2527 ( .A(n3921), .B(n3922), .C(n3923), .D(n3924), .Y(n3911) );
  AOI22XL U2528 ( .A0(n3755), .A1(SHA256_result[200]), .B0(n3756), .B1(
        SHA256_result[204]), .Y(n3923) );
  NAND4X1 U2529 ( .A(n3857), .B(n3858), .C(n3859), .D(n3860), .Y(n3851) );
  AOI22XL U2530 ( .A0(n3755), .A1(SHA256_result[201]), .B0(n3756), .B1(
        SHA256_result[205]), .Y(n3859) );
  NAND4X1 U2531 ( .A(n3815), .B(n3816), .C(n3817), .D(n3818), .Y(n3809) );
  AOI22XL U2532 ( .A0(n3755), .A1(SHA256_result[202]), .B0(n3756), .B1(
        SHA256_result[206]), .Y(n3817) );
  NAND4X1 U2533 ( .A(n3749), .B(n3750), .C(n3751), .D(n3752), .Y(n3735) );
  AOI22XL U2534 ( .A0(n3755), .A1(SHA256_result[203]), .B0(n3756), .B1(
        SHA256_result[207]), .Y(n3751) );
  NAND4X1 U2535 ( .A(n3903), .B(n3904), .C(n3905), .D(n3906), .Y(n3871) );
  AOI22X1 U2536 ( .A0(n3729), .A1(SHA256_result[16]), .B0(n3730), .B1(
        SHA256_result[20]), .Y(n3904) );
  AOI22X1 U2537 ( .A0(n3731), .A1(SHA256_result[24]), .B0(n3732), .B1(
        SHA256_result[28]), .Y(n3903) );
  NAND4X1 U2538 ( .A(n3845), .B(n3846), .C(n3847), .D(n3848), .Y(n3829) );
  AOI22X1 U2539 ( .A0(n3729), .A1(SHA256_result[17]), .B0(n3730), .B1(
        SHA256_result[21]), .Y(n3846) );
  AOI22X1 U2540 ( .A0(n3731), .A1(SHA256_result[25]), .B0(n3732), .B1(
        SHA256_result[29]), .Y(n3845) );
  NAND4X1 U2541 ( .A(n3803), .B(n3804), .C(n3805), .D(n3806), .Y(n3787) );
  AOI22X1 U2542 ( .A0(n3729), .A1(SHA256_result[18]), .B0(n3730), .B1(
        SHA256_result[22]), .Y(n3804) );
  AOI22X1 U2543 ( .A0(n3731), .A1(SHA256_result[26]), .B0(n3732), .B1(
        SHA256_result[30]), .Y(n3803) );
  NAND4X1 U2544 ( .A(n3722), .B(n3723), .C(n3724), .D(n3725), .Y(n3682) );
  AOI22X1 U2545 ( .A0(n3729), .A1(SHA256_result[19]), .B0(n3730), .B1(
        SHA256_result[23]), .Y(n3723) );
  AOI22X1 U2546 ( .A0(n3731), .A1(SHA256_result[27]), .B0(n3732), .B1(
        SHA256_result[31]), .Y(n3722) );
  NOR2X1 U2547 ( .A(read_counter[5]), .B(read_counter[0]), .Y(n3893) );
  NOR2X1 U2548 ( .A(read_counter[4]), .B(read_counter[1]), .Y(n3907) );
  NOR2X1 U2549 ( .A(n1431), .B(read_counter[0]), .Y(n3926) );
  NOR2X1 U2550 ( .A(n1429), .B(read_counter[4]), .Y(n3908) );
  OAI21XL U2551 ( .A0(n4205), .A1(n2925), .B0(n4206), .Y(n4204) );
  AOI211X1 U2552 ( .A0(n258), .A1(n429), .B0(n3946), .C0(n4122), .Y(n4205) );
  OAI21XL U2553 ( .A0(n1265), .A1(n249), .B0(n4055), .Y(n4206) );
  NAND2X1 U2554 ( .A(n4039), .B(n2938), .Y(n4173) );
  MX2X1 U2555 ( .A(SHA256_result[29]), .B(SHA256_result[61]), .S0(
        mux_control_0_), .Y(mux2[29]) );
  AOI22XL U2556 ( .A0(n3741), .A1(n222), .B0(n3742), .B1(n219), .Y(n3740) );
  AOI22XL U2557 ( .A0(n3741), .A1(n317), .B0(n3742), .B1(n88), .Y(n3916) );
  AOI22XL U2558 ( .A0(n3753), .A1(n96), .B0(n3754), .B1(SHA256_result[196]), 
        .Y(n3924) );
  AOI22XL U2559 ( .A0(n3753), .A1(SHA256_result[194]), .B0(n3754), .B1(
        SHA256_result[198]), .Y(n3818) );
  AOI22XL U2560 ( .A0(n3753), .A1(n100), .B0(n3754), .B1(SHA256_result[199]), 
        .Y(n3752) );
  AOI22XL U2561 ( .A0(n3765), .A1(SHA256_result[160]), .B0(n3766), .B1(
        SHA256_result[164]), .Y(n3930) );
  AOI22XL U2562 ( .A0(n3753), .A1(SHA256_result[193]), .B0(n3754), .B1(
        SHA256_result[197]), .Y(n3860) );
  AOI22XL U2563 ( .A0(n3765), .A1(SHA256_result[161]), .B0(n3766), .B1(
        SHA256_result[165]), .Y(n3864) );
  AOI22XL U2564 ( .A0(n3765), .A1(SHA256_result[162]), .B0(n3766), .B1(
        SHA256_result[166]), .Y(n3822) );
  AOI22XL U2565 ( .A0(n3765), .A1(SHA256_result[163]), .B0(n3766), .B1(
        SHA256_result[167]), .Y(n3764) );
  AOI22X1 U2566 ( .A0(n3781), .A1(SHA256_result[144]), .B0(n3782), .B1(
        SHA256_result[148]), .Y(n3936) );
  AOI22X1 U2567 ( .A0(n3781), .A1(SHA256_result[145]), .B0(n3782), .B1(
        SHA256_result[149]), .Y(n3866) );
  AOI22X1 U2568 ( .A0(n3781), .A1(SHA256_result[146]), .B0(n3782), .B1(
        SHA256_result[150]), .Y(n3824) );
  AOI22X1 U2569 ( .A0(n3781), .A1(SHA256_result[147]), .B0(n3782), .B1(
        SHA256_result[151]), .Y(n3774) );
  AOI22X1 U2570 ( .A0(n3783), .A1(SHA256_result[152]), .B0(n3784), .B1(
        SHA256_result[156]), .Y(n3935) );
  AOI22X1 U2571 ( .A0(n3783), .A1(SHA256_result[153]), .B0(n3784), .B1(
        SHA256_result[157]), .Y(n3865) );
  AOI22X1 U2572 ( .A0(n3783), .A1(SHA256_result[154]), .B0(n3784), .B1(
        SHA256_result[158]), .Y(n3823) );
  AOI22X1 U2573 ( .A0(n3783), .A1(SHA256_result[155]), .B0(n3784), .B1(
        SHA256_result[159]), .Y(n3773) );
  OAI2BB2X1 U2574 ( .B0(n4121), .B1(n1306), .A0N(n260), .A1N(n3964), .Y(n4119)
         );
  AOI211X1 U2575 ( .A0(n425), .A1(n2938), .B0(n4027), .C0(n4122), .Y(n4121) );
  MX2X1 U2576 ( .A(SHA256_result[28]), .B(SHA256_result[60]), .S0(
        mux_control_0_), .Y(mux2[28]) );
  INVX1 U2577 ( .A(read_counter[2]), .Y(n1430) );
  INVX1 U2578 ( .A(read_counter[1]), .Y(n1429) );
  INVX1 U2579 ( .A(read_counter[5]), .Y(n1431) );
  INVXL U2580 ( .A(n18), .Y(n1164) );
  INVXL U2581 ( .A(SHA256_result[228]), .Y(n1181) );
  INVXL U2582 ( .A(SHA256_result[200]), .Y(n1312) );
  INVXL U2583 ( .A(SHA256_result[193]), .Y(n1307) );
  INVXL U2584 ( .A(SHA256_result[206]), .Y(n1316) );
  INVXL U2585 ( .A(SHA256_result[204]), .Y(n1314) );
  INVXL U2586 ( .A(SHA256_result[198]), .Y(n1311) );
  INVXL U2587 ( .A(SHA256_result[197]), .Y(n1310) );
  INVXL U2588 ( .A(SHA256_result[196]), .Y(n1309) );
  INVXL U2589 ( .A(SHA256_result[118]), .Y(n722) );
  INVXL U2590 ( .A(SHA256_result[117]), .Y(n1370) );
  INVXL U2591 ( .A(SHA256_result[116]), .Y(n1369) );
  INVXL U2592 ( .A(SHA256_result[171]), .Y(n937) );
  INVX1 U2593 ( .A(SHA256_result[63]), .Y(n1403) );
  INVX1 U2594 ( .A(SHA256_result[222]), .Y(n1238) );
  INVX1 U2595 ( .A(SHA256_result[191]), .Y(n1328) );
  INVX1 U2596 ( .A(SHA256_result[190]), .Y(n1345) );
  INVXL U2597 ( .A(SHA256_result[51]), .Y(n1392) );
  INVXL U2598 ( .A(SHA256_result[50]), .Y(n1391) );
  INVXL U2599 ( .A(SHA256_result[52]), .Y(n1393) );
  INVX1 U2600 ( .A(SHA256_result[61]), .Y(n1401) );
  INVXL U2601 ( .A(SHA256_result[83]), .Y(n1375) );
  INVX1 U2602 ( .A(SHA256_result[94]), .Y(n1386) );
  INVXL U2603 ( .A(SHA256_result[86]), .Y(n1378) );
  INVXL U2604 ( .A(SHA256_result[85]), .Y(n1377) );
  INVXL U2605 ( .A(SHA256_result[84]), .Y(n1376) );
  INVX1 U2606 ( .A(SHA256_result[93]), .Y(n1385) );
  INVXL U2607 ( .A(SHA256_result[68]), .Y(n668) );
  INVXL U2608 ( .A(n94), .Y(n705) );
  INVXL U2609 ( .A(SHA256_result[207]), .Y(n1317) );
  INVXL U2610 ( .A(SHA256_result[205]), .Y(n1315) );
  INVXL U2611 ( .A(SHA256_result[201]), .Y(n1313) );
  INVX1 U2612 ( .A(SHA256_result[221]), .Y(n1237) );
  INVX1 U2613 ( .A(SHA256_result[220]), .Y(n1236) );
  INVX1 U2614 ( .A(SHA256_result[189]), .Y(n1344) );
  INVXL U2615 ( .A(SHA256_result[175]), .Y(n1331) );
  INVXL U2616 ( .A(SHA256_result[174]), .Y(n1330) );
  INVXL U2617 ( .A(SHA256_result[173]), .Y(n1329) );
  INVX1 U2618 ( .A(SHA256_result[188]), .Y(n1343) );
  INVXL U2619 ( .A(SHA256_result[172]), .Y(n933) );
  INVXL U2620 ( .A(SHA256_result[49]), .Y(n1390) );
  INVXL U2621 ( .A(SHA256_result[48]), .Y(n1389) );
  INVXL U2622 ( .A(SHA256_result[82]), .Y(n1374) );
  INVX1 U2623 ( .A(SHA256_result[95]), .Y(n1387) );
  AOI22XL U2624 ( .A0(n3694), .A1(n111), .B0(n3695), .B1(n90), .Y(n3687) );
  XOR3X2 U2625 ( .A(n136), .B(n111), .C(n102), .Y(f4_E_32[13]) );
  NAND2XL U2626 ( .A(SHA256_result[73]), .B(n323), .Y(n655) );
  AOI22XL U2627 ( .A0(n3704), .A1(SHA256_result[73]), .B0(n3705), .B1(
        SHA256_result[77]), .Y(n3839) );
  AOI21XL U2628 ( .A0(n232), .A1(n343), .B0(n327), .Y(n603) );
  NAND2XL U2629 ( .A(n85), .B(n323), .Y(n658) );
  AOI22XL U2630 ( .A0(n3704), .A1(n85), .B0(n3705), .B1(SHA256_result[76]), 
        .Y(n3887) );
  MX2XL U2631 ( .A(SHA256_result[14]), .B(SHA256_result[46]), .S0(
        mux_control_0_), .Y(mux2[14]) );
  AOI22XL U2632 ( .A0(n3704), .A1(SHA256_result[74]), .B0(n3705), .B1(
        SHA256_result[78]), .Y(n3797) );
  AOI21XL U2633 ( .A0(n207), .A1(n341), .B0(n328), .Y(n671) );
  INVX8 U2634 ( .A(SHA256_result[38]), .Y(n1206) );
  INVXL U2635 ( .A(n210), .Y(n768) );
  AOI22XL U2636 ( .A0(n3692), .A1(n210), .B0(n3693), .B1(n147), .Y(n3877) );
  XOR3X2 U2637 ( .A(n210), .B(SHA256_result[117]), .C(n118), .Y(f4_E_32[15])
         );
  XOR3X2 U2638 ( .A(n210), .B(n171), .C(n122), .Y(f4_E_32[2]) );
  XOR3X2 U2639 ( .A(n150), .B(n202), .C(n103), .Y(f4_E_32[31]) );
  XOR3X2 U2640 ( .A(n202), .B(n90), .C(n94), .Y(f4_E_32[17]) );
  INVXL U2641 ( .A(n283), .Y(n784) );
  AOI21XL U2642 ( .A0(n283), .A1(n341), .B0(n329), .Y(n785) );
  AOI21XL U2643 ( .A0(n213), .A1(n341), .B0(n328), .Y(n673) );
  AOI22XL U2644 ( .A0(n3702), .A1(n213), .B0(n3703), .B1(n84), .Y(n3798) );
  AOI22XL U2645 ( .A0(n3692), .A1(n139), .B0(n3693), .B1(n280), .Y(n3688) );
  XOR3X2 U2646 ( .A(n139), .B(SHA256_result[112]), .C(n114), .Y(f4_E_32[5]) );
  AOI22XL U2647 ( .A0(n3704), .A1(SHA256_result[75]), .B0(n3705), .B1(
        SHA256_result[79]), .Y(n3700) );
  AOI21XL U2648 ( .A0(n184), .A1(n342), .B0(n327), .Y(n584) );
  MX2XL U2649 ( .A(SHA256_result[8]), .B(n184), .S0(mux_control_0_), .Y(
        mux2[8]) );
  AOI22XL U2650 ( .A0(n3716), .A1(n184), .B0(n3717), .B1(SHA256_result[44]), 
        .Y(n3897) );
  AOI21XL U2651 ( .A0(n134), .A1(n342), .B0(n327), .Y(n586) );
  MX2XL U2652 ( .A(SHA256_result[7]), .B(n134), .S0(mux_control_0_), .Y(
        mux2[7]) );
  AOI21XL U2653 ( .A0(n167), .A1(n341), .B0(n328), .Y(n659) );
  AOI22XL U2654 ( .A0(n3702), .A1(n207), .B0(n3703), .B1(n167), .Y(n3701) );
  NAND2XL U2655 ( .A(n203), .B(n345), .Y(n747) );
  AOI22XL U2656 ( .A0(n3692), .A1(n202), .B0(n3693), .B1(n203), .Y(n3793) );
  NAND2BXL U2657 ( .AN(n332), .B(n209), .Y(n712) );
  NAND2XL U2658 ( .A(n74), .B(n323), .Y(n595) );
  AOI22XL U2659 ( .A0(n3714), .A1(n232), .B0(n3715), .B1(n74), .Y(n3898) );
  INVX8 U2660 ( .A(n231), .Y(n1217) );
  NAND2XL U2661 ( .A(n159), .B(n323), .Y(n580) );
  MX2XL U2662 ( .A(SHA256_result[10]), .B(n159), .S0(mux_control_0_), .Y(
        mux2[10]) );
  AOI22XL U2663 ( .A0(n3716), .A1(n159), .B0(n3717), .B1(SHA256_result[46]), 
        .Y(n3801) );
  AOI21XL U2664 ( .A0(SHA256_result[43]), .A1(n342), .B0(n327), .Y(n576) );
  MX2XL U2665 ( .A(SHA256_result[11]), .B(SHA256_result[43]), .S0(
        mux_control_0_), .Y(mux2[11]) );
  AOI22XL U2666 ( .A0(n3716), .A1(SHA256_result[43]), .B0(n3717), .B1(
        SHA256_result[47]), .Y(n3712) );
  NAND2XL U2667 ( .A(n165), .B(n323), .Y(n583) );
  MX2XL U2668 ( .A(SHA256_result[9]), .B(n165), .S0(mux_control_0_), .Y(
        mux2[9]) );
  AOI22XL U2669 ( .A0(n3716), .A1(n165), .B0(n3717), .B1(SHA256_result[45]), 
        .Y(n3843) );
  INVXL U2670 ( .A(n281), .Y(n763) );
  NAND2XL U2671 ( .A(n281), .B(n345), .Y(n764) );
  AOI22XL U2672 ( .A0(n3692), .A1(n281), .B0(n3693), .B1(n171), .Y(n3835) );
  XOR3X2 U2673 ( .A(n292), .B(n281), .C(n90), .Y(f4_E_32[30]) );
  XOR3X2 U2674 ( .A(n281), .B(SHA256_result[118]), .C(n123), .Y(f4_E_32[16])
         );
  XOR3X2 U2675 ( .A(n281), .B(n203), .C(n93), .Y(f4_E_32[3]) );
  AOI22XL U2676 ( .A0(n3696), .A1(n244), .B0(n3697), .B1(n110), .Y(n3833) );
  MX2XL U2677 ( .A(SHA256_result[61]), .B(SHA256_result[93]), .S0(n110), .Y(
        f1_EFG_32[29]) );
  XOR3X2 U2678 ( .A(n126), .B(n280), .C(n109), .Y(f4_E_32[4]) );
  XOR3X2 U2679 ( .A(n139), .B(n103), .C(n110), .Y(f4_E_32[18]) );
  NAND4X1 U2680 ( .A(n3833), .B(n3834), .C(n3835), .D(n3836), .Y(n3832) );
  OAI21XL U2681 ( .A0(n420), .A1(n703), .B0(n702), .Y(n4509) );
  OAI211X1 U2682 ( .A0(n332), .A1(n703), .B0(n611), .C0(n610), .Y(n4414) );
  OAI21XL U2683 ( .A0(n420), .A1(n141), .B0(n598), .Y(n4377) );
  NAND2XL U2684 ( .A(n234), .B(n323), .Y(n600) );
  MXI2XL U2685 ( .A(n1215), .B(n141), .S0(mux_control_0_), .Y(mux2[2]) );
  AOI22XL U2686 ( .A0(n3690), .A1(n283), .B0(n3691), .B1(n154), .Y(n3689) );
  XOR3X2 U2687 ( .A(n154), .B(SHA256_result[116]), .C(n244), .Y(f4_E_32[14])
         );
  NAND2XL U2688 ( .A(n181), .B(n323), .Y(n677) );
  AOI22XL U2689 ( .A0(n3702), .A1(n181), .B0(n3703), .B1(n129), .Y(n3840) );
  AOI21XL U2690 ( .A0(n185), .A1(n341), .B0(n329), .Y(n789) );
  AOI22XL U2691 ( .A0(n3690), .A1(n185), .B0(n3691), .B1(n136), .Y(n3794) );
  XOR3X2 U2692 ( .A(n185), .B(n154), .C(SHA256_result[117]), .Y(f4_E_32[28])
         );
  XOR3X2 U2693 ( .A(n185), .B(SHA256_result[112]), .C(n110), .Y(f4_E_32[23])
         );
  XOR3X2 U2694 ( .A(n282), .B(n280), .C(SHA256_result[116]), .Y(f4_E_32[9]) );
  XOR3X2 U2695 ( .A(n283), .B(n210), .C(SHA256_result[118]), .Y(f4_E_32[29])
         );
  MXI2XL U2696 ( .A(n1218), .B(n1217), .S0(mux_control_0_), .Y(mux2[0]) );
  AOI21XL U2697 ( .A0(n158), .A1(n341), .B0(n329), .Y(n792) );
  AOI22XL U2698 ( .A0(n3690), .A1(n158), .B0(n3691), .B1(n150), .Y(n3836) );
  XOR3X2 U2699 ( .A(n158), .B(n136), .C(SHA256_result[116]), .Y(f4_E_32[27])
         );
  XOR3X2 U2700 ( .A(n158), .B(n280), .C(n94), .Y(f4_E_32[22]) );
  XOR3X2 U2701 ( .A(n158), .B(n203), .C(n111), .Y(f4_E_32[8]) );
  XOR3X2 U2702 ( .A(n283), .B(SHA256_result[112]), .C(SHA256_result[117]), .Y(
        f4_E_32[10]) );
  XOR3X2 U2703 ( .A(n283), .B(SHA256_result[113]), .C(n115), .Y(f4_E_32[24])
         );
  NAND2XL U2704 ( .A(n239), .B(n323), .Y(n680) );
  AOI22XL U2705 ( .A0(n3702), .A1(n239), .B0(n3703), .B1(SHA256_result[68]), 
        .Y(n3888) );
  INVX4 U2706 ( .A(n238), .Y(n699) );
  NAND2BXL U2707 ( .AN(n331), .B(next_E[29]), .Y(n704) );
  NAND2XL U2708 ( .A(n143), .B(n323), .Y(n590) );
  AOI22XL U2709 ( .A0(n3714), .A1(n234), .B0(n3715), .B1(n143), .Y(n3802) );
  AOI21XL U2710 ( .A0(n285), .A1(n341), .B0(n799), .Y(n801) );
  AOI22XL U2711 ( .A0(n3690), .A1(n285), .B0(n3691), .B1(n292), .Y(n3878) );
  XOR3X2 U2712 ( .A(n285), .B(n150), .C(n111), .Y(f4_E_32[26]) );
  XOR3X2 U2713 ( .A(n285), .B(n203), .C(n123), .Y(f4_E_32[21]) );
  XOR3X2 U2714 ( .A(n285), .B(n171), .C(n291), .Y(f4_E_32[7]) );
  AOI22XL U2715 ( .A0(n3714), .A1(n208), .B0(n3715), .B1(n134), .Y(n3713) );
  NAND2BXL U2716 ( .AN(n332), .B(n188), .Y(n714) );
  AOI21XL U2717 ( .A0(n164), .A1(n342), .B0(n327), .Y(n601) );
  AOI22XL U2718 ( .A0(n3714), .A1(n164), .B0(n3715), .B1(n174), .Y(n3844) );
  NAND2BXL U2719 ( .AN(n330), .B(next_E[21]), .Y(n725) );
  MX2X4 U2720 ( .A(SHA256_result[50]), .B(SHA256_result[82]), .S0(n291), .Y(
        f1_EFG_32[18]) );
  MX2X4 U2721 ( .A(SHA256_result[49]), .B(SHA256_result[81]), .S0(
        SHA256_result[113]), .Y(f1_EFG_32[17]) );
  MX2X4 U2722 ( .A(SHA256_result[48]), .B(SHA256_result[80]), .S0(
        SHA256_result[112]), .Y(f1_EFG_32[16]) );
  MX2X4 U2723 ( .A(SHA256_result[47]), .B(SHA256_result[79]), .S0(n280), .Y(
        f1_EFG_32[15]) );
  MXI2X4 U2724 ( .A(n682), .B(n681), .S0(SHA256_result[110]), .Y(f1_EFG_32[14]) );
  MXI2X4 U2725 ( .A(n686), .B(n685), .S0(n146), .Y(f1_EFG_32[12]) );
  MXI2X4 U2726 ( .A(n688), .B(n687), .S0(n138), .Y(f1_EFG_32[11]) );
  MXI2X4 U2727 ( .A(n160), .B(n689), .S0(n126), .Y(f1_EFG_32[10]) );
  MXI2X4 U2728 ( .A(n166), .B(n690), .S0(SHA256_result[105]), .Y(f1_EFG_32[9])
         );
  MXI2X4 U2729 ( .A(n183), .B(n691), .S0(SHA256_result[104]), .Y(f1_EFG_32[8])
         );
  MXI2X4 U2730 ( .A(n692), .B(n168), .S0(n153), .Y(f1_EFG_32[7]) );
  NAND2X4 U2731 ( .A(SHA256_result[102]), .B(n83), .Y(n693) );
  OAI21X4 U2732 ( .A0(SHA256_result[102]), .A1(n1206), .B0(n693), .Y(
        f1_EFG_32[6]) );
  NAND2X4 U2733 ( .A(n129), .B(n149), .Y(n694) );
  OAI21X4 U2734 ( .A0(n149), .A1(n1208), .B0(n694), .Y(f1_EFG_32[5]) );
  NAND2X4 U2735 ( .A(SHA256_result[68]), .B(SHA256_result[100]), .Y(n695) );
  OAI21X4 U2736 ( .A0(SHA256_result[100]), .A1(n1210), .B0(n695), .Y(
        f1_EFG_32[4]) );
  MXI2X4 U2737 ( .A(n1212), .B(n696), .S0(n68), .Y(f1_EFG_32[3]) );
  MXI2X4 U2738 ( .A(n1214), .B(n697), .S0(SHA256_result[98]), .Y(f1_EFG_32[2])
         );
  MXI2X4 U2739 ( .A(n182), .B(n698), .S0(n157), .Y(f1_EFG_32[1]) );
  MXI2X4 U2740 ( .A(n1217), .B(n699), .S0(SHA256_result[96]), .Y(f1_EFG_32[0])
         );
  NAND2X4 U2741 ( .A(N948), .B(n807), .Y(n759) );
  OAI2BB1X4 U2742 ( .A0N(SHA256_result[205]), .A1N(SHA256_result[237]), .B0(
        n1070), .Y(f2_ABC_32[13]) );
  OAI2BB1X4 U2743 ( .A0N(SHA256_result[204]), .A1N(SHA256_result[236]), .B0(
        n1071), .Y(f2_ABC_32[12]) );
  OAI2BB1X4 U2744 ( .A0N(SHA256_result[203]), .A1N(n16), .B0(n1072), .Y(
        f2_ABC_32[11]) );
  OAI21X4 U2745 ( .A0(n311), .A1(SHA256_result[202]), .B0(SHA256_result[170]), 
        .Y(n1073) );
  OAI2BB1X4 U2746 ( .A0N(SHA256_result[202]), .A1N(n311), .B0(n1073), .Y(
        f2_ABC_32[10]) );
  OAI21X4 U2747 ( .A0(n312), .A1(SHA256_result[201]), .B0(SHA256_result[169]), 
        .Y(n1074) );
  OAI21X4 U2748 ( .A0(n218), .A1(SHA256_result[199]), .B0(SHA256_result[167]), 
        .Y(n1076) );
  OAI21X4 U2749 ( .A0(SHA256_result[198]), .A1(n313), .B0(SHA256_result[166]), 
        .Y(n1077) );
  OAI2BB1X4 U2750 ( .A0N(SHA256_result[198]), .A1N(n313), .B0(n1077), .Y(
        f2_ABC_32[6]) );
  OAI21X4 U2751 ( .A0(SHA256_result[197]), .A1(n314), .B0(SHA256_result[165]), 
        .Y(n1078) );
  OAI2BB1X4 U2752 ( .A0N(SHA256_result[197]), .A1N(n314), .B0(n1078), .Y(
        f2_ABC_32[5]) );
  OAI2BB1X4 U2753 ( .A0N(SHA256_result[196]), .A1N(SHA256_result[228]), .B0(
        n1079), .Y(f2_ABC_32[4]) );
  OAI2BB1X4 U2754 ( .A0N(SHA256_result[194]), .A1N(n315), .B0(n1081), .Y(
        f2_ABC_32[2]) );
  OAI2BB1X4 U2755 ( .A0N(n96), .A1N(n317), .B0(n1083), .Y(f2_ABC_32[0]) );
  OAI2BB1X1 U2756 ( .A0N(read_counter[0]), .A1N(read_counter[1]), .B0(n1239), 
        .Y(N3564) );
  OR2X1 U2757 ( .A(n1239), .B(read_counter[2]), .Y(n1240) );
  OAI2BB1X1 U2758 ( .A0N(n1239), .A1N(read_counter[2]), .B0(n1240), .Y(N3565)
         );
  OR2X1 U2759 ( .A(n1240), .B(read_counter[3]), .Y(n1241) );
  OAI2BB1X1 U2760 ( .A0N(n1240), .A1N(read_counter[3]), .B0(n1241), .Y(N3566)
         );
  NOR2X1 U2761 ( .A(read_counter[4]), .B(n1241), .Y(n1242) );
endmodule


module controller_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module controller_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module controller ( clk, reset, first_block, last_block, output_enable, busy, 
        inner_busy, first_block_core );
  input clk, reset, first_block, last_block;
  output output_enable, busy, inner_busy, first_block_core;
  wire   N13, N14, N24, N25, N26, N27, N28, N29, N30, N45, N46, N47, N48, N49,
         N50, N51, N52, n26, n27, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38;
  wire   [1:0] state;
  wire   [7:0] counter2;
  wire   [6:0] counter1;

  CLKINVX4 U29 ( .A(reset), .Y(n27) );
  controller_DW01_inc_0 add_97 ( .A(counter2), .SUM({N52, N51, N50, N49, N48, 
        N47, N46, N45}) );
  controller_DW01_inc_1 add_83 ( .A(counter1), .SUM({N30, N29, N28, N27, N26, 
        N25, N24}) );
  DFFTRX1 counter2_reg_0_ ( .D(N45), .RN(n37), .CK(clk), .Q(counter2[0]), .QN(
        n26) );
  DFFTRX1 counter1_reg_2_ ( .D(N26), .RN(n38), .CK(clk), .Q(counter1[2]), .QN(
        n2) );
  DFFTRX1 counter1_reg_3_ ( .D(N27), .RN(n38), .CK(clk), .Q(counter1[3]), .QN(
        n1) );
  DFFTRX1 counter1_reg_4_ ( .D(N28), .RN(n38), .CK(clk), .Q(counter1[4]), .QN(
        n14) );
  DFFTRX1 counter1_reg_5_ ( .D(N29), .RN(n38), .CK(clk), .Q(counter1[5]), .QN(
        n13) );
  DFFTRX1 counter1_reg_0_ ( .D(N24), .RN(n38), .CK(clk), .Q(counter1[0]), .QN(
        n4) );
  DFFTRX1 counter1_reg_6_ ( .D(N30), .RN(n38), .CK(clk), .Q(counter1[6]), .QN(
        n12) );
  DFFTRX1 counter1_reg_1_ ( .D(N25), .RN(n38), .CK(clk), .Q(counter1[1]), .QN(
        n3) );
  DFFTRX1 counter2_reg_3_ ( .D(N48), .RN(n37), .CK(clk), .Q(counter2[3]), .QN(
        n9) );
  DFFTRX1 counter2_reg_5_ ( .D(N50), .RN(n37), .CK(clk), .Q(counter2[5]), .QN(
        n7) );
  DFFTRX1 counter2_reg_4_ ( .D(N49), .RN(n37), .CK(clk), .Q(counter2[4]), .QN(
        n8) );
  DFFTRX1 counter2_reg_1_ ( .D(N46), .RN(n37), .CK(clk), .Q(counter2[1]), .QN(
        n11) );
  DFFHQX1 state_reg_0_ ( .D(N13), .CK(clk), .Q(state[0]) );
  DFFTRX1 counter2_reg_2_ ( .D(N47), .RN(n37), .CK(clk), .Q(counter2[2]), .QN(
        n10) );
  DFFTRX1 counter2_reg_6_ ( .D(N51), .RN(n37), .CK(clk), .Q(counter2[6]), .QN(
        n6) );
  DFFTRX1 counter2_reg_7_ ( .D(N52), .RN(n37), .CK(clk), .Q(counter2[7]), .QN(
        n5) );
  DFFXL state_reg_1_ ( .D(N14), .CK(clk), .Q(state[1]), .QN(n34) );
  NAND3X1 U3 ( .A(n8), .B(n7), .C(n9), .Y(n19) );
  NOR2X1 U4 ( .A(n34), .B(state[0]), .Y(inner_busy) );
  NOR2X1 U5 ( .A(n5), .B(n15), .Y(output_enable) );
  MXI2X1 U6 ( .A(n16), .B(n17), .S0(n6), .Y(n15) );
  NOR2X1 U7 ( .A(n11), .B(n10), .Y(n18) );
  MXI2XL U8 ( .A(n23), .B(n24), .S0(n6), .Y(n21) );
  NAND2BXL U9 ( .AN(n5), .B(n18), .Y(n23) );
  NOR2XL U10 ( .A(state[1]), .B(state[0]), .Y(n28) );
  NAND3XL U11 ( .A(n27), .B(n34), .C(state[0]), .Y(n32) );
  OR2X1 U12 ( .A(n18), .B(n19), .Y(n17) );
  NOR2X1 U13 ( .A(n18), .B(n19), .Y(n16) );
  AOI31X1 U14 ( .A0(n26), .A1(n20), .A2(n21), .B0(n22), .Y(n37) );
  INVX1 U15 ( .A(n27), .Y(n22) );
  NAND4BXL U16 ( .AN(last_block), .B(n5), .C(n11), .D(n10), .Y(n24) );
  AND4X1 U17 ( .A(n13), .B(n14), .C(n25), .D(n2), .Y(first_block_core) );
  NOR4BX1 U18 ( .AN(n1), .B(n3), .C(n4), .D(n12), .Y(n25) );
  INVX1 U19 ( .A(n28), .Y(busy) );
  OAI32X1 U20 ( .A0(n29), .A1(reset), .A2(n30), .B0(n31), .B1(n32), .Y(N14) );
  AND4X1 U21 ( .A(n33), .B(n20), .C(n11), .D(n6), .Y(n30) );
  INVX1 U22 ( .A(n19), .Y(n20) );
  NOR3X1 U23 ( .A(n5), .B(n26), .C(n10), .Y(n33) );
  INVX1 U24 ( .A(inner_busy), .Y(n29) );
  OAI2BB1X1 U25 ( .A0N(n31), .A1N(n38), .B0(n35), .Y(N13) );
  NAND3X1 U26 ( .A(n27), .B(n28), .C(first_block), .Y(n35) );
  INVX1 U27 ( .A(n32), .Y(n38) );
  NAND4X1 U28 ( .A(n14), .B(n13), .C(n4), .D(n36), .Y(n31) );
  NOR4BBX1 U30 ( .AN(n1), .BN(n2), .C(n12), .D(n3), .Y(n36) );
endmodule


module top ( clk, reset, data, write_enable, last_block, first_block, busy, 
        digest, output_valid );
  input [7:0] data;
  output [3:0] digest;
  input clk, reset, write_enable, last_block, first_block;
  output busy, output_valid;
  wire   inner_busy, first_block_core, output_enable;
  wire   [31:0] Wt;

  message_schedule our_message_schedule ( .clk(clk), .reset(reset), .data(data), .write_enable(write_enable), .inner_busy(inner_busy), .Wt(Wt) );
  hash_core our_hash_core ( .clk(clk), .reset(reset), .Wt(Wt), .inner_busy(
        inner_busy), .first_block_core(first_block_core), .output_enable(
        output_enable), .digest(digest), .output_valid(output_valid) );
  controller our_controller ( .clk(clk), .reset(reset), .first_block(
        first_block), .last_block(last_block), .output_enable(output_enable), 
        .busy(busy), .inner_busy(inner_busy), .first_block_core(
        first_block_core) );
endmodule


module sha256_chip ( clk, reset, data, write_enable, last_block, first_block, 
        busy, digest, output_valid );
  input [7:0] data;
  output [3:0] digest;
  input clk, reset, write_enable, last_block, first_block;
  output busy, output_valid;
  wire   net_clk, net_reset, net_write_enable, net_last_block, net_first_block,
         net_busy, net_output_valid;
  wire   [7:0] net_data;
  wire   [3:0] net_digest;

  PIW PIW_clk ( .PAD(clk), .C(net_clk) );
  PIW PIW_reset ( .PAD(reset), .C(net_reset) );
  PIW PIW_data0 ( .PAD(data[0]), .C(net_data[0]) );
  PIW PIW_data1 ( .PAD(data[1]), .C(net_data[1]) );
  PIW PIW_data2 ( .PAD(data[2]), .C(net_data[2]) );
  PIW PIW_data3 ( .PAD(data[3]), .C(net_data[3]) );
  PIW PIW_data4 ( .PAD(data[4]), .C(net_data[4]) );
  PIW PIW_data5 ( .PAD(data[5]), .C(net_data[5]) );
  PIW PIW_data6 ( .PAD(data[6]), .C(net_data[6]) );
  PIW PIW_data7 ( .PAD(data[7]), .C(net_data[7]) );
  PIW PIW_write_enable ( .PAD(write_enable), .C(net_write_enable) );
  PIW PIW_last_block ( .PAD(last_block), .C(net_last_block) );
  PIW PIW_first_block ( .PAD(first_block), .C(net_first_block) );
  PO8W PO8W_busy ( .I(net_busy), .PAD(busy) );
  PO8W PO8W_digest0 ( .I(net_digest[0]), .PAD(digest[0]) );
  PO8W PO8W_digest1 ( .I(net_digest[1]), .PAD(digest[1]) );
  PO8W PO8W_digest2 ( .I(net_digest[2]), .PAD(digest[2]) );
  PO8W PO8W_digest3 ( .I(net_digest[3]), .PAD(digest[3]) );
  PO8W PO8W_output_valid ( .I(net_output_valid), .PAD(output_valid) );
  top inst_top ( .clk(net_clk), .reset(net_reset), .data(net_data), 
        .write_enable(net_write_enable), .last_block(net_last_block), 
        .first_block(net_first_block), .busy(net_busy), .digest(net_digest), 
        .output_valid(net_output_valid) );
endmodule

